* NGSPICE file created from mkQF100SPI.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

.subckt mkQF100SPI CLK RST_N VGND VPWR slave_ack_o slave_adr_i[0] slave_adr_i[10]
+ slave_adr_i[11] slave_adr_i[12] slave_adr_i[13] slave_adr_i[14] slave_adr_i[15]
+ slave_adr_i[16] slave_adr_i[17] slave_adr_i[18] slave_adr_i[19] slave_adr_i[1] slave_adr_i[20]
+ slave_adr_i[21] slave_adr_i[22] slave_adr_i[23] slave_adr_i[24] slave_adr_i[25]
+ slave_adr_i[26] slave_adr_i[27] slave_adr_i[28] slave_adr_i[29] slave_adr_i[2] slave_adr_i[30]
+ slave_adr_i[31] slave_adr_i[3] slave_adr_i[4] slave_adr_i[5] slave_adr_i[6] slave_adr_i[7]
+ slave_adr_i[8] slave_adr_i[9] slave_cyc_i slave_dat_i[0] slave_dat_i[10] slave_dat_i[11]
+ slave_dat_i[12] slave_dat_i[13] slave_dat_i[14] slave_dat_i[15] slave_dat_i[16]
+ slave_dat_i[17] slave_dat_i[18] slave_dat_i[19] slave_dat_i[1] slave_dat_i[20] slave_dat_i[21]
+ slave_dat_i[22] slave_dat_i[23] slave_dat_i[24] slave_dat_i[25] slave_dat_i[26]
+ slave_dat_i[27] slave_dat_i[28] slave_dat_i[29] slave_dat_i[2] slave_dat_i[30] slave_dat_i[31]
+ slave_dat_i[3] slave_dat_i[4] slave_dat_i[5] slave_dat_i[6] slave_dat_i[7] slave_dat_i[8]
+ slave_dat_i[9] slave_dat_o[0] slave_dat_o[10] slave_dat_o[11] slave_dat_o[12] slave_dat_o[13]
+ slave_dat_o[14] slave_dat_o[15] slave_dat_o[16] slave_dat_o[17] slave_dat_o[18]
+ slave_dat_o[19] slave_dat_o[1] slave_dat_o[20] slave_dat_o[21] slave_dat_o[22] slave_dat_o[23]
+ slave_dat_o[24] slave_dat_o[25] slave_dat_o[26] slave_dat_o[27] slave_dat_o[28]
+ slave_dat_o[29] slave_dat_o[2] slave_dat_o[30] slave_dat_o[31] slave_dat_o[3] slave_dat_o[4]
+ slave_dat_o[5] slave_dat_o[6] slave_dat_o[7] slave_dat_o[8] slave_dat_o[9] slave_err_o
+ slave_rty_o slave_sel_i[0] slave_sel_i[1] slave_sel_i[2] slave_sel_i[3] slave_stb_i
+ slave_we_i spiMaster_miso spiMaster_mosi spiMaster_mosi_oe spiMaster_sclk
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1270_ _1521_/A _1270_/B VGND VGND VPWR VPWR _1271_/A sky130_fd_sc_hd__and2_1
X_1606_ _1606_/A _1606_/B _1606_/C VGND VGND VPWR VPWR _1607_/A sky130_fd_sc_hd__and3_1
X_0985_ _0985_/A VGND VGND VPWR VPWR _0985_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1537_ _1551_/A _1585_/B VGND VGND VPWR VPWR _1538_/S sky130_fd_sc_hd__nor2_1
X_1468_ _1626_/Q _1608_/B VGND VGND VPWR VPWR _1468_/X sky130_fd_sc_hd__or2_1
X_1399_ _1429_/B VGND VGND VPWR VPWR _1459_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_42_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1322_ _1321_/A _1321_/B _1321_/C VGND VGND VPWR VPWR _1323_/C sky130_fd_sc_hd__o21ai_1
X_1253_ input20/X _1231_/X _1102_/A _1667_/Q VGND VGND VPWR VPWR _1254_/B sky130_fd_sc_hd__o22a_1
X_1184_ _1184_/A VGND VGND VPWR VPWR _1647_/D sky130_fd_sc_hd__clkbuf_1
X_0968_ _1709_/Q _1069_/A _0967_/X _1693_/Q VGND VGND VPWR VPWR _1418_/A sky130_fd_sc_hd__a22oi_2
X_0899_ _1568_/B _0891_/X _0896_/X _1551_/A VGND VGND VPWR VPWR _0900_/C sky130_fd_sc_hd__a211o_1
XFILLER_23_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0822_ _1682_/Q _1337_/A _1331_/A _1681_/Q VGND VGND VPWR VPWR _0841_/B sky130_fd_sc_hd__a22o_1
XFILLER_9_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1305_ _1305_/A _1305_/B VGND VGND VPWR VPWR _1677_/D sky130_fd_sc_hd__nor2_1
X_1236_ _1251_/A _1236_/B VGND VGND VPWR VPWR _1237_/A sky130_fd_sc_hd__and2_1
X_1098_ _1098_/A VGND VGND VPWR VPWR _1411_/A sky130_fd_sc_hd__clkbuf_2
X_1167_ input24/X _1159_/X _1139_/X _1643_/Q VGND VGND VPWR VPWR _1168_/B sky130_fd_sc_hd__o22a_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1021_ _1726_/Q _1029_/B _1029_/C VGND VGND VPWR VPWR _1022_/A sky130_fd_sc_hd__and3_1
X_0805_ _1289_/A VGND VGND VPWR VPWR _1509_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1219_ _1233_/A _1219_/B VGND VGND VPWR VPWR _1220_/A sky130_fd_sc_hd__or2_1
XFILLER_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_5 slave_adr_i[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1570_ _1759_/Q _1542_/X _1569_/X _1546_/X VGND VGND VPWR VPWR _1571_/B sky130_fd_sc_hd__a22o_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1004_ _1004_/A VGND VGND VPWR VPWR _1004_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1699_ _1730_/CLK _1699_/D VGND VGND VPWR VPWR _1699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput64 _1004_/X VGND VGND VPWR VPWR slave_dat_o[18] sky130_fd_sc_hd__buf_2
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput75 _1028_/X VGND VGND VPWR VPWR slave_dat_o[28] sky130_fd_sc_hd__buf_2
XFILLER_48_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput86 _0974_/X VGND VGND VPWR VPWR slave_dat_o[9] sky130_fd_sc_hd__buf_2
XFILLER_31_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1622_ _1767_/CLK _1622_/D VGND VGND VPWR VPWR _1622_/Q sky130_fd_sc_hd__dfxtp_1
X_1553_ _1756_/Q _1542_/X _1552_/X _1546_/X VGND VGND VPWR VPWR _1554_/B sky130_fd_sc_hd__a22o_1
X_1484_ _1743_/Q _1480_/Y _1744_/Q VGND VGND VPWR VPWR _1484_/X sky130_fd_sc_hd__a21o_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_5_0_CLK clkbuf_4_5_0_CLK/A VGND VGND VPWR VPWR _1740_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0984_ _1424_/A _1005_/C VGND VGND VPWR VPWR _0985_/A sky130_fd_sc_hd__and2b_1
X_1536_ _1536_/A _1550_/A _1600_/B _1536_/D VGND VGND VPWR VPWR _1585_/B sky130_fd_sc_hd__or4_1
X_1605_ _1735_/Q _1442_/A _1509_/B _1766_/Q VGND VGND VPWR VPWR _1606_/C sky130_fd_sc_hd__a31o_1
X_1398_ input1/X _1427_/B VGND VGND VPWR VPWR _1429_/B sky130_fd_sc_hd__nand2_1
X_1467_ _0879_/B _1080_/X _1466_/X _1279_/X VGND VGND VPWR VPWR _1737_/D sky130_fd_sc_hd__o211a_1
XFILLER_10_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1321_ _1321_/A _1321_/B _1321_/C VGND VGND VPWR VPWR _1333_/A sky130_fd_sc_hd__or3_2
X_1252_ _1252_/A VGND VGND VPWR VPWR _1666_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1183_ _1197_/A _1183_/B VGND VGND VPWR VPWR _1184_/A sky130_fd_sc_hd__or2_1
X_0967_ _0967_/A VGND VGND VPWR VPWR _0967_/X sky130_fd_sc_hd__buf_2
X_0898_ _1557_/D VGND VGND VPWR VPWR _1551_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1519_ _1508_/X _1751_/Q _1519_/S VGND VGND VPWR VPWR _1519_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0821_ _1681_/Q _1331_/A _1325_/A _1680_/Q VGND VGND VPWR VPWR _0841_/A sky130_fd_sc_hd__o22a_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1304_ _1298_/X _1300_/X _1302_/Y _1342_/B VGND VGND VPWR VPWR _1305_/B sky130_fd_sc_hd__o22a_1
X_1235_ input15/X _1206_/X _1207_/X _1662_/Q VGND VGND VPWR VPWR _1236_/B sky130_fd_sc_hd__a22o_1
X_1166_ _1411_/A VGND VGND VPWR VPWR _1197_/A sky130_fd_sc_hd__clkbuf_1
X_1097_ _1097_/A VGND VGND VPWR VPWR _1624_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1020_ _1020_/A VGND VGND VPWR VPWR _1029_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0804_ _1749_/Q VGND VGND VPWR VPWR _1289_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1218_ input9/X _1195_/X _1211_/X _1657_/Q VGND VGND VPWR VPWR _1219_/B sky130_fd_sc_hd__o22a_1
X_1149_ _1256_/A VGND VGND VPWR VPWR _1180_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_6 slave_adr_i[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1003_ _1719_/Q _1433_/A _1005_/C VGND VGND VPWR VPWR _1004_/A sky130_fd_sc_hd__and3_1
X_1767_ _1767_/CLK _1767_/D VGND VGND VPWR VPWR _1767_/Q sky130_fd_sc_hd__dfxtp_1
X_1698_ _1730_/CLK _1698_/D VGND VGND VPWR VPWR _1698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput65 _1006_/X VGND VGND VPWR VPWR slave_dat_o[19] sky130_fd_sc_hd__buf_2
XFILLER_0_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput54 _1411_/B VGND VGND VPWR VPWR slave_ack_o sky130_fd_sc_hd__buf_2
Xoutput76 _1030_/X VGND VGND VPWR VPWR slave_dat_o[29] sky130_fd_sc_hd__buf_2
Xoutput87 _0901_/X VGND VGND VPWR VPWR spiMaster_mosi sky130_fd_sc_hd__buf_2
XFILLER_48_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1552_ _1756_/Q _1524_/X _1552_/S VGND VGND VPWR VPWR _1552_/X sky130_fd_sc_hd__mux2_1
X_1621_ _1733_/CLK _1621_/D VGND VGND VPWR VPWR _1621_/Q sky130_fd_sc_hd__dfxtp_1
X_1483_ _1480_/Y _1482_/Y _1083_/X VGND VGND VPWR VPWR _1743_/D sky130_fd_sc_hd__o21a_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0983_ _1020_/A VGND VGND VPWR VPWR _1005_/C sky130_fd_sc_hd__clkbuf_1
X_1604_ _1604_/A VGND VGND VPWR VPWR _1765_/D sky130_fd_sc_hd__clkbuf_1
X_1535_ _1535_/A VGND VGND VPWR VPWR _1753_/D sky130_fd_sc_hd__clkbuf_1
X_1397_ _1397_/A VGND VGND VPWR VPWR _1701_/D sky130_fd_sc_hd__clkbuf_1
X_1466_ _1631_/Q _1608_/B VGND VGND VPWR VPWR _1466_/X sky130_fd_sc_hd__or2_1
XFILLER_35_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1320_ _1680_/Q _1319_/Y _1486_/A VGND VGND VPWR VPWR _1321_/C sky130_fd_sc_hd__mux2_1
Xclkbuf_4_4_0_CLK clkbuf_4_5_0_CLK/A VGND VGND VPWR VPWR _1742_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_5_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1251_ _1251_/A _1251_/B VGND VGND VPWR VPWR _1252_/A sky130_fd_sc_hd__and2_1
X_1182_ input30/X _1159_/X _1175_/X _1647_/Q VGND VGND VPWR VPWR _1183_/B sky130_fd_sc_hd__o22a_1
XFILLER_24_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0897_ _1301_/A _0897_/B _0897_/C VGND VGND VPWR VPWR _1557_/D sky130_fd_sc_hd__nor3_2
X_0966_ _0966_/A VGND VGND VPWR VPWR _1069_/A sky130_fd_sc_hd__buf_2
X_1518_ _1531_/A _1568_/B _1590_/C _1551_/A VGND VGND VPWR VPWR _1519_/S sky130_fd_sc_hd__or4_1
X_1449_ _1726_/Q _1433_/X _1434_/X VGND VGND VPWR VPWR _1726_/D sky130_fd_sc_hd__a21o_1
XFILLER_15_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0820_ _0946_/A _0828_/A _0826_/A VGND VGND VPWR VPWR _1325_/A sky130_fd_sc_hd__or3b_2
X_1303_ _1338_/S VGND VGND VPWR VPWR _1342_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1234_ _1234_/A VGND VGND VPWR VPWR _1661_/D sky130_fd_sc_hd__clkbuf_1
X_1096_ _1107_/A _1096_/B VGND VGND VPWR VPWR _1097_/A sky130_fd_sc_hd__and2_1
X_1165_ _1165_/A VGND VGND VPWR VPWR _1642_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0949_ _0949_/A VGND VGND VPWR VPWR _0949_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_47_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0803_ _1395_/A VGND VGND VPWR VPWR _1411_/B sky130_fd_sc_hd__inv_2
XFILLER_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1217_ _1217_/A VGND VGND VPWR VPWR _1656_/D sky130_fd_sc_hd__clkbuf_1
X_1079_ _1346_/A _1079_/B _1079_/C VGND VGND VPWR VPWR _1080_/A sky130_fd_sc_hd__and3_1
X_1148_ _1148_/A VGND VGND VPWR VPWR _1637_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_7 slave_adr_i[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1002_ _1002_/A VGND VGND VPWR VPWR _1002_/X sky130_fd_sc_hd__clkbuf_1
X_1766_ _1766_/CLK _1766_/D VGND VGND VPWR VPWR _1766_/Q sky130_fd_sc_hd__dfxtp_1
X_1697_ _1730_/CLK _1697_/D VGND VGND VPWR VPWR _1697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput88 _0903_/Y VGND VGND VPWR VPWR spiMaster_mosi_oe sky130_fd_sc_hd__buf_2
Xoutput77 _0939_/X VGND VGND VPWR VPWR slave_dat_o[2] sky130_fd_sc_hd__buf_2
Xoutput55 _0926_/X VGND VGND VPWR VPWR slave_dat_o[0] sky130_fd_sc_hd__buf_2
XFILLER_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput66 _0931_/X VGND VGND VPWR VPWR slave_dat_o[1] sky130_fd_sc_hd__buf_2
XFILLER_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1551_ _1551_/A _1595_/B VGND VGND VPWR VPWR _1552_/S sky130_fd_sc_hd__nor2_1
X_1482_ _1491_/A _1509_/B _1471_/Y _1481_/Y VGND VGND VPWR VPWR _1482_/Y sky130_fd_sc_hd__a31oi_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1620_ _1742_/CLK _1620_/D VGND VGND VPWR VPWR _1620_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1749_ _1766_/CLK _1749_/D VGND VGND VPWR VPWR _1749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0982_ _1713_/Q _1069_/A _0967_/X _1697_/Q VGND VGND VPWR VPWR _1424_/A sky130_fd_sc_hd__a22oi_4
X_1534_ _1554_/A _1534_/B VGND VGND VPWR VPWR _1535_/A sky130_fd_sc_hd__and2_1
X_1603_ _1603_/A _1603_/B VGND VGND VPWR VPWR _1604_/A sky130_fd_sc_hd__and2_1
X_1465_ _1736_/Q _1080_/X _1464_/X _1279_/X VGND VGND VPWR VPWR _1736_/D sky130_fd_sc_hd__o211a_1
XFILLER_27_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1396_ _1402_/A _1427_/B _1396_/C VGND VGND VPWR VPWR _1397_/A sky130_fd_sc_hd__and3_1
XFILLER_10_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1250_ input19/X _1242_/X _1243_/X _1666_/Q VGND VGND VPWR VPWR _1251_/B sky130_fd_sc_hd__a22o_1
X_1181_ _1181_/A VGND VGND VPWR VPWR _1646_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0896_ _1563_/C _0892_/X _0895_/X _1590_/B VGND VGND VPWR VPWR _0896_/X sky130_fd_sc_hd__o211a_1
X_0965_ _0965_/A VGND VGND VPWR VPWR _0965_/X sky130_fd_sc_hd__clkbuf_1
X_1517_ _1517_/A VGND VGND VPWR VPWR _1750_/D sky130_fd_sc_hd__clkbuf_1
X_1448_ _1448_/A VGND VGND VPWR VPWR _1725_/D sky130_fd_sc_hd__clkbuf_1
X_1379_ _1759_/Q _1368_/X _1378_/X _1633_/Q _1375_/X VGND VGND VPWR VPWR _1379_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1302_ _0844_/X _1536_/A _0833_/X VGND VGND VPWR VPWR _1302_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1233_ _1233_/A _1233_/B VGND VGND VPWR VPWR _1234_/A sky130_fd_sc_hd__or2_1
X_1095_ input35/X _1092_/X _1094_/X _1624_/Q VGND VGND VPWR VPWR _1096_/B sky130_fd_sc_hd__a22o_1
X_1164_ _1180_/A _1164_/B VGND VGND VPWR VPWR _1165_/A sky130_fd_sc_hd__and2_1
X_0948_ _0948_/A _1407_/C VGND VGND VPWR VPWR _0949_/A sky130_fd_sc_hd__and2_1
X_0879_ _1746_/Q _0879_/B VGND VGND VPWR VPWR _1536_/D sky130_fd_sc_hd__xnor2_1
XFILLER_34_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_3_0_CLK clkbuf_4_3_0_CLK/A VGND VGND VPWR VPWR _1733_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_34_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0802_ _1734_/Q _1093_/A _1673_/Q VGND VGND VPWR VPWR _1395_/A sky130_fd_sc_hd__o21ai_2
X_1216_ _1216_/A _1216_/B VGND VGND VPWR VPWR _1217_/A sky130_fd_sc_hd__and2_1
XFILLER_37_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1147_ _1161_/A _1147_/B VGND VGND VPWR VPWR _1148_/A sky130_fd_sc_hd__or2_1
X_1078_ _1070_/Y _1074_/X _1305_/A VGND VGND VPWR VPWR _1621_/D sky130_fd_sc_hd__a21oi_1
XFILLER_29_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_8 slave_adr_i[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1001_ _1718_/Q _1433_/A _1005_/C VGND VGND VPWR VPWR _1002_/A sky130_fd_sc_hd__and3_1
XFILLER_19_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1765_ _1765_/CLK _1765_/D VGND VGND VPWR VPWR _1765_/Q sky130_fd_sc_hd__dfxtp_1
X_1696_ _1765_/CLK _1696_/D VGND VGND VPWR VPWR _1696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput89 _0854_/X VGND VGND VPWR VPWR spiMaster_sclk sky130_fd_sc_hd__buf_2
Xoutput67 _1010_/X VGND VGND VPWR VPWR slave_dat_o[20] sky130_fd_sc_hd__buf_2
Xoutput56 _0977_/X VGND VGND VPWR VPWR slave_dat_o[10] sky130_fd_sc_hd__buf_2
Xoutput78 _1033_/X VGND VGND VPWR VPWR slave_dat_o[30] sky130_fd_sc_hd__buf_2
XFILLER_16_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1481_ _1743_/Q VGND VGND VPWR VPWR _1481_/Y sky130_fd_sc_hd__inv_2
X_1550_ _1550_/A _1600_/B _1550_/C VGND VGND VPWR VPWR _1595_/B sky130_fd_sc_hd__or3_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1748_ _1766_/CLK _1748_/D VGND VGND VPWR VPWR _1748_/Q sky130_fd_sc_hd__dfxtp_1
X_1679_ _1740_/CLK _1679_/D VGND VGND VPWR VPWR _1679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0981_ _0981_/A VGND VGND VPWR VPWR _0981_/X sky130_fd_sc_hd__clkbuf_1
X_1602_ _1765_/Q _1573_/A _1601_/X _1576_/A VGND VGND VPWR VPWR _1603_/B sky130_fd_sc_hd__a22o_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1533_ _1753_/Q _1507_/X _1532_/X _1514_/X VGND VGND VPWR VPWR _1534_/B sky130_fd_sc_hd__a22o_1
X_1464_ _1635_/Q _1608_/B VGND VGND VPWR VPWR _1464_/X sky130_fd_sc_hd__or2_1
X_1395_ _1395_/A VGND VGND VPWR VPWR _1427_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1180_ _1180_/A _1180_/B VGND VGND VPWR VPWR _1181_/A sky130_fd_sc_hd__and2_1
X_0964_ _0980_/A _1415_/A VGND VGND VPWR VPWR _0965_/A sky130_fd_sc_hd__and2_1
X_1516_ _1521_/A _1516_/B VGND VGND VPWR VPWR _1517_/A sky130_fd_sc_hd__and2_1
X_0895_ _1687_/Q _0892_/S _0893_/X _1550_/C VGND VGND VPWR VPWR _0895_/X sky130_fd_sc_hd__a211o_1
X_1447_ _1725_/Q _1456_/B _1456_/C VGND VGND VPWR VPWR _1448_/A sky130_fd_sc_hd__and3_1
X_1378_ _1378_/A VGND VGND VPWR VPWR _1378_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1301_ _1301_/A VGND VGND VPWR VPWR _1536_/A sky130_fd_sc_hd__clkbuf_2
X_1232_ input14/X _1231_/X _1211_/X _1661_/Q VGND VGND VPWR VPWR _1233_/B sky130_fd_sc_hd__o22a_1
X_1094_ _1243_/A VGND VGND VPWR VPWR _1094_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1163_ input13/X _1134_/X _1135_/X _1642_/Q VGND VGND VPWR VPWR _1164_/B sky130_fd_sc_hd__a22o_1
X_0947_ _1705_/Q _0997_/A _0967_/A _1689_/Q _0946_/X VGND VGND VPWR VPWR _1407_/C
+ sky130_fd_sc_hd__a221o_1
X_0878_ _1696_/Q _1695_/Q _0892_/S VGND VGND VPWR VPWR _0878_/X sky130_fd_sc_hd__mux2_1
X_0801_ _1348_/A VGND VGND VPWR VPWR _1093_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1146_ input39/X _1123_/X _1139_/X _1637_/Q VGND VGND VPWR VPWR _1147_/B sky130_fd_sc_hd__o22a_1
X_1215_ input8/X _1206_/X _1207_/X _1656_/Q VGND VGND VPWR VPWR _1216_/B sky130_fd_sc_hd__a22o_1
XFILLER_37_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1077_ _1502_/A VGND VGND VPWR VPWR _1305_/A sky130_fd_sc_hd__buf_2
XFILLER_45_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_9 slave_adr_i[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1000_ _1000_/A VGND VGND VPWR VPWR _1000_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1764_ _1765_/CLK _1764_/D VGND VGND VPWR VPWR _1764_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_4_2_0_CLK clkbuf_4_3_0_CLK/A VGND VGND VPWR VPWR _1671_/CLK sky130_fd_sc_hd__clkbuf_2
X_1695_ _1730_/CLK _1695_/D VGND VGND VPWR VPWR _1695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1129_ _1129_/A VGND VGND VPWR VPWR _1632_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput57 _0981_/X VGND VGND VPWR VPWR slave_dat_o[11] sky130_fd_sc_hd__buf_2
XFILLER_0_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput79 _1035_/X VGND VGND VPWR VPWR slave_dat_o[31] sky130_fd_sc_hd__buf_2
Xoutput68 _1012_/X VGND VGND VPWR VPWR slave_dat_o[21] sky130_fd_sc_hd__buf_2
X_1480_ _1623_/Q _1622_/Q _1606_/B VGND VGND VPWR VPWR _1480_/Y sky130_fd_sc_hd__a21oi_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1678_ _1740_/CLK _1678_/D VGND VGND VPWR VPWR _1678_/Q sky130_fd_sc_hd__dfxtp_1
X_1747_ _1752_/CLK _1747_/D VGND VGND VPWR VPWR _1747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0980_ _0980_/A _1422_/A VGND VGND VPWR VPWR _0981_/A sky130_fd_sc_hd__and2_1
XFILLER_16_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1532_ _1508_/X _1753_/Q _1532_/S VGND VGND VPWR VPWR _1532_/X sky130_fd_sc_hd__mux2_1
X_1601_ _1562_/X _1765_/Q _1601_/S VGND VGND VPWR VPWR _1601_/X sky130_fd_sc_hd__mux2_1
X_1463_ _1461_/X _1462_/Y _1083_/X VGND VGND VPWR VPWR _1735_/D sky130_fd_sc_hd__o21a_1
X_1394_ _1700_/Q _1381_/A _1393_/X VGND VGND VPWR VPWR _1700_/D sky130_fd_sc_hd__o21a_1
XFILLER_41_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0894_ _0894_/A _1536_/D VGND VGND VPWR VPWR _1550_/C sky130_fd_sc_hd__nand2_1
XFILLER_32_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0963_ _1708_/Q _1272_/B _0961_/X _0962_/X VGND VGND VPWR VPWR _1415_/A sky130_fd_sc_hd__o22a_1
X_1515_ _1750_/Q _1507_/X _1512_/X _1514_/X VGND VGND VPWR VPWR _1516_/B sky130_fd_sc_hd__a22o_1
X_1377_ _1693_/Q _1367_/X _1376_/X VGND VGND VPWR VPWR _1693_/D sky130_fd_sc_hd__o21a_1
X_1446_ _1724_/Q _1433_/X _1434_/X VGND VGND VPWR VPWR _1724_/D sky130_fd_sc_hd__a21o_1
XFILLER_23_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1300_ _1477_/A _1475_/A _1473_/A _1338_/S _1299_/X VGND VGND VPWR VPWR _1300_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_1_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1231_ _1231_/A VGND VGND VPWR VPWR _1231_/X sky130_fd_sc_hd__clkbuf_2
X_1162_ _1162_/A VGND VGND VPWR VPWR _1641_/D sky130_fd_sc_hd__clkbuf_1
X_1093_ _1093_/A _1093_/B VGND VGND VPWR VPWR _1243_/A sky130_fd_sc_hd__nor2_2
X_0877_ _1600_/D VGND VGND VPWR VPWR _1595_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0946_ _0946_/A _0993_/B _0993_/C VGND VGND VPWR VPWR _0946_/X sky130_fd_sc_hd__and3_1
X_1429_ _1429_/A _1429_/B VGND VGND VPWR VPWR _1430_/A sky130_fd_sc_hd__or2_1
XFILLER_18_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0800_ _0787_/Y _0798_/X _1079_/B VGND VGND VPWR VPWR _1348_/A sky130_fd_sc_hd__o21a_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1214_ _1214_/A VGND VGND VPWR VPWR _1655_/D sky130_fd_sc_hd__clkbuf_1
X_1145_ _1145_/A VGND VGND VPWR VPWR _1636_/D sky130_fd_sc_hd__clkbuf_1
X_1076_ _1098_/A VGND VGND VPWR VPWR _1502_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0929_ _1702_/Q _0928_/X _0955_/A VGND VGND VPWR VPWR _1400_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1763_ _1765_/CLK _1763_/D VGND VGND VPWR VPWR _1763_/Q sky130_fd_sc_hd__dfxtp_1
X_1694_ _1765_/CLK _1694_/D VGND VGND VPWR VPWR _1694_/Q sky130_fd_sc_hd__dfxtp_1
X_1128_ _1144_/A _1128_/B VGND VGND VPWR VPWR _1129_/A sky130_fd_sc_hd__and2_1
X_1059_ _1402_/A _1616_/Q _1274_/B VGND VGND VPWR VPWR _1060_/A sky130_fd_sc_hd__and3_1
XFILLER_0_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput58 _0985_/X VGND VGND VPWR VPWR slave_dat_o[12] sky130_fd_sc_hd__buf_2
Xoutput69 _1014_/X VGND VGND VPWR VPWR slave_dat_o[22] sky130_fd_sc_hd__buf_2
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1746_ _1766_/CLK _1746_/D VGND VGND VPWR VPWR _1746_/Q sky130_fd_sc_hd__dfxtp_2
X_1677_ _1766_/CLK _1677_/D VGND VGND VPWR VPWR _1677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_1_0_CLK clkbuf_4_1_0_CLK/A VGND VGND VPWR VPWR _1650_/CLK sky130_fd_sc_hd__clkbuf_2
X_1531_ _1531_/A _1568_/B _1580_/C _1557_/D VGND VGND VPWR VPWR _1532_/S sky130_fd_sc_hd__or4_1
X_1462_ _1462_/A _1462_/B VGND VGND VPWR VPWR _1462_/Y sky130_fd_sc_hd__nor2_1
X_1600_ _1600_/A _1600_/B _1600_/C _1600_/D VGND VGND VPWR VPWR _1601_/S sky130_fd_sc_hd__or4_1
X_1393_ _1765_/Q _1382_/A _1378_/A _1639_/Q _1048_/A VGND VGND VPWR VPWR _1393_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1729_ _1732_/CLK _1729_/D VGND VGND VPWR VPWR _1729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0893_ _1688_/Q _0900_/A _1550_/A VGND VGND VPWR VPWR _0893_/X sky130_fd_sc_hd__and3_1
X_0962_ _0879_/B _1079_/C _0927_/B _1509_/A _0966_/A VGND VGND VPWR VPWR _0962_/X
+ sky130_fd_sc_hd__a221o_1
X_1445_ _1445_/A VGND VGND VPWR VPWR _1723_/D sky130_fd_sc_hd__clkbuf_1
X_1514_ _1576_/A VGND VGND VPWR VPWR _1514_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1376_ _1758_/Q _1368_/X _1364_/X _1632_/Q _1375_/X VGND VGND VPWR VPWR _1376_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_23_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1230_ _1230_/A VGND VGND VPWR VPWR _1660_/D sky130_fd_sc_hd__clkbuf_1
X_1161_ _1161_/A _1161_/B VGND VGND VPWR VPWR _1162_/A sky130_fd_sc_hd__or2_1
X_1092_ _1242_/A VGND VGND VPWR VPWR _1092_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0876_ _1301_/A _0897_/B _0897_/C VGND VGND VPWR VPWR _1600_/D sky130_fd_sc_hd__or3_2
X_0945_ _0945_/A VGND VGND VPWR VPWR _0945_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1428_ _1428_/A VGND VGND VPWR VPWR _1715_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1359_ _1752_/Q _1352_/X _1462_/B _1626_/Q _1469_/A VGND VGND VPWR VPWR _1359_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1213_ _1233_/A _1213_/B VGND VGND VPWR VPWR _1214_/A sky130_fd_sc_hd__or2_1
XFILLER_37_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1075_ input1/X VGND VGND VPWR VPWR _1098_/A sky130_fd_sc_hd__inv_2
X_1144_ _1144_/A _1144_/B VGND VGND VPWR VPWR _1145_/A sky130_fd_sc_hd__and2_1
X_0859_ _1737_/Q VGND VGND VPWR VPWR _0879_/B sky130_fd_sc_hd__clkbuf_2
X_0928_ _1686_/Q _0961_/B _0989_/C _1675_/Q _0927_/X VGND VGND VPWR VPWR _0928_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1762_ _1762_/CLK _1762_/D VGND VGND VPWR VPWR _1762_/Q sky130_fd_sc_hd__dfxtp_1
X_1693_ _1765_/CLK _1693_/D VGND VGND VPWR VPWR _1693_/Q sky130_fd_sc_hd__dfxtp_1
X_1058_ _1058_/A VGND VGND VPWR VPWR _1615_/D sky130_fd_sc_hd__clkbuf_1
X_1127_ input49/X _1092_/X _1094_/X _1632_/Q VGND VGND VPWR VPWR _1128_/B sky130_fd_sc_hd__a22o_1
Xoutput59 _0988_/X VGND VGND VPWR VPWR slave_dat_o[13] sky130_fd_sc_hd__buf_2
XFILLER_16_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1745_ _1766_/CLK _1745_/D VGND VGND VPWR VPWR _1745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1676_ _1766_/CLK _1676_/D VGND VGND VPWR VPWR _1676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1530_ _1530_/A VGND VGND VPWR VPWR _1752_/D sky130_fd_sc_hd__clkbuf_1
X_1461_ _1766_/Q _1272_/B _1462_/A _1735_/Q VGND VGND VPWR VPWR _1461_/X sky130_fd_sc_hd__o31a_1
X_1392_ _1699_/Q _1381_/X _1391_/X VGND VGND VPWR VPWR _1699_/D sky130_fd_sc_hd__o21a_1
XFILLER_35_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1728_ _1730_/CLK _1728_/D VGND VGND VPWR VPWR _1728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1659_ _1662_/CLK _1659_/D VGND VGND VPWR VPWR _1659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0961_ _1692_/Q _0961_/B VGND VGND VPWR VPWR _0961_/X sky130_fd_sc_hd__and2_1
XFILLER_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0892_ _1686_/Q _1685_/Q _0892_/S VGND VGND VPWR VPWR _0892_/X sky130_fd_sc_hd__mux2_1
X_1513_ _1513_/A _1536_/A VGND VGND VPWR VPWR _1576_/A sky130_fd_sc_hd__nor2_2
XFILLER_4_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1444_ _1723_/Q _1456_/B _1456_/C VGND VGND VPWR VPWR _1445_/A sky130_fd_sc_hd__and3_1
X_1375_ _1375_/A VGND VGND VPWR VPWR _1375_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_0_0_CLK clkbuf_4_1_0_CLK/A VGND VGND VPWR VPWR _1662_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_14_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1160_ input2/X _1159_/X _1139_/X _1641_/Q VGND VGND VPWR VPWR _1161_/B sky130_fd_sc_hd__o22a_1
X_1091_ _1093_/B VGND VGND VPWR VPWR _1242_/A sky130_fd_sc_hd__clkbuf_2
X_0944_ _0948_/A _1405_/A VGND VGND VPWR VPWR _0945_/A sky130_fd_sc_hd__and2_1
XFILLER_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0875_ _1748_/Q _1737_/Q VGND VGND VPWR VPWR _0897_/C sky130_fd_sc_hd__and2b_1
X_1358_ _1686_/Q _1351_/X _1357_/X VGND VGND VPWR VPWR _1686_/D sky130_fd_sc_hd__o21a_1
X_1427_ _1606_/A _1427_/B _1427_/C VGND VGND VPWR VPWR _1428_/A sky130_fd_sc_hd__and3_1
X_1289_ _1289_/A _1289_/B _1766_/Q VGND VGND VPWR VPWR _1289_/X sky130_fd_sc_hd__or3b_2
XFILLER_11_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_7_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_3_7_0_CLK/X sky130_fd_sc_hd__clkbuf_2
X_1212_ input7/X _1195_/X _1211_/X _1655_/Q VGND VGND VPWR VPWR _1213_/B sky130_fd_sc_hd__o22a_1
XFILLER_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1074_ _1195_/A VGND VGND VPWR VPWR _1074_/X sky130_fd_sc_hd__clkbuf_2
X_1143_ input38/X _1134_/X _1135_/X _1636_/Q VGND VGND VPWR VPWR _1144_/B sky130_fd_sc_hd__a22o_1
X_0927_ _1735_/Q _0927_/B VGND VGND VPWR VPWR _0927_/X sky130_fd_sc_hd__and2b_1
X_0858_ _1747_/Q VGND VGND VPWR VPWR _1498_/A sky130_fd_sc_hd__buf_2
XFILLER_20_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0789_ _1644_/Q _1643_/Q _0789_/C VGND VGND VPWR VPWR _1353_/A sky130_fd_sc_hd__nand3_1
XFILLER_45_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1761_ _1762_/CLK _1761_/D VGND VGND VPWR VPWR _1761_/Q sky130_fd_sc_hd__dfxtp_1
X_1692_ _1765_/CLK _1692_/D VGND VGND VPWR VPWR _1692_/Q sky130_fd_sc_hd__dfxtp_1
X_1126_ _1126_/A VGND VGND VPWR VPWR _1631_/D sky130_fd_sc_hd__clkbuf_1
X_1057_ _1615_/Q _1063_/B VGND VGND VPWR VPWR _1058_/A sky130_fd_sc_hd__or2_1
XFILLER_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1744_ _1767_/CLK _1744_/D VGND VGND VPWR VPWR _1744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1675_ _1766_/CLK _1675_/D VGND VGND VPWR VPWR _1675_/Q sky130_fd_sc_hd__dfxtp_1
X_1109_ input44/X _1074_/X _1102_/X _1627_/Q VGND VGND VPWR VPWR _1110_/B sky130_fd_sc_hd__o22a_1
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1460_ _1734_/Q _1272_/B _1439_/C VGND VGND VPWR VPWR _1734_/D sky130_fd_sc_hd__o21a_1
X_1391_ _1764_/Q _1382_/X _1378_/A _1638_/Q _1048_/A VGND VGND VPWR VPWR _1391_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_35_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1658_ _1662_/CLK _1658_/D VGND VGND VPWR VPWR _1658_/Q sky130_fd_sc_hd__dfxtp_1
X_1727_ _1732_/CLK _1727_/D VGND VGND VPWR VPWR _1727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1589_ _1589_/A VGND VGND VPWR VPWR _1762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0960_ _0960_/A VGND VGND VPWR VPWR _0960_/X sky130_fd_sc_hd__clkbuf_1
X_1512_ _1508_/X _1750_/Q _1512_/S VGND VGND VPWR VPWR _1512_/X sky130_fd_sc_hd__mux2_1
X_0891_ _0888_/X _0889_/X _1563_/C VGND VGND VPWR VPWR _0891_/X sky130_fd_sc_hd__mux2_1
X_1443_ _1443_/A VGND VGND VPWR VPWR _1456_/C sky130_fd_sc_hd__clkbuf_1
X_1374_ _1692_/Q _1367_/X _1373_/X VGND VGND VPWR VPWR _1692_/D sky130_fd_sc_hd__o21a_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1090_ _1621_/Q _0909_/A _1071_/Y VGND VGND VPWR VPWR _1093_/B sky130_fd_sc_hd__a21oi_1
X_0874_ _1737_/Q _1288_/B VGND VGND VPWR VPWR _0897_/B sky130_fd_sc_hd__and2b_1
XFILLER_9_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0943_ _1704_/Q _0940_/X _0934_/X _1688_/Q _0942_/X VGND VGND VPWR VPWR _1405_/A
+ sky130_fd_sc_hd__a221o_1
X_1288_ _1747_/Q _1288_/B _1498_/B VGND VGND VPWR VPWR _1288_/X sky130_fd_sc_hd__and3_1
X_1426_ _1426_/A VGND VGND VPWR VPWR _1714_/D sky130_fd_sc_hd__clkbuf_1
X_1357_ _1751_/Q _1352_/X _1462_/B _1625_/Q _1469_/A VGND VGND VPWR VPWR _1357_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1211_ _1211_/A VGND VGND VPWR VPWR _1211_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1142_ _1142_/A VGND VGND VPWR VPWR _1635_/D sky130_fd_sc_hd__clkbuf_1
X_1073_ _1231_/A VGND VGND VPWR VPWR _1195_/A sky130_fd_sc_hd__clkbuf_2
X_0857_ _0894_/A VGND VGND VPWR VPWR _0900_/A sky130_fd_sc_hd__clkbuf_2
X_0926_ _0926_/A VGND VGND VPWR VPWR _0926_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0788_ _1648_/Q _1647_/Q _1646_/Q _1645_/Q VGND VGND VPWR VPWR _0789_/C sky130_fd_sc_hd__nor4_1
X_1409_ _1409_/A _1422_/B VGND VGND VPWR VPWR _1410_/A sky130_fd_sc_hd__or2_1
XFILLER_45_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1760_ _1762_/CLK _1760_/D VGND VGND VPWR VPWR _1760_/Q sky130_fd_sc_hd__dfxtp_1
X_1691_ _1765_/CLK _1691_/D VGND VGND VPWR VPWR _1691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1125_ _1504_/A _1125_/B VGND VGND VPWR VPWR _1126_/A sky130_fd_sc_hd__or2_1
X_1056_ _1056_/A VGND VGND VPWR VPWR _1614_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0909_ _0909_/A VGND VGND VPWR VPWR _1347_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_3_6_0_CLK/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1674_ _1767_/CLK _1674_/D VGND VGND VPWR VPWR _1674_/Q sky130_fd_sc_hd__dfxtp_1
X_1743_ _1767_/CLK _1743_/D VGND VGND VPWR VPWR _1743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1108_ _1108_/A VGND VGND VPWR VPWR _1626_/D sky130_fd_sc_hd__clkbuf_1
X_1039_ _1346_/A _1079_/B VGND VGND VPWR VPWR _1353_/D sky130_fd_sc_hd__nand2_1
XFILLER_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1390_ _1698_/Q _1381_/X _1389_/X VGND VGND VPWR VPWR _1698_/D sky130_fd_sc_hd__o21a_1
XFILLER_35_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1588_ _1603_/A _1588_/B VGND VGND VPWR VPWR _1589_/A sky130_fd_sc_hd__and2_1
X_1657_ _1662_/CLK _1657_/D VGND VGND VPWR VPWR _1657_/Q sky130_fd_sc_hd__dfxtp_1
X_1726_ _1732_/CLK _1726_/D VGND VGND VPWR VPWR _1726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0890_ _1301_/A _1600_/C VGND VGND VPWR VPWR _1563_/C sky130_fd_sc_hd__nor2_1
XFILLER_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1442_ _1442_/A VGND VGND VPWR VPWR _1456_/B sky130_fd_sc_hd__clkbuf_1
X_1511_ _1563_/A _1557_/D _1563_/C _1563_/D VGND VGND VPWR VPWR _1512_/S sky130_fd_sc_hd__or4_1
XFILLER_4_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1373_ _1757_/Q _1368_/X _1364_/X _1631_/Q _1361_/X VGND VGND VPWR VPWR _1373_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_23_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1709_ _1730_/CLK _1709_/D VGND VGND VPWR VPWR _1709_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0873_ _1748_/Q _1736_/Q VGND VGND VPWR VPWR _1288_/B sky130_fd_sc_hd__xnor2_1
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0942_ _0942_/A _0955_/A _1079_/C VGND VGND VPWR VPWR _0942_/X sky130_fd_sc_hd__and3_1
X_1425_ _1425_/A _1429_/B VGND VGND VPWR VPWR _1426_/A sky130_fd_sc_hd__or2_1
X_1287_ _1289_/A _1746_/Q _1745_/Q VGND VGND VPWR VPWR _1498_/B sky130_fd_sc_hd__and3_1
X_1356_ _1685_/Q _1351_/X _1355_/X VGND VGND VPWR VPWR _1685_/D sky130_fd_sc_hd__o21a_1
XFILLER_18_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1210_ _1210_/A VGND VGND VPWR VPWR _1654_/D sky130_fd_sc_hd__clkbuf_1
X_1141_ _1161_/A _1141_/B VGND VGND VPWR VPWR _1142_/A sky130_fd_sc_hd__or2_1
X_1072_ _1621_/Q _0909_/A _1071_/Y VGND VGND VPWR VPWR _1231_/A sky130_fd_sc_hd__a21o_1
X_0856_ _1491_/A _1289_/B VGND VGND VPWR VPWR _0894_/A sky130_fd_sc_hd__nor2_1
X_0925_ _0948_/A _1396_/C VGND VGND VPWR VPWR _0926_/A sky130_fd_sc_hd__and2_1
X_0787_ _1739_/Q VGND VGND VPWR VPWR _0787_/Y sky130_fd_sc_hd__inv_2
X_1408_ _1408_/A VGND VGND VPWR VPWR _1705_/D sky130_fd_sc_hd__clkbuf_1
X_1339_ _1339_/A _1339_/B VGND VGND VPWR VPWR _1339_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1690_ _1765_/CLK _1690_/D VGND VGND VPWR VPWR _1690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1124_ input48/X _1123_/X _1102_/X _1631_/Q VGND VGND VPWR VPWR _1125_/B sky130_fd_sc_hd__o22a_1
X_1055_ _1402_/A _1614_/Q _1274_/B VGND VGND VPWR VPWR _1056_/A sky130_fd_sc_hd__and3_1
XFILLER_33_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0839_ _1473_/A _0825_/X _0830_/A _0951_/A _1475_/A VGND VGND VPWR VPWR _0839_/X
+ sky130_fd_sc_hd__a2111o_1
X_0908_ _0787_/Y _0798_/X _1079_/B VGND VGND VPWR VPWR _0909_/A sky130_fd_sc_hd__o21ai_1
XFILLER_16_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1742_ _1742_/CLK _1742_/D VGND VGND VPWR VPWR _1742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1673_ _1733_/CLK _1673_/D VGND VGND VPWR VPWR _1673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1107_ _1107_/A _1107_/B VGND VGND VPWR VPWR _1108_/A sky130_fd_sc_hd__and2_1
X_1038_ _1640_/Q VGND VGND VPWR VPWR _1346_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1725_ _1732_/CLK _1725_/D VGND VGND VPWR VPWR _1725_/Q sky130_fd_sc_hd__dfxtp_1
X_1587_ _1762_/Q _1573_/X _1586_/X _1576_/X VGND VGND VPWR VPWR _1588_/B sky130_fd_sc_hd__a22o_1
X_1656_ _1671_/CLK _1656_/D VGND VGND VPWR VPWR _1656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_5_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_3_5_0_CLK/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1510_ _1536_/A _1600_/B VGND VGND VPWR VPWR _1563_/D sky130_fd_sc_hd__nor2_1
X_1441_ _1722_/Q _1433_/X _1434_/X VGND VGND VPWR VPWR _1722_/D sky130_fd_sc_hd__a21o_1
XFILLER_4_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1372_ _1691_/Q _1367_/X _1371_/X VGND VGND VPWR VPWR _1691_/D sky130_fd_sc_hd__o21a_1
X_1708_ _1712_/CLK _1708_/D VGND VGND VPWR VPWR _1708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1639_ _1732_/CLK _1639_/D VGND VGND VPWR VPWR _1639_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_14_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0941_ _0989_/C VGND VGND VPWR VPWR _1079_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_0872_ _1289_/A _1509_/B VGND VGND VPWR VPWR _1301_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1424_ _1424_/A _1459_/B VGND VGND VPWR VPWR _1713_/D sky130_fd_sc_hd__nor2_1
X_1355_ _1750_/Q _1352_/X _1462_/B _1624_/Q _1469_/A VGND VGND VPWR VPWR _1355_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_48_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1286_ _1286_/A _1286_/B _1286_/C _1285_/X VGND VGND VPWR VPWR _1348_/B sky130_fd_sc_hd__or4b_2
XFILLER_40_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1140_ input37/X _1123_/X _1139_/X _1635_/Q VGND VGND VPWR VPWR _1141_/B sky130_fd_sc_hd__o22a_1
X_1071_ _1673_/Q _1071_/B _1071_/C VGND VGND VPWR VPWR _1071_/Y sky130_fd_sc_hd__nand3b_1
X_0924_ _1701_/Q _0955_/A _0918_/X _0923_/X VGND VGND VPWR VPWR _1396_/C sky130_fd_sc_hd__o22a_1
X_0855_ _1289_/A VGND VGND VPWR VPWR _1491_/A sky130_fd_sc_hd__inv_2
X_1338_ _0808_/X _1337_/Y _1338_/S VGND VGND VPWR VPWR _1339_/B sky130_fd_sc_hd__mux2_1
XFILLER_29_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1407_ _1606_/A _1427_/B _1407_/C VGND VGND VPWR VPWR _1408_/A sky130_fd_sc_hd__and3_1
X_1269_ input26/X _1242_/X _1243_/X _1672_/Q VGND VGND VPWR VPWR _1270_/B sky130_fd_sc_hd__a22o_1
XFILLER_3_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1123_ _1195_/A VGND VGND VPWR VPWR _1123_/X sky130_fd_sc_hd__clkbuf_2
X_1054_ _1276_/A VGND VGND VPWR VPWR _1274_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_0907_ _0921_/A _1640_/Q _0916_/A VGND VGND VPWR VPWR _0907_/X sky130_fd_sc_hd__a21o_1
X_0838_ _0838_/A VGND VGND VPWR VPWR _1475_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1741_ _1742_/CLK _1741_/D VGND VGND VPWR VPWR _1741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1672_ _1717_/CLK _1672_/D VGND VGND VPWR VPWR _1672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1106_ input43/X _1092_/X _1094_/X _1626_/Q VGND VGND VPWR VPWR _1107_/B sky130_fd_sc_hd__a22o_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1037_ _1375_/A VGND VGND VPWR VPWR _1048_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1724_ _1732_/CLK _1724_/D VGND VGND VPWR VPWR _1724_/Q sky130_fd_sc_hd__dfxtp_1
X_1586_ _1762_/Q _1524_/X _1586_/S VGND VGND VPWR VPWR _1586_/X sky130_fd_sc_hd__mux2_1
X_1655_ _1662_/CLK _1655_/D VGND VGND VPWR VPWR _1655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1440_ _1440_/A VGND VGND VPWR VPWR _1721_/D sky130_fd_sc_hd__clkbuf_1
X_1371_ _1756_/Q _1368_/X _1364_/X _1630_/Q _1361_/X VGND VGND VPWR VPWR _1371_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_15_0_CLK clkbuf_3_7_0_CLK/X VGND VGND VPWR VPWR _1762_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_31_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1707_ _1734_/CLK _1707_/D VGND VGND VPWR VPWR _1707_/Q sky130_fd_sc_hd__dfxtp_1
X_1638_ _1734_/CLK _1638_/D VGND VGND VPWR VPWR _1638_/Q sky130_fd_sc_hd__dfxtp_2
X_1569_ _1562_/X _1759_/Q _1569_/S VGND VGND VPWR VPWR _1569_/X sky130_fd_sc_hd__mux2_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_4_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_4_9_0_CLK/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0940_ _0966_/A VGND VGND VPWR VPWR _0940_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0871_ _1767_/Q _1738_/Q VGND VGND VPWR VPWR _1509_/B sky130_fd_sc_hd__and2_1
XFILLER_9_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1285_ _1767_/Q _1766_/Q _1749_/Q _1738_/Q VGND VGND VPWR VPWR _1285_/X sky130_fd_sc_hd__and4_1
X_1423_ _1423_/A VGND VGND VPWR VPWR _1712_/D sky130_fd_sc_hd__clkbuf_1
X_1354_ _1378_/A VGND VGND VPWR VPWR _1462_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1070_ _1621_/Q _1070_/B VGND VGND VPWR VPWR _1070_/Y sky130_fd_sc_hd__nand2_1
X_0854_ _0854_/A VGND VGND VPWR VPWR _0854_/X sky130_fd_sc_hd__clkbuf_1
X_0923_ _1674_/Q _0993_/C _0927_/B _1743_/Q _0966_/A VGND VGND VPWR VPWR _0923_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_45_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1337_ _1337_/A VGND VGND VPWR VPWR _1337_/Y sky130_fd_sc_hd__clkinv_2
X_1268_ _1268_/A VGND VGND VPWR VPWR _1671_/D sky130_fd_sc_hd__clkbuf_1
X_1406_ _1406_/A VGND VGND VPWR VPWR _1704_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1199_ input4/X _1170_/X _1171_/X _1652_/Q VGND VGND VPWR VPWR _1200_/B sky130_fd_sc_hd__a22o_1
XFILLER_3_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1122_ _1122_/A VGND VGND VPWR VPWR _1630_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1053_ _1556_/A VGND VGND VPWR VPWR _1402_/A sky130_fd_sc_hd__clkbuf_2
X_0837_ _0833_/X _0834_/X _0846_/C VGND VGND VPWR VPWR _0837_/X sky130_fd_sc_hd__o21a_1
X_0906_ _1353_/B _1353_/C _0906_/C VGND VGND VPWR VPWR _0916_/A sky130_fd_sc_hd__or3_1
XFILLER_24_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1740_ _1740_/CLK _1740_/D VGND VGND VPWR VPWR _1740_/Q sky130_fd_sc_hd__dfxtp_1
X_1671_ _1671_/CLK _1671_/D VGND VGND VPWR VPWR _1671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1105_ _1105_/A VGND VGND VPWR VPWR _1625_/D sky130_fd_sc_hd__clkbuf_1
X_1036_ input1/X VGND VGND VPWR VPWR _1375_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1654_ _1662_/CLK _1654_/D VGND VGND VPWR VPWR _1654_/Q sky130_fd_sc_hd__dfxtp_1
X_1723_ _1732_/CLK _1723_/D VGND VGND VPWR VPWR _1723_/Q sky130_fd_sc_hd__dfxtp_1
X_1585_ _1595_/A _1585_/B VGND VGND VPWR VPWR _1586_/S sky130_fd_sc_hd__nor2_1
X_1019_ _1442_/A VGND VGND VPWR VPWR _1029_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_5_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1370_ _1690_/Q _1367_/X _1369_/X VGND VGND VPWR VPWR _1690_/D sky130_fd_sc_hd__o21a_1
XFILLER_16_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1637_ _1732_/CLK _1637_/D VGND VGND VPWR VPWR _1637_/Q sky130_fd_sc_hd__dfxtp_1
X_1706_ _1765_/CLK _1706_/D VGND VGND VPWR VPWR _1706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1499_ _1509_/A _1748_/Q _1498_/Y VGND VGND VPWR VPWR _1499_/Y sky130_fd_sc_hd__a21oi_1
X_1568_ _1590_/A _1568_/B _1590_/C _1595_/A VGND VGND VPWR VPWR _1569_/S sky130_fd_sc_hd__or4_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0870_ _0865_/X _0867_/X _1580_/C VGND VGND VPWR VPWR _0870_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1422_ _1422_/A _1422_/B VGND VGND VPWR VPWR _1423_/A sky130_fd_sc_hd__or2_1
X_1284_ _1286_/A _1286_/B _1286_/C VGND VGND VPWR VPWR _1284_/X sky130_fd_sc_hd__or3_1
X_1353_ _1353_/A _1353_/B _1353_/C _1353_/D VGND VGND VPWR VPWR _1378_/A sky130_fd_sc_hd__or4_4
X_0999_ _1717_/Q _1433_/A _1005_/C VGND VGND VPWR VPWR _1000_/A sky130_fd_sc_hd__and3_1
XFILLER_46_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_14_0_CLK clkbuf_3_7_0_CLK/X VGND VGND VPWR VPWR _1765_/CLK sky130_fd_sc_hd__clkbuf_2
X_0853_ _0851_/X _0853_/B VGND VGND VPWR VPWR _0854_/A sky130_fd_sc_hd__and2b_1
X_0922_ _1347_/D VGND VGND VPWR VPWR _0966_/A sky130_fd_sc_hd__clkbuf_2
X_1405_ _1405_/A _1422_/B VGND VGND VPWR VPWR _1406_/A sky130_fd_sc_hd__or2_1
X_1336_ _1323_/A _1339_/A _1334_/Y _1335_/Y VGND VGND VPWR VPWR _1682_/D sky130_fd_sc_hd__a31oi_1
XFILLER_28_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput1 RST_N VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_4
X_1267_ _1267_/A _1267_/B VGND VGND VPWR VPWR _1268_/A sky130_fd_sc_hd__or2_1
X_1198_ _1198_/A VGND VGND VPWR VPWR _1651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_4_7_0_CLK/A sky130_fd_sc_hd__clkbuf_2
X_1121_ _1144_/A _1121_/B VGND VGND VPWR VPWR _1122_/A sky130_fd_sc_hd__and2_1
X_1052_ input1/X VGND VGND VPWR VPWR _1556_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0836_ _0833_/X _0834_/X _0835_/X _1676_/Q VGND VGND VPWR VPWR _0846_/C sky130_fd_sc_hd__a22o_1
X_0905_ _1643_/Q _0789_/C VGND VGND VPWR VPWR _0906_/C sky130_fd_sc_hd__or2b_1
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1319_ _1319_/A VGND VGND VPWR VPWR _1319_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1670_ _1671_/CLK _1670_/D VGND VGND VPWR VPWR _1670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1104_ _1504_/A _1104_/B VGND VGND VPWR VPWR _1105_/A sky130_fd_sc_hd__or2_1
X_1035_ _1035_/A VGND VGND VPWR VPWR _1035_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0819_ _1741_/Q VGND VGND VPWR VPWR _0946_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1584_ _1584_/A VGND VGND VPWR VPWR _1761_/D sky130_fd_sc_hd__clkbuf_1
X_1722_ _1732_/CLK _1722_/D VGND VGND VPWR VPWR _1722_/Q sky130_fd_sc_hd__dfxtp_1
X_1653_ _1662_/CLK _1653_/D VGND VGND VPWR VPWR _1653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1018_ _1018_/A VGND VGND VPWR VPWR _1018_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1705_ _1734_/CLK _1705_/D VGND VGND VPWR VPWR _1705_/Q sky130_fd_sc_hd__dfxtp_1
X_1567_ _1567_/A VGND VGND VPWR VPWR _1758_/D sky130_fd_sc_hd__clkbuf_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1636_ _1732_/CLK _1636_/D VGND VGND VPWR VPWR _1636_/Q sky130_fd_sc_hd__dfxtp_1
X_1498_ _1498_/A _1498_/B VGND VGND VPWR VPWR _1498_/Y sky130_fd_sc_hd__nand2_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1421_ _1421_/A _1421_/B VGND VGND VPWR VPWR _1711_/D sky130_fd_sc_hd__nor2_1
X_1283_ _1684_/Q _1681_/Q _1677_/Q _1676_/Q VGND VGND VPWR VPWR _1286_/C sky130_fd_sc_hd__or4_1
X_1352_ _1382_/A VGND VGND VPWR VPWR _1352_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0998_ _1442_/A VGND VGND VPWR VPWR _1433_/A sky130_fd_sc_hd__clkbuf_1
X_1619_ _1650_/CLK _1619_/D VGND VGND VPWR VPWR _1619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0921_ _0921_/A _1040_/B VGND VGND VPWR VPWR _0927_/B sky130_fd_sc_hd__nor2_1
X_0852_ _0806_/X _0847_/Y _0848_/X _1675_/Q VGND VGND VPWR VPWR _0853_/B sky130_fd_sc_hd__a31o_1
X_1335_ _1682_/Q _1323_/A _1107_/A VGND VGND VPWR VPWR _1335_/Y sky130_fd_sc_hd__o21ai_1
X_1404_ _1429_/B VGND VGND VPWR VPWR _1422_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 slave_adr_i[0] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
X_1197_ _1197_/A _1197_/B VGND VGND VPWR VPWR _1198_/A sky130_fd_sc_hd__or2_1
X_1266_ input25/X _1195_/A _1102_/A _1671_/Q VGND VGND VPWR VPWR _1267_/B sky130_fd_sc_hd__o22a_1
XFILLER_10_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1051_ _1051_/A VGND VGND VPWR VPWR _1613_/D sky130_fd_sc_hd__clkbuf_1
X_1120_ input47/X _1092_/X _1094_/X _1630_/Q VGND VGND VPWR VPWR _1121_/B sky130_fd_sc_hd__a22o_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0904_ _1644_/Q VGND VGND VPWR VPWR _0921_/A sky130_fd_sc_hd__inv_2
X_0835_ _0951_/A _0946_/A _0942_/A VGND VGND VPWR VPWR _0835_/X sky130_fd_sc_hd__or3_1
X_1318_ _0830_/A _1294_/X _1317_/X _1279_/X VGND VGND VPWR VPWR _1679_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_4_13_0_CLK clkbuf_3_6_0_CLK/X VGND VGND VPWR VPWR _1752_/CLK sky130_fd_sc_hd__clkbuf_2
X_1249_ _1249_/A VGND VGND VPWR VPWR _1665_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_40 _1411_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1034_ _1732_/Q _1439_/B _1034_/C VGND VGND VPWR VPWR _1035_/A sky130_fd_sc_hd__and3_1
X_1103_ input42/X _1074_/X _1102_/X _1625_/Q VGND VGND VPWR VPWR _1104_/B sky130_fd_sc_hd__o22a_1
Xclkbuf_3_2_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_4_5_0_CLK/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0818_ _1741_/Q _0828_/A _0951_/A VGND VGND VPWR VPWR _1331_/A sky130_fd_sc_hd__nand3b_2
XFILLER_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1721_ _1732_/CLK _1721_/D VGND VGND VPWR VPWR _1721_/Q sky130_fd_sc_hd__dfxtp_1
X_1583_ _1583_/A _1583_/B VGND VGND VPWR VPWR _1584_/A sky130_fd_sc_hd__and2_1
X_1652_ _1662_/CLK _1652_/D VGND VGND VPWR VPWR _1652_/Q sky130_fd_sc_hd__dfxtp_1
X_1017_ _1725_/Q _1017_/B _1017_/C VGND VGND VPWR VPWR _1018_/A sky130_fd_sc_hd__and3_1
XFILLER_43_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1704_ _1734_/CLK _1704_/D VGND VGND VPWR VPWR _1704_/Q sky130_fd_sc_hd__dfxtp_1
X_1497_ _1498_/A _1488_/X _1491_/X _1496_/Y _1305_/A VGND VGND VPWR VPWR _1747_/D
+ sky130_fd_sc_hd__a311oi_1
X_1566_ _1583_/A _1566_/B VGND VGND VPWR VPWR _1567_/A sky130_fd_sc_hd__and2_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1635_ _1717_/CLK _1635_/D VGND VGND VPWR VPWR _1635_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1420_ _1420_/A VGND VGND VPWR VPWR _1710_/D sky130_fd_sc_hd__clkbuf_1
X_1351_ _1381_/A VGND VGND VPWR VPWR _1351_/X sky130_fd_sc_hd__clkbuf_2
X_1282_ _1683_/Q _1682_/Q VGND VGND VPWR VPWR _1286_/B sky130_fd_sc_hd__or2_1
X_1618_ _1742_/CLK _1618_/D VGND VGND VPWR VPWR _1618_/Q sky130_fd_sc_hd__dfxtp_1
X_0997_ _0997_/A VGND VGND VPWR VPWR _1442_/A sky130_fd_sc_hd__buf_2
X_1549_ _1549_/A VGND VGND VPWR VPWR _1755_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0920_ _0989_/C VGND VGND VPWR VPWR _0993_/C sky130_fd_sc_hd__clkbuf_1
X_0851_ _0806_/X _1675_/Q _0847_/Y _0848_/X _1462_/A VGND VGND VPWR VPWR _0851_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1334_ _1333_/A _1333_/B _1333_/C VGND VGND VPWR VPWR _1334_/Y sky130_fd_sc_hd__o21ai_1
X_1265_ _1265_/A VGND VGND VPWR VPWR _1670_/D sky130_fd_sc_hd__clkbuf_1
X_1403_ _1403_/A VGND VGND VPWR VPWR _1703_/D sky130_fd_sc_hd__clkbuf_1
Xinput3 slave_adr_i[10] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1196_ input3/X _1195_/X _1175_/X _1651_/Q VGND VGND VPWR VPWR _1197_/B sky130_fd_sc_hd__o22a_1
XFILLER_27_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1050_ _1613_/Q _1063_/B VGND VGND VPWR VPWR _1051_/A sky130_fd_sc_hd__or2_1
XFILLER_18_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0834_ _0951_/A _0946_/A _0942_/A VGND VGND VPWR VPWR _0834_/X sky130_fd_sc_hd__or3b_1
X_0903_ _1086_/A _1622_/Q _1462_/A VGND VGND VPWR VPWR _0903_/Y sky130_fd_sc_hd__a21oi_2
X_1317_ _1317_/A _1317_/B _1316_/Y VGND VGND VPWR VPWR _1317_/X sky130_fd_sc_hd__or3b_1
X_1248_ _1267_/A _1248_/B VGND VGND VPWR VPWR _1249_/A sky130_fd_sc_hd__or2_1
X_1179_ input29/X _1170_/X _1171_/X _1646_/Q VGND VGND VPWR VPWR _1180_/B sky130_fd_sc_hd__a22o_1
XFILLER_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_30 slave_dat_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 slave_adr_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1102_ _1102_/A VGND VGND VPWR VPWR _1102_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1033_ _1033_/A VGND VGND VPWR VPWR _1033_/X sky130_fd_sc_hd__clkbuf_1
Xinput50 slave_dat_i[9] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_1
X_0817_ _0826_/A VGND VGND VPWR VPWR _0951_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1720_ _1732_/CLK _1720_/D VGND VGND VPWR VPWR _1720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1651_ _1662_/CLK _1651_/D VGND VGND VPWR VPWR _1651_/Q sky130_fd_sc_hd__dfxtp_1
X_1582_ _1761_/Q _1573_/X _1581_/X _1576_/X VGND VGND VPWR VPWR _1583_/B sky130_fd_sc_hd__a22o_1
Xclkbuf_4_12_0_CLK clkbuf_3_6_0_CLK/X VGND VGND VPWR VPWR _1712_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1016_ _1016_/A VGND VGND VPWR VPWR _1016_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_4_3_0_CLK/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1634_ _1730_/CLK _1634_/D VGND VGND VPWR VPWR _1634_/Q sky130_fd_sc_hd__dfxtp_1
X_1703_ _1734_/CLK _1703_/D VGND VGND VPWR VPWR _1703_/Q sky130_fd_sc_hd__dfxtp_1
X_1496_ _1498_/B _1488_/X _1498_/A VGND VGND VPWR VPWR _1496_/Y sky130_fd_sc_hd__a21oi_1
X_1565_ _1758_/Q _1542_/X _1564_/X _1546_/X VGND VGND VPWR VPWR _1566_/B sky130_fd_sc_hd__a22o_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1281_ _1680_/Q _1679_/Q _1678_/Q VGND VGND VPWR VPWR _1286_/A sky130_fd_sc_hd__or3_1
X_1350_ _1346_/Y _1347_/X _1382_/A VGND VGND VPWR VPWR _1381_/A sky130_fd_sc_hd__o21ai_4
X_0996_ _0996_/A VGND VGND VPWR VPWR _0996_/X sky130_fd_sc_hd__clkbuf_1
X_1617_ _1742_/CLK _1617_/D VGND VGND VPWR VPWR _1617_/Q sky130_fd_sc_hd__dfxtp_1
X_1548_ _1554_/A _1548_/B VGND VGND VPWR VPWR _1549_/A sky130_fd_sc_hd__and2_1
XFILLER_39_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1479_ _1479_/A VGND VGND VPWR VPWR _1606_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_24_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0850_ _1289_/B VGND VGND VPWR VPWR _1462_/A sky130_fd_sc_hd__clkbuf_2
X_1402_ _1402_/A _1427_/B _1402_/C VGND VGND VPWR VPWR _1403_/A sky130_fd_sc_hd__and3_1
Xinput4 slave_adr_i[11] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
X_1333_ _1333_/A _1333_/B _1333_/C VGND VGND VPWR VPWR _1339_/A sky130_fd_sc_hd__or3_2
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1264_ _1521_/A _1264_/B VGND VGND VPWR VPWR _1265_/A sky130_fd_sc_hd__and2_1
X_1195_ _1195_/A VGND VGND VPWR VPWR _1195_/X sky130_fd_sc_hd__clkbuf_2
X_0979_ _1712_/Q _0940_/X _0934_/X _1696_/Q _0978_/X VGND VGND VPWR VPWR _1422_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_19_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0833_ _1677_/Q VGND VGND VPWR VPWR _0833_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0902_ _1623_/Q VGND VGND VPWR VPWR _1086_/A sky130_fd_sc_hd__inv_2
X_1316_ _1321_/A _1321_/B VGND VGND VPWR VPWR _1316_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1247_ input18/X _1231_/X _1102_/A _1665_/Q VGND VGND VPWR VPWR _1248_/B sky130_fd_sc_hd__o22a_1
X_1178_ _1178_/A VGND VGND VPWR VPWR _1645_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_31 slave_dat_i[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_20 slave_adr_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1032_ _1731_/Q _1439_/B _1034_/C VGND VGND VPWR VPWR _1033_/A sky130_fd_sc_hd__and3_1
X_1101_ _1211_/A VGND VGND VPWR VPWR _1102_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput40 slave_dat_i[14] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_1
Xinput51 slave_stb_i VGND VGND VPWR VPWR _1071_/B sky130_fd_sc_hd__clkbuf_1
X_0816_ _0808_/X _1342_/A _1337_/A _1682_/Q VGND VGND VPWR VPWR _0824_/A sky130_fd_sc_hd__o22a_1
XFILLER_29_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1581_ _1562_/X _1761_/Q _1581_/S VGND VGND VPWR VPWR _1581_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1650_ _1650_/CLK _1650_/D VGND VGND VPWR VPWR _1650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1015_ _1724_/Q _1017_/B _1017_/C VGND VGND VPWR VPWR _1016_/A sky130_fd_sc_hd__and3_1
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1564_ _1562_/X _1758_/Q _1564_/S VGND VGND VPWR VPWR _1564_/X sky130_fd_sc_hd__mux2_1
X_1633_ _1717_/CLK _1633_/D VGND VGND VPWR VPWR _1633_/Q sky130_fd_sc_hd__dfxtp_1
X_1702_ _1733_/CLK _1702_/D VGND VGND VPWR VPWR _1702_/Q sky130_fd_sc_hd__dfxtp_1
X_1495_ _1488_/X _1493_/Y _1494_/X _1305_/A VGND VGND VPWR VPWR _1746_/D sky130_fd_sc_hd__a211o_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_11_0_CLK clkbuf_3_5_0_CLK/X VGND VGND VPWR VPWR _1730_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_48_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1280_ _1675_/Q _1080_/X _1277_/X _1279_/X VGND VGND VPWR VPWR _1675_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0995_ _0995_/A _1429_/A VGND VGND VPWR VPWR _0996_/A sky130_fd_sc_hd__and2_1
X_1547_ _1755_/Q _1542_/X _1545_/X _1546_/X VGND VGND VPWR VPWR _1548_/B sky130_fd_sc_hd__a22o_1
X_1616_ _1742_/CLK _1616_/D VGND VGND VPWR VPWR _1616_/Q sky130_fd_sc_hd__dfxtp_1
X_1478_ _1629_/Q _1086_/B _1477_/Y _1469_/X VGND VGND VPWR VPWR _1742_/D sky130_fd_sc_hd__o211a_1
XFILLER_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_0_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_4_1_0_CLK/A sky130_fd_sc_hd__clkbuf_2
X_1401_ _1401_/A VGND VGND VPWR VPWR _1702_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput5 slave_adr_i[12] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
X_1332_ _1682_/Q _1331_/Y _1486_/A VGND VGND VPWR VPWR _1333_/C sky130_fd_sc_hd__mux2_1
XFILLER_36_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1263_ input23/X _1242_/X _1243_/X _1670_/Q VGND VGND VPWR VPWR _1264_/B sky130_fd_sc_hd__a22o_1
X_1194_ _1194_/A VGND VGND VPWR VPWR _1650_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0978_ _1736_/Q _0993_/B _0993_/C VGND VGND VPWR VPWR _0978_/X sky130_fd_sc_hd__and3_1
XFILLER_10_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0832_ _0825_/X _1313_/A _0830_/Y _0831_/X VGND VGND VPWR VPWR _0846_/B sky130_fd_sc_hd__a211o_1
X_0901_ _0901_/A VGND VGND VPWR VPWR _0901_/X sky130_fd_sc_hd__clkbuf_1
X_1315_ _1321_/A _1321_/B VGND VGND VPWR VPWR _1317_/B sky130_fd_sc_hd__nor2_1
XFILLER_2_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1246_ _1246_/A VGND VGND VPWR VPWR _1664_/D sky130_fd_sc_hd__clkbuf_1
X_1177_ _1197_/A _1177_/B VGND VGND VPWR VPWR _1178_/A sky130_fd_sc_hd__or2_1
XANTENNA_32 slave_dat_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 slave_cyc_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 slave_adr_i[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1031_ _1442_/A VGND VGND VPWR VPWR _1439_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1100_ _1347_/D _1231_/A VGND VGND VPWR VPWR _1211_/A sky130_fd_sc_hd__nand2_2
XFILLER_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput41 slave_dat_i[15] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_1
Xinput30 slave_adr_i[6] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_1
X_0815_ _0828_/A _1741_/Q _0826_/A VGND VGND VPWR VPWR _1337_/A sky130_fd_sc_hd__nand3b_2
Xinput52 slave_we_i VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__clkbuf_2
X_1229_ _1251_/A _1229_/B VGND VGND VPWR VPWR _1230_/A sky130_fd_sc_hd__and2_1
XFILLER_32_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1580_ _1590_/A _1580_/B _1580_/C _1600_/D VGND VGND VPWR VPWR _1581_/S sky130_fd_sc_hd__or4_1
XFILLER_7_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1014_ _1014_/A VGND VGND VPWR VPWR _1014_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1701_ _1733_/CLK _1701_/D VGND VGND VPWR VPWR _1701_/Q sky130_fd_sc_hd__dfxtp_1
X_1494_ _1746_/Q _1504_/B _1606_/B VGND VGND VPWR VPWR _1494_/X sky130_fd_sc_hd__and3_1
X_1563_ _1563_/A _1600_/D _1563_/C _1563_/D VGND VGND VPWR VPWR _1564_/S sky130_fd_sc_hd__or4_1
X_1632_ _1717_/CLK _1632_/D VGND VGND VPWR VPWR _1632_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0994_ _1716_/Q _0997_/A _0934_/X _1700_/Q _0993_/X VGND VGND VPWR VPWR _1429_/A
+ sky130_fd_sc_hd__a221o_1
X_1546_ _1576_/A VGND VGND VPWR VPWR _1546_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1477_ _1477_/A _1477_/B VGND VGND VPWR VPWR _1477_/Y sky130_fd_sc_hd__nand2_1
X_1615_ _1742_/CLK _1615_/D VGND VGND VPWR VPWR _1615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1331_ _1331_/A VGND VGND VPWR VPWR _1331_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1400_ _1400_/A _1459_/B VGND VGND VPWR VPWR _1401_/A sky130_fd_sc_hd__or2_1
Xinput6 slave_adr_i[13] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1193_ _1216_/A _1193_/B VGND VGND VPWR VPWR _1194_/A sky130_fd_sc_hd__and2_1
X_1262_ _1262_/A VGND VGND VPWR VPWR _1669_/D sky130_fd_sc_hd__clkbuf_1
X_0977_ _0977_/A VGND VGND VPWR VPWR _0977_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1529_ _1554_/A _1529_/B VGND VGND VPWR VPWR _1530_/A sky130_fd_sc_hd__and2_1
Xclkbuf_4_10_0_CLK clkbuf_3_5_0_CLK/X VGND VGND VPWR VPWR _1732_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_19_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ _0900_/A _0900_/B _0900_/C VGND VGND VPWR VPWR _0901_/A sky130_fd_sc_hd__and3_1
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0831_ _0825_/X _1313_/A _1319_/A _0830_/A VGND VGND VPWR VPWR _0831_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1314_ _0830_/A _1313_/Y _1314_/S VGND VGND VPWR VPWR _1321_/B sky130_fd_sc_hd__mux2_1
X_1245_ _1251_/A _1245_/B VGND VGND VPWR VPWR _1246_/A sky130_fd_sc_hd__and2_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1176_ input28/X _1159_/X _1175_/X _1645_/Q VGND VGND VPWR VPWR _1177_/B sky130_fd_sc_hd__o22a_1
XFILLER_24_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_33 slave_dat_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 slave_dat_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_11 slave_adr_i[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1030_ _1030_/A VGND VGND VPWR VPWR _1030_/X sky130_fd_sc_hd__clkbuf_1
Xinput31 slave_adr_i[7] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_1
Xinput20 slave_adr_i[26] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__clkbuf_1
X_0814_ _1742_/Q VGND VGND VPWR VPWR _0826_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput42 slave_dat_i[1] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_1
Xinput53 spiMaster_miso VGND VGND VPWR VPWR _1562_/A sky130_fd_sc_hd__clkbuf_2
X_1228_ input12/X _1206_/X _1207_/X _1660_/Q VGND VGND VPWR VPWR _1229_/B sky130_fd_sc_hd__a22o_1
X_1159_ _1195_/A VGND VGND VPWR VPWR _1159_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1013_ _1723_/Q _1017_/B _1017_/C VGND VGND VPWR VPWR _1014_/A sky130_fd_sc_hd__and3_1
XFILLER_27_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1631_ _1717_/CLK _1631_/D VGND VGND VPWR VPWR _1631_/Q sky130_fd_sc_hd__dfxtp_2
X_1700_ _1730_/CLK _1700_/D VGND VGND VPWR VPWR _1700_/Q sky130_fd_sc_hd__dfxtp_1
X_1493_ _1491_/X _1492_/Y _1342_/B VGND VGND VPWR VPWR _1493_/Y sky130_fd_sc_hd__o21ai_1
X_1562_ _1562_/A VGND VGND VPWR VPWR _1562_/X sky130_fd_sc_hd__clkbuf_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0993_ _1622_/Q _0993_/B _0993_/C VGND VGND VPWR VPWR _0993_/X sky130_fd_sc_hd__and3_1
X_1614_ _1742_/CLK _1614_/D VGND VGND VPWR VPWR _1614_/Q sky130_fd_sc_hd__dfxtp_1
X_1545_ _1508_/X _1755_/Q _1545_/S VGND VGND VPWR VPWR _1545_/X sky130_fd_sc_hd__mux2_1
X_1476_ _1628_/Q _1086_/B _1475_/Y _1469_/X VGND VGND VPWR VPWR _1741_/D sky130_fd_sc_hd__o211a_1
XFILLER_40_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1330_ _1681_/Q _1294_/X _1327_/Y _1328_/X _1329_/X VGND VGND VPWR VPWR _1681_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_5_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1261_ _1267_/A _1261_/B VGND VGND VPWR VPWR _1262_/A sky130_fd_sc_hd__or2_1
Xinput7 slave_adr_i[14] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1192_ input33/X _1170_/X _1171_/X _1650_/Q VGND VGND VPWR VPWR _1193_/B sky130_fd_sc_hd__a22o_1
X_0976_ _1421_/A _0995_/A VGND VGND VPWR VPWR _0977_/A sky130_fd_sc_hd__and2b_1
X_1528_ _1752_/Q _1507_/X _1527_/X _1514_/X VGND VGND VPWR VPWR _1529_/B sky130_fd_sc_hd__a22o_1
X_1459_ _1459_/A _1459_/B VGND VGND VPWR VPWR _1733_/D sky130_fd_sc_hd__nor2_1
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0830_ _0830_/A _1319_/A VGND VGND VPWR VPWR _0830_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1313_ _1313_/A VGND VGND VPWR VPWR _1313_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1244_ input17/X _1242_/X _1243_/X _1664_/Q VGND VGND VPWR VPWR _1245_/B sky130_fd_sc_hd__a22o_1
X_1175_ _1211_/A VGND VGND VPWR VPWR _1175_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_23 slave_dat_i[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 slave_dat_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_12 slave_adr_i[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0959_ _0980_/A _1413_/A VGND VGND VPWR VPWR _0960_/A sky130_fd_sc_hd__and2_1
XFILLER_47_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput21 slave_adr_i[27] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_1
Xinput43 slave_dat_i[2] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_1
Xinput32 slave_adr_i[8] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__clkbuf_1
X_0813_ _1740_/Q VGND VGND VPWR VPWR _0828_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput10 slave_adr_i[17] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_1
X_1227_ _1227_/A VGND VGND VPWR VPWR _1659_/D sky130_fd_sc_hd__clkbuf_1
X_1158_ _1158_/A VGND VGND VPWR VPWR _1640_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1089_ _1606_/A VGND VGND VPWR VPWR _1107_/A sky130_fd_sc_hd__buf_2
XFILLER_20_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1012_ _1012_/A VGND VGND VPWR VPWR _1012_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1630_ _1717_/CLK _1630_/D VGND VGND VPWR VPWR _1630_/Q sky130_fd_sc_hd__dfxtp_1
X_1492_ _1746_/Q _1745_/Q VGND VGND VPWR VPWR _1492_/Y sky130_fd_sc_hd__nor2_1
X_1561_ _1561_/A VGND VGND VPWR VPWR _1757_/D sky130_fd_sc_hd__clkbuf_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1759_ _1762_/CLK _1759_/D VGND VGND VPWR VPWR _1759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0992_ _0992_/A VGND VGND VPWR VPWR _0992_/X sky130_fd_sc_hd__clkbuf_1
X_1544_ _1590_/A _1590_/B _1590_/C _1557_/D VGND VGND VPWR VPWR _1545_/S sky130_fd_sc_hd__or4_1
X_1613_ _1742_/CLK _1613_/D VGND VGND VPWR VPWR _1613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1475_ _1475_/A _1477_/B VGND VGND VPWR VPWR _1475_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 slave_adr_i[15] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1260_ input22/X _1231_/X _1102_/A _1669_/Q VGND VGND VPWR VPWR _1261_/B sky130_fd_sc_hd__o22a_1
X_1191_ _1191_/A VGND VGND VPWR VPWR _1649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0975_ _1711_/Q _1069_/A _0967_/X _1695_/Q VGND VGND VPWR VPWR _1421_/A sky130_fd_sc_hd__a22oi_4
X_1527_ _1752_/Q _1524_/X _1527_/S VGND VGND VPWR VPWR _1527_/X sky130_fd_sc_hd__mux2_1
X_1458_ _1732_/Q _1070_/B _1421_/B VGND VGND VPWR VPWR _1732_/D sky130_fd_sc_hd__a21o_1
XFILLER_19_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1389_ _1763_/Q _1382_/X _1378_/X _1637_/Q _1048_/A VGND VGND VPWR VPWR _1389_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_35_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1312_ _1321_/A _1309_/Y _1311_/Y VGND VGND VPWR VPWR _1678_/D sky130_fd_sc_hd__a21oi_1
X_1243_ _1243_/A VGND VGND VPWR VPWR _1243_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1174_ _1174_/A VGND VGND VPWR VPWR _1644_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_13 slave_adr_i[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_24 slave_dat_i[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 slave_dat_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0889_ _1692_/Q _1691_/Q _1531_/A VGND VGND VPWR VPWR _0889_/X sky130_fd_sc_hd__mux2_1
X_0958_ _1707_/Q _1272_/B _0956_/X _0957_/X VGND VGND VPWR VPWR _1413_/A sky130_fd_sc_hd__o22a_1
XFILLER_46_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput44 slave_dat_i[3] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_1
Xinput33 slave_adr_i[9] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_1
X_0812_ _1477_/A _0838_/A _1473_/A VGND VGND VPWR VPWR _1342_/A sky130_fd_sc_hd__or3_2
Xinput11 slave_adr_i[18] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__clkbuf_1
Xinput22 slave_adr_i[28] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1226_ _1233_/A _1226_/B VGND VGND VPWR VPWR _1227_/A sky130_fd_sc_hd__or2_1
X_1157_ _1180_/A _1157_/B VGND VGND VPWR VPWR _1158_/A sky130_fd_sc_hd__and2_1
XFILLER_32_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1088_ input1/X VGND VGND VPWR VPWR _1606_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1011_ _1722_/Q _1017_/B _1017_/C VGND VGND VPWR VPWR _1012_/A sky130_fd_sc_hd__and3_1
XFILLER_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1209_ _1216_/A _1209_/B VGND VGND VPWR VPWR _1210_/A sky130_fd_sc_hd__and2_1
XFILLER_40_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1560_ _1583_/A _1560_/B VGND VGND VPWR VPWR _1561_/A sky130_fd_sc_hd__and2_1
XFILLER_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1491_ _1491_/A _1498_/B VGND VGND VPWR VPWR _1491_/X sky130_fd_sc_hd__or2_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1758_ _1762_/CLK _1758_/D VGND VGND VPWR VPWR _1758_/Q sky130_fd_sc_hd__dfxtp_1
X_1689_ _1712_/CLK _1689_/D VGND VGND VPWR VPWR _1689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0991_ _0995_/A _1427_/C VGND VGND VPWR VPWR _0992_/A sky130_fd_sc_hd__and2_1
X_1543_ _1600_/A VGND VGND VPWR VPWR _1590_/A sky130_fd_sc_hd__clkbuf_1
X_1474_ _1627_/Q _1086_/B _1473_/Y _1469_/X VGND VGND VPWR VPWR _1740_/D sky130_fd_sc_hd__o211a_1
X_1612_ _1742_/CLK _1612_/D VGND VGND VPWR VPWR _1612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 slave_adr_i[16] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
X_1190_ _1197_/A _1190_/B VGND VGND VPWR VPWR _1191_/A sky130_fd_sc_hd__or2_1
XFILLER_44_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0974_ _0974_/A VGND VGND VPWR VPWR _0974_/X sky130_fd_sc_hd__clkbuf_1
X_1526_ _1551_/A _1574_/B VGND VGND VPWR VPWR _1527_/S sky130_fd_sc_hd__nor2_1
X_1457_ _1457_/A VGND VGND VPWR VPWR _1731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1388_ _1697_/Q _1381_/X _1387_/X VGND VGND VPWR VPWR _1697_/D sky130_fd_sc_hd__o21a_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1311_ _0825_/X _1323_/A _1107_/A VGND VGND VPWR VPWR _1311_/Y sky130_fd_sc_hd__o21ai_1
X_1242_ _1242_/A VGND VGND VPWR VPWR _1242_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1173_ _1180_/A _1173_/B VGND VGND VPWR VPWR _1174_/A sky130_fd_sc_hd__and2_1
XANTENNA_36 slave_dat_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 slave_dat_i[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_14 slave_adr_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0957_ _1767_/Q _1079_/C _0927_/B _1744_/Q _0966_/A VGND VGND VPWR VPWR _0957_/X
+ sky130_fd_sc_hd__a221o_1
X_0888_ _1690_/Q _1689_/Q _1531_/A VGND VGND VPWR VPWR _0888_/X sky130_fd_sc_hd__mux2_1
X_1509_ _1509_/A _1509_/B _1509_/C VGND VGND VPWR VPWR _1563_/A sky130_fd_sc_hd__and3_1
XFILLER_15_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput45 slave_dat_i[4] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__clkbuf_1
Xinput34 slave_cyc_i VGND VGND VPWR VPWR _1071_/C sky130_fd_sc_hd__clkbuf_1
Xinput23 slave_adr_i[29] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_1
X_0811_ _1740_/Q VGND VGND VPWR VPWR _1473_/A sky130_fd_sc_hd__inv_2
Xinput12 slave_adr_i[19] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1087_ _1638_/Q _1086_/B _1086_/Y _1083_/X VGND VGND VPWR VPWR _1623_/D sky130_fd_sc_hd__o211a_1
X_1225_ input11/X _1195_/X _1211_/X _1659_/Q VGND VGND VPWR VPWR _1226_/B sky130_fd_sc_hd__o22a_1
X_1156_ input52/X _1134_/X _1135_/X _1346_/A VGND VGND VPWR VPWR _1157_/B sky130_fd_sc_hd__a22o_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1010_ _1010_/A VGND VGND VPWR VPWR _1010_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1208_ input6/X _1206_/X _1207_/X _1654_/Q VGND VGND VPWR VPWR _1209_/B sky130_fd_sc_hd__a22o_1
X_1139_ _1211_/A VGND VGND VPWR VPWR _1139_/X sky130_fd_sc_hd__buf_2
XFILLER_16_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1490_ _1745_/Q _1488_/X _1489_/Y _1329_/X VGND VGND VPWR VPWR _1745_/D sky130_fd_sc_hd__o211a_1
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1757_ _1762_/CLK _1757_/D VGND VGND VPWR VPWR _1757_/Q sky130_fd_sc_hd__dfxtp_1
X_1688_ _1712_/CLK _1688_/D VGND VGND VPWR VPWR _1688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1611_ _1742_/CLK _1611_/D VGND VGND VPWR VPWR _1611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0990_ _1715_/Q _0997_/A _0967_/A _1699_/Q _0989_/X VGND VGND VPWR VPWR _1427_/C
+ sky130_fd_sc_hd__a221o_1
X_1542_ _1573_/A VGND VGND VPWR VPWR _1542_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1473_ _1473_/A _1477_/B VGND VGND VPWR VPWR _1473_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0973_ _0980_/A _1419_/A VGND VGND VPWR VPWR _0974_/A sky130_fd_sc_hd__and2_1
X_1525_ _1550_/A _1580_/B _1550_/C VGND VGND VPWR VPWR _1574_/B sky130_fd_sc_hd__or3_1
X_1456_ _1731_/Q _1456_/B _1456_/C VGND VGND VPWR VPWR _1457_/A sky130_fd_sc_hd__and3_1
X_1387_ _1762_/Q _1382_/X _1378_/X _1636_/Q _1375_/X VGND VGND VPWR VPWR _1387_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_35_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1310_ _1310_/A VGND VGND VPWR VPWR _1323_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1241_ _1241_/A VGND VGND VPWR VPWR _1663_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1172_ input27/X _1170_/X _1171_/X _1644_/Q VGND VGND VPWR VPWR _1173_/B sky130_fd_sc_hd__a22o_1
XFILLER_24_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_26 slave_dat_i[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 slave_dat_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_15 slave_adr_i[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0956_ _1691_/Q _0961_/B VGND VGND VPWR VPWR _0956_/X sky130_fd_sc_hd__and2_1
X_0887_ _1568_/B _0870_/X _1595_/A _0886_/X VGND VGND VPWR VPWR _0900_/B sky130_fd_sc_hd__a211o_1
X_1508_ _1562_/A VGND VGND VPWR VPWR _1508_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1439_ _1721_/Q _1439_/B _1439_/C VGND VGND VPWR VPWR _1440_/A sky130_fd_sc_hd__and3_1
XFILLER_23_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput13 slave_adr_i[1] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_1
X_0810_ _1741_/Q VGND VGND VPWR VPWR _0838_/A sky130_fd_sc_hd__inv_2
XFILLER_14_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput46 slave_dat_i[5] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__clkbuf_1
Xinput35 slave_dat_i[0] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_1
Xinput24 slave_adr_i[2] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1224_ _1224_/A VGND VGND VPWR VPWR _1658_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1086_ _1086_/A _1086_/B VGND VGND VPWR VPWR _1086_/Y sky130_fd_sc_hd__nand2_1
X_1155_ _1155_/A VGND VGND VPWR VPWR _1639_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0939_ _0939_/A VGND VGND VPWR VPWR _0939_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1207_ _1243_/A VGND VGND VPWR VPWR _1207_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1069_ _1069_/A VGND VGND VPWR VPWR _1070_/B sky130_fd_sc_hd__buf_2
X_1138_ _1138_/A VGND VGND VPWR VPWR _1634_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1756_ _1762_/CLK _1756_/D VGND VGND VPWR VPWR _1756_/Q sky130_fd_sc_hd__dfxtp_1
X_1687_ _1752_/CLK _1687_/D VGND VGND VPWR VPWR _1687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1610_ _1742_/CLK _1610_/D VGND VGND VPWR VPWR _1610_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1541_ _1541_/A VGND VGND VPWR VPWR _1754_/D sky130_fd_sc_hd__clkbuf_1
X_1472_ _0806_/X _1462_/A _1471_/Y _1469_/X VGND VGND VPWR VPWR _1739_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1739_ _1767_/CLK _1739_/D VGND VGND VPWR VPWR _1739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0972_ _1710_/Q _0940_/X _0967_/X _1694_/Q VGND VGND VPWR VPWR _1419_/A sky130_fd_sc_hd__a22o_1
X_1524_ _1562_/A VGND VGND VPWR VPWR _1524_/X sky130_fd_sc_hd__clkbuf_2
X_1455_ _1730_/Q _1070_/B _1421_/B VGND VGND VPWR VPWR _1730_/D sky130_fd_sc_hd__a21o_1
X_1386_ _1696_/Q _1381_/X _1385_/X VGND VGND VPWR VPWR _1696_/D sky130_fd_sc_hd__o21a_1
XFILLER_18_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_CLK CLK VGND VGND VPWR VPWR clkbuf_0_CLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1240_ _1267_/A _1240_/B VGND VGND VPWR VPWR _1241_/A sky130_fd_sc_hd__or2_1
X_1171_ _1243_/A VGND VGND VPWR VPWR _1171_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_27 slave_dat_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 slave_stb_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_16 slave_adr_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0886_ _1580_/C _0878_/X _0883_/X _1590_/B VGND VGND VPWR VPWR _0886_/X sky130_fd_sc_hd__o211a_1
X_0955_ _0955_/A VGND VGND VPWR VPWR _1272_/B sky130_fd_sc_hd__clkbuf_2
X_1507_ _1573_/A VGND VGND VPWR VPWR _1507_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1369_ _1755_/Q _1368_/X _1364_/X _1629_/Q _1361_/X VGND VGND VPWR VPWR _1369_/X
+ sky130_fd_sc_hd__o221a_1
X_1438_ _1720_/Q _1433_/X _1434_/X VGND VGND VPWR VPWR _1720_/D sky130_fd_sc_hd__a21o_1
XFILLER_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput36 slave_dat_i[10] VGND VGND VPWR VPWR input36/X sky130_fd_sc_hd__clkbuf_1
Xinput14 slave_adr_i[20] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_1
Xinput25 slave_adr_i[30] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_1
Xinput47 slave_dat_i[6] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1223_ _1251_/A _1223_/B VGND VGND VPWR VPWR _1224_/A sky130_fd_sc_hd__and2_1
X_1154_ _1161_/A _1154_/B VGND VGND VPWR VPWR _1155_/A sky130_fd_sc_hd__or2_1
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1085_ _1276_/A VGND VGND VPWR VPWR _1086_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0869_ _1600_/C VGND VGND VPWR VPWR _1580_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_0938_ _0948_/A _1402_/C VGND VGND VPWR VPWR _0939_/A sky130_fd_sc_hd__and2_1
XFILLER_11_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1206_ _1242_/A VGND VGND VPWR VPWR _1206_/X sky130_fd_sc_hd__clkbuf_2
X_1137_ _1144_/A _1137_/B VGND VGND VPWR VPWR _1138_/A sky130_fd_sc_hd__and2_1
XFILLER_33_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1068_ _1068_/A VGND VGND VPWR VPWR _1620_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1755_ _1762_/CLK _1755_/D VGND VGND VPWR VPWR _1755_/Q sky130_fd_sc_hd__dfxtp_1
X_1686_ _1712_/CLK _1686_/D VGND VGND VPWR VPWR _1686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1540_ _1554_/A _1540_/B VGND VGND VPWR VPWR _1541_/A sky130_fd_sc_hd__and2_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1471_ _1346_/A _1347_/X _0787_/Y VGND VGND VPWR VPWR _1471_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_40_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1738_ _1766_/CLK _1738_/D VGND VGND VPWR VPWR _1738_/Q sky130_fd_sc_hd__dfxtp_1
X_1669_ _1671_/CLK _1669_/D VGND VGND VPWR VPWR _1669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0971_ _0971_/A VGND VGND VPWR VPWR _0971_/X sky130_fd_sc_hd__clkbuf_1
X_1454_ _1454_/A VGND VGND VPWR VPWR _1729_/D sky130_fd_sc_hd__clkbuf_1
X_1523_ _1556_/A VGND VGND VPWR VPWR _1554_/A sky130_fd_sc_hd__clkbuf_1
X_1385_ _1761_/Q _1382_/X _1378_/X _1635_/Q _1375_/X VGND VGND VPWR VPWR _1385_/X
+ sky130_fd_sc_hd__o221a_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1170_ _1242_/A VGND VGND VPWR VPWR _1170_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_28 slave_dat_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_17 slave_adr_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0885_ _1600_/B VGND VGND VPWR VPWR _1590_/B sky130_fd_sc_hd__clkbuf_2
X_1769__91 VGND VGND VPWR VPWR _1769__91/HI slave_rty_o sky130_fd_sc_hd__conb_1
XANTENNA_39 _1265_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0954_ _0954_/A VGND VGND VPWR VPWR _0954_/X sky130_fd_sc_hd__clkbuf_1
X_1437_ _1437_/A VGND VGND VPWR VPWR _1719_/D sky130_fd_sc_hd__clkbuf_1
X_1506_ _1513_/A _1536_/A _1289_/X VGND VGND VPWR VPWR _1573_/A sky130_fd_sc_hd__o21a_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1299_ _0833_/X _0844_/X _1348_/B _1288_/X _1289_/X VGND VGND VPWR VPWR _1299_/X
+ sky130_fd_sc_hd__o221a_1
X_1368_ _1382_/A VGND VGND VPWR VPWR _1368_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput37 slave_dat_i[11] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_1
Xinput48 slave_dat_i[7] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_1
Xinput26 slave_adr_i[31] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_1
Xinput15 slave_adr_i[21] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1084_ _1622_/Q _1080_/X _1081_/X _1083_/X VGND VGND VPWR VPWR _1622_/D sky130_fd_sc_hd__o211a_1
X_1222_ input10/X _1206_/X _1207_/X _1658_/Q VGND VGND VPWR VPWR _1223_/B sky130_fd_sc_hd__a22o_1
X_1153_ input41/X _1123_/X _1139_/X _1639_/Q VGND VGND VPWR VPWR _1154_/B sky130_fd_sc_hd__o22a_1
X_0868_ _1746_/Q _0879_/B VGND VGND VPWR VPWR _1600_/C sky130_fd_sc_hd__xor2_1
X_0799_ _1734_/Q _1621_/Q VGND VGND VPWR VPWR _1079_/B sky130_fd_sc_hd__nor2b_2
X_0937_ _1703_/Q _0997_/A _0934_/X _1687_/Q _0936_/X VGND VGND VPWR VPWR _1402_/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_28_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1205_ _1205_/A VGND VGND VPWR VPWR _1653_/D sky130_fd_sc_hd__clkbuf_1
X_1136_ input36/X _1134_/X _1135_/X _1634_/Q VGND VGND VPWR VPWR _1137_/B sky130_fd_sc_hd__a22o_1
X_1067_ _1620_/Q _1067_/B VGND VGND VPWR VPWR _1068_/A sky130_fd_sc_hd__or2_1
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1754_ _1762_/CLK _1754_/D VGND VGND VPWR VPWR _1754_/Q sky130_fd_sc_hd__dfxtp_1
X_1685_ _1712_/CLK _1685_/D VGND VGND VPWR VPWR _1685_/Q sky130_fd_sc_hd__dfxtp_1
X_1119_ _1119_/A VGND VGND VPWR VPWR _1629_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1470_ _1738_/Q _1080_/A _1468_/X _1469_/X VGND VGND VPWR VPWR _1738_/D sky130_fd_sc_hd__o211a_1
XFILLER_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1599_ _1599_/A VGND VGND VPWR VPWR _1764_/D sky130_fd_sc_hd__clkbuf_1
X_1737_ _1752_/CLK _1737_/D VGND VGND VPWR VPWR _1737_/Q sky130_fd_sc_hd__dfxtp_2
X_1668_ _1671_/CLK _1668_/D VGND VGND VPWR VPWR _1668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0970_ _1418_/A _0995_/A VGND VGND VPWR VPWR _0971_/A sky130_fd_sc_hd__and2b_1
X_1522_ _1522_/A VGND VGND VPWR VPWR _1751_/D sky130_fd_sc_hd__clkbuf_1
X_1453_ _1729_/Q _1456_/B _1456_/C VGND VGND VPWR VPWR _1454_/A sky130_fd_sc_hd__and3_1
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1384_ _1695_/Q _1381_/X _1383_/X VGND VGND VPWR VPWR _1695_/D sky130_fd_sc_hd__o21a_1
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_29 slave_dat_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_18 slave_adr_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_0884_ _1498_/A _1737_/Q VGND VGND VPWR VPWR _1600_/B sky130_fd_sc_hd__xor2_2
X_0953_ _0980_/A _1409_/A VGND VGND VPWR VPWR _0954_/A sky130_fd_sc_hd__and2_1
X_1505_ _0806_/X _1107_/A _1606_/B _1504_/Y VGND VGND VPWR VPWR _1749_/D sky130_fd_sc_hd__a31o_1
X_1367_ _1381_/A VGND VGND VPWR VPWR _1367_/X sky130_fd_sc_hd__clkbuf_2
X_1436_ _1719_/Q _1439_/B _1439_/C VGND VGND VPWR VPWR _1437_/A sky130_fd_sc_hd__and3_1
X_1298_ _1317_/A VGND VGND VPWR VPWR _1298_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput49 slave_dat_i[8] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_1
Xinput38 slave_dat_i[12] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__clkbuf_1
Xinput27 slave_adr_i[3] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__clkbuf_1
Xinput16 slave_adr_i[22] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__clkbuf_1
X_1221_ _1256_/A VGND VGND VPWR VPWR _1251_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1083_ _1469_/A VGND VGND VPWR VPWR _1083_/X sky130_fd_sc_hd__clkbuf_2
X_1152_ _1152_/A VGND VGND VPWR VPWR _1638_/D sky130_fd_sc_hd__clkbuf_1
X_0936_ _1738_/Q _0993_/B _0993_/C VGND VGND VPWR VPWR _0936_/X sky130_fd_sc_hd__and3_1
XFILLER_9_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0798_ _1640_/Q _1353_/A _1353_/B _1353_/C VGND VGND VPWR VPWR _0798_/X sky130_fd_sc_hd__or4_1
X_0867_ _1698_/Q _1697_/Q _1531_/A VGND VGND VPWR VPWR _0867_/X sky130_fd_sc_hd__mux2_1
X_1419_ _1419_/A _1422_/B VGND VGND VPWR VPWR _1420_/A sky130_fd_sc_hd__or2_1
XFILLER_43_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1204_ _1233_/A _1204_/B VGND VGND VPWR VPWR _1205_/A sky130_fd_sc_hd__or2_1
X_1135_ _1243_/A VGND VGND VPWR VPWR _1135_/X sky130_fd_sc_hd__clkbuf_2
X_1066_ _1066_/A VGND VGND VPWR VPWR _1619_/D sky130_fd_sc_hd__clkbuf_1
X_0919_ _1644_/Q _1040_/B VGND VGND VPWR VPWR _0989_/C sky130_fd_sc_hd__nor2_1
XFILLER_33_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1753_ _1762_/CLK _1753_/D VGND VGND VPWR VPWR _1753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1684_ _1766_/CLK _1684_/D VGND VGND VPWR VPWR _1684_/Q sky130_fd_sc_hd__dfxtp_1
X_1049_ _1049_/A VGND VGND VPWR VPWR _1612_/D sky130_fd_sc_hd__clkbuf_1
X_1118_ _1504_/A _1118_/B VGND VGND VPWR VPWR _1119_/A sky130_fd_sc_hd__or2_1
XFILLER_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1736_ _1752_/CLK _1736_/D VGND VGND VPWR VPWR _1736_/Q sky130_fd_sc_hd__dfxtp_1
X_1598_ _1603_/A _1598_/B VGND VGND VPWR VPWR _1599_/A sky130_fd_sc_hd__and2_1
X_1667_ _1671_/CLK _1667_/D VGND VGND VPWR VPWR _1667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1521_ _1521_/A _1521_/B VGND VGND VPWR VPWR _1522_/A sky130_fd_sc_hd__and2_1
XFILLER_4_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1452_ _1728_/Q _1070_/B _1421_/B VGND VGND VPWR VPWR _1728_/D sky130_fd_sc_hd__a21o_1
X_1383_ _1760_/Q _1382_/X _1378_/X _1634_/Q _1375_/X VGND VGND VPWR VPWR _1383_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1719_ _1732_/CLK _1719_/D VGND VGND VPWR VPWR _1719_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_19 slave_adr_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0952_ _1706_/Q _0940_/X _0934_/X _1690_/Q _0951_/X VGND VGND VPWR VPWR _1409_/A
+ sky130_fd_sc_hd__a221o_1
X_1504_ _1504_/A _1504_/B VGND VGND VPWR VPWR _1504_/Y sky130_fd_sc_hd__nor2_1
X_0883_ _1693_/Q _0892_/S _1590_/C _0882_/X VGND VGND VPWR VPWR _0883_/X sky130_fd_sc_hd__a211o_1
X_1435_ _1718_/Q _1433_/X _1434_/X VGND VGND VPWR VPWR _1718_/D sky130_fd_sc_hd__a21o_1
X_1366_ _1689_/Q _1351_/X _1365_/X VGND VGND VPWR VPWR _1689_/D sky130_fd_sc_hd__o21a_1
X_1297_ _0900_/A _1284_/X _1338_/S VGND VGND VPWR VPWR _1317_/A sky130_fd_sc_hd__a21oi_1
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput39 slave_dat_i[13] VGND VGND VPWR VPWR input39/X sky130_fd_sc_hd__clkbuf_1
Xinput17 slave_adr_i[23] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__clkbuf_1
Xinput28 slave_adr_i[4] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1220_ _1220_/A VGND VGND VPWR VPWR _1657_/D sky130_fd_sc_hd__clkbuf_1
X_1151_ _1180_/A _1151_/B VGND VGND VPWR VPWR _1152_/A sky130_fd_sc_hd__and2_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1082_ _1556_/A VGND VGND VPWR VPWR _1469_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_0866_ _1600_/A VGND VGND VPWR VPWR _1531_/A sky130_fd_sc_hd__clkbuf_2
X_0935_ _1093_/A VGND VGND VPWR VPWR _0993_/B sky130_fd_sc_hd__clkbuf_1
X_0797_ _0797_/A _0797_/B _0797_/C _0797_/D VGND VGND VPWR VPWR _1353_/C sky130_fd_sc_hd__or4_2
X_1418_ _1418_/A _1421_/B VGND VGND VPWR VPWR _1709_/D sky130_fd_sc_hd__nor2_1
X_1349_ _1623_/Q _1622_/Q _1479_/A VGND VGND VPWR VPWR _1382_/A sky130_fd_sc_hd__a21o_2
XFILLER_28_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1203_ input5/X _1195_/X _1175_/X _1653_/Q VGND VGND VPWR VPWR _1204_/B sky130_fd_sc_hd__o22a_1
X_1134_ _1242_/A VGND VGND VPWR VPWR _1134_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1065_ _1402_/A _1619_/Q _1274_/B VGND VGND VPWR VPWR _1066_/A sky130_fd_sc_hd__and3_1
X_0849_ _1767_/Q _1738_/Q VGND VGND VPWR VPWR _1289_/B sky130_fd_sc_hd__nand2_1
X_0918_ _1685_/Q _0961_/B VGND VGND VPWR VPWR _0918_/X sky130_fd_sc_hd__and2_1
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1752_ _1752_/CLK _1752_/D VGND VGND VPWR VPWR _1752_/Q sky130_fd_sc_hd__dfxtp_1
X_1683_ _1740_/CLK _1683_/D VGND VGND VPWR VPWR _1683_/Q sky130_fd_sc_hd__dfxtp_1
X_1117_ input46/X _1074_/X _1102_/X _1629_/Q VGND VGND VPWR VPWR _1118_/B sky130_fd_sc_hd__o22a_1
X_1048_ _1048_/A _1612_/Q _1477_/B VGND VGND VPWR VPWR _1049_/A sky130_fd_sc_hd__and3_1
XFILLER_21_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1735_ _1752_/CLK _1735_/D VGND VGND VPWR VPWR _1735_/Q sky130_fd_sc_hd__dfxtp_1
X_1666_ _1671_/CLK _1666_/D VGND VGND VPWR VPWR _1666_/Q sky130_fd_sc_hd__dfxtp_1
X_1597_ _1764_/Q _1573_/X _1596_/X _1576_/X VGND VGND VPWR VPWR _1598_/B sky130_fd_sc_hd__a22o_1
XFILLER_14_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1520_ _1751_/Q _1507_/X _1519_/X _1514_/X VGND VGND VPWR VPWR _1521_/B sky130_fd_sc_hd__a22o_1
X_1451_ _1451_/A VGND VGND VPWR VPWR _1727_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1382_ _1382_/A VGND VGND VPWR VPWR _1382_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1718_ _1732_/CLK _1718_/D VGND VGND VPWR VPWR _1718_/Q sky130_fd_sc_hd__dfxtp_1
X_1649_ _1650_/CLK _1649_/D VGND VGND VPWR VPWR _1649_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0882_ _1694_/Q _0900_/A _1550_/A VGND VGND VPWR VPWR _0882_/X sky130_fd_sc_hd__and3_1
X_0951_ _0951_/A _0955_/A _1079_/C VGND VGND VPWR VPWR _0951_/X sky130_fd_sc_hd__and3_1
X_1503_ _1503_/A VGND VGND VPWR VPWR _1748_/D sky130_fd_sc_hd__clkbuf_1
X_1296_ _0844_/X _1294_/X _1295_/X VGND VGND VPWR VPWR _1676_/D sky130_fd_sc_hd__o21ba_1
X_1365_ _1754_/Q _1352_/X _1364_/X _1628_/Q _1361_/X VGND VGND VPWR VPWR _1365_/X
+ sky130_fd_sc_hd__o221a_1
X_1434_ _1459_/B VGND VGND VPWR VPWR _1434_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 slave_adr_i[24] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_1
Xinput29 slave_adr_i[5] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1150_ input40/X _1134_/X _1135_/X _1638_/Q VGND VGND VPWR VPWR _1151_/B sky130_fd_sc_hd__a22o_1
X_1081_ _1639_/Q _1274_/B VGND VGND VPWR VPWR _1081_/X sky130_fd_sc_hd__or2_1
XFILLER_20_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0934_ _0967_/A VGND VGND VPWR VPWR _0934_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0865_ _1700_/Q _1699_/Q _0892_/S VGND VGND VPWR VPWR _0865_/X sky130_fd_sc_hd__mux2_1
X_0796_ _1672_/Q _1671_/Q _1670_/Q _1669_/Q VGND VGND VPWR VPWR _0797_/D sky130_fd_sc_hd__or4_1
X_1417_ _1459_/B VGND VGND VPWR VPWR _1421_/B sky130_fd_sc_hd__clkbuf_2
X_1279_ _1603_/A VGND VGND VPWR VPWR _1279_/X sky130_fd_sc_hd__clkbuf_2
X_1348_ _1348_/A _1348_/B _1288_/X VGND VGND VPWR VPWR _1479_/A sky130_fd_sc_hd__or3b_1
XFILLER_47_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1064_ _1064_/A VGND VGND VPWR VPWR _1618_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1202_ _1411_/A VGND VGND VPWR VPWR _1233_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1133_ _1133_/A VGND VGND VPWR VPWR _1633_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0848_ _0847_/A _0847_/C _1513_/A _1674_/Q VGND VGND VPWR VPWR _0848_/X sky130_fd_sc_hd__a31o_1
X_0917_ _1040_/B VGND VGND VPWR VPWR _0961_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1751_ _1752_/CLK _1751_/D VGND VGND VPWR VPWR _1751_/Q sky130_fd_sc_hd__dfxtp_1
X_1682_ _1740_/CLK _1682_/D VGND VGND VPWR VPWR _1682_/Q sky130_fd_sc_hd__dfxtp_1
X_1047_ _1047_/A VGND VGND VPWR VPWR _1611_/D sky130_fd_sc_hd__clkbuf_1
X_1116_ _1116_/A VGND VGND VPWR VPWR _1628_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1596_ _1764_/Q _1562_/A _1596_/S VGND VGND VPWR VPWR _1596_/X sky130_fd_sc_hd__mux2_1
X_1665_ _1671_/CLK _1665_/D VGND VGND VPWR VPWR _1665_/Q sky130_fd_sc_hd__dfxtp_1
X_1734_ _1734_/CLK _1734_/D VGND VGND VPWR VPWR _1734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1450_ _1727_/Q _1456_/B _1456_/C VGND VGND VPWR VPWR _1451_/A sky130_fd_sc_hd__and3_1
X_1381_ _1381_/A VGND VGND VPWR VPWR _1381_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1579_ _1579_/A VGND VGND VPWR VPWR _1760_/D sky130_fd_sc_hd__clkbuf_1
X_1717_ _1717_/CLK _1717_/D VGND VGND VPWR VPWR _1717_/Q sky130_fd_sc_hd__dfxtp_1
X_1648_ _1650_/CLK _1648_/D VGND VGND VPWR VPWR _1648_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0881_ _1509_/C VGND VGND VPWR VPWR _1550_/A sky130_fd_sc_hd__clkbuf_1
X_0950_ _1034_/C VGND VGND VPWR VPWR _0980_/A sky130_fd_sc_hd__clkbuf_1
X_1502_ _1502_/A _1502_/B VGND VGND VPWR VPWR _1503_/A sky130_fd_sc_hd__or2_1
X_1433_ _1433_/A VGND VGND VPWR VPWR _1433_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1295_ _0806_/X _0844_/X _1310_/A _1502_/A VGND VGND VPWR VPWR _1295_/X sky130_fd_sc_hd__a31o_1
X_1364_ _1378_/A VGND VGND VPWR VPWR _1364_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput19 slave_adr_i[25] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1080_ _1080_/A VGND VGND VPWR VPWR _1080_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0864_ _1600_/A VGND VGND VPWR VPWR _0892_/S sky130_fd_sc_hd__clkbuf_2
X_0795_ _1664_/Q _1663_/Q _1662_/Q _1661_/Q VGND VGND VPWR VPWR _0797_/C sky130_fd_sc_hd__or4_1
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0933_ _1093_/A _1040_/B VGND VGND VPWR VPWR _0967_/A sky130_fd_sc_hd__and2_1
X_1416_ _1416_/A VGND VGND VPWR VPWR _1708_/D sky130_fd_sc_hd__clkbuf_1
X_1347_ _1353_/A _1353_/B _1353_/C _1347_/D VGND VGND VPWR VPWR _1347_/X sky130_fd_sc_hd__or4_2
XFILLER_36_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1278_ _1556_/A VGND VGND VPWR VPWR _1603_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1201_ _1201_/A VGND VGND VPWR VPWR _1652_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1063_ _1618_/Q _1063_/B VGND VGND VPWR VPWR _1064_/A sky130_fd_sc_hd__or2_1
X_1132_ _1161_/A _1132_/B VGND VGND VPWR VPWR _1133_/A sky130_fd_sc_hd__or2_1
XFILLER_33_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0916_ _0916_/A VGND VGND VPWR VPWR _1040_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_0847_ _0847_/A _1674_/Q _0847_/C _1513_/A VGND VGND VPWR VPWR _0847_/Y sky130_fd_sc_hd__nand4_1
XFILLER_33_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1750_ _1752_/CLK _1750_/D VGND VGND VPWR VPWR _1750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1681_ _1740_/CLK _1681_/D VGND VGND VPWR VPWR _1681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1046_ _1611_/Q _1063_/B VGND VGND VPWR VPWR _1047_/A sky130_fd_sc_hd__or2_1
X_1115_ _1144_/A _1115_/B VGND VGND VPWR VPWR _1116_/A sky130_fd_sc_hd__and2_1
XFILLER_21_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1733_ _1733_/CLK _1733_/D VGND VGND VPWR VPWR _1733_/Q sky130_fd_sc_hd__dfxtp_1
X_1595_ _1595_/A _1595_/B VGND VGND VPWR VPWR _1596_/S sky130_fd_sc_hd__nor2_1
X_1664_ _1671_/CLK _1664_/D VGND VGND VPWR VPWR _1664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1029_ _1730_/Q _1029_/B _1029_/C VGND VGND VPWR VPWR _1030_/A sky130_fd_sc_hd__and3_1
XFILLER_30_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1380_ _1694_/Q _1367_/X _1379_/X VGND VGND VPWR VPWR _1694_/D sky130_fd_sc_hd__o21a_1
X_1716_ _1734_/CLK _1716_/D VGND VGND VPWR VPWR _1716_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1578_ _1583_/A _1578_/B VGND VGND VPWR VPWR _1579_/A sky130_fd_sc_hd__and2_1
XFILLER_6_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1647_ _1650_/CLK _1647_/D VGND VGND VPWR VPWR _1647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0880_ _1536_/D VGND VGND VPWR VPWR _1590_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_1501_ _1748_/Q _1488_/A _1499_/Y _1500_/X VGND VGND VPWR VPWR _1502_/B sky130_fd_sc_hd__o22a_1
X_1432_ _1432_/A VGND VGND VPWR VPWR _1717_/D sky130_fd_sc_hd__clkbuf_1
X_1363_ _1688_/Q _1351_/X _1362_/X VGND VGND VPWR VPWR _1688_/D sky130_fd_sc_hd__o21a_1
XFILLER_48_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1294_ _1310_/A VGND VGND VPWR VPWR _1294_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0932_ _1347_/D VGND VGND VPWR VPWR _0997_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_0863_ _0894_/A _1509_/C VGND VGND VPWR VPWR _1600_/A sky130_fd_sc_hd__nand2_1
X_0794_ _1660_/Q _1659_/Q _1658_/Q _1657_/Q VGND VGND VPWR VPWR _0797_/B sky130_fd_sc_hd__or4_1
X_1346_ _1346_/A VGND VGND VPWR VPWR _1346_/Y sky130_fd_sc_hd__inv_2
X_1415_ _1415_/A _1422_/B VGND VGND VPWR VPWR _1416_/A sky130_fd_sc_hd__or2_1
X_1277_ _1625_/Q _1608_/B VGND VGND VPWR VPWR _1277_/X sky130_fd_sc_hd__or2_1
XFILLER_42_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1200_ _1216_/A _1200_/B VGND VGND VPWR VPWR _1201_/A sky130_fd_sc_hd__and2_1
XFILLER_33_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1062_ _1062_/A VGND VGND VPWR VPWR _1617_/D sky130_fd_sc_hd__clkbuf_1
X_1131_ input50/X _1123_/X _1102_/X _1633_/Q VGND VGND VPWR VPWR _1132_/B sky130_fd_sc_hd__o22a_1
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0915_ _1093_/A VGND VGND VPWR VPWR _0955_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_0846_ _0846_/A _0846_/B _0846_/C _0845_/X VGND VGND VPWR VPWR _1513_/A sky130_fd_sc_hd__or4b_2
X_1329_ _1606_/A VGND VGND VPWR VPWR _1329_/X sky130_fd_sc_hd__buf_2
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1680_ _1740_/CLK _1680_/D VGND VGND VPWR VPWR _1680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1114_ input45/X _1092_/X _1094_/X _1628_/Q VGND VGND VPWR VPWR _1115_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1045_ _1067_/B VGND VGND VPWR VPWR _1063_/B sky130_fd_sc_hd__clkbuf_1
X_0829_ _0826_/A _0946_/A _0942_/A VGND VGND VPWR VPWR _1319_/A sky130_fd_sc_hd__nand3b_1
XFILLER_9_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1663_ _1671_/CLK _1663_/D VGND VGND VPWR VPWR _1663_/Q sky130_fd_sc_hd__dfxtp_1
X_1732_ _1732_/CLK _1732_/D VGND VGND VPWR VPWR _1732_/Q sky130_fd_sc_hd__dfxtp_1
X_1594_ _1594_/A VGND VGND VPWR VPWR _1763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1028_ _1028_/A VGND VGND VPWR VPWR _1028_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1715_ _1734_/CLK _1715_/D VGND VGND VPWR VPWR _1715_/Q sky130_fd_sc_hd__dfxtp_1
X_1646_ _1650_/CLK _1646_/D VGND VGND VPWR VPWR _1646_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1577_ _1760_/Q _1573_/X _1575_/X _1576_/X VGND VGND VPWR VPWR _1578_/B sky130_fd_sc_hd__a22o_1
XFILLER_41_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1500_ _1509_/A _1748_/Q _1498_/Y _1504_/B VGND VGND VPWR VPWR _1500_/X sky130_fd_sc_hd__a31o_1
X_1293_ _0900_/A _1284_/X _1338_/S VGND VGND VPWR VPWR _1310_/A sky130_fd_sc_hd__a21o_1
X_1362_ _1753_/Q _1352_/X _1462_/B _1627_/Q _1361_/X VGND VGND VPWR VPWR _1362_/X
+ sky130_fd_sc_hd__o221a_1
X_1431_ _1717_/Q _1439_/B _1439_/C VGND VGND VPWR VPWR _1432_/A sky130_fd_sc_hd__and3_1
X_1629_ _1717_/CLK _1629_/D VGND VGND VPWR VPWR _1629_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_46_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0862_ _1745_/Q _1737_/Q VGND VGND VPWR VPWR _1509_/C sky130_fd_sc_hd__xnor2_1
X_0931_ _0931_/A VGND VGND VPWR VPWR _0931_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0793_ _1668_/Q _1667_/Q _1666_/Q _1665_/Q VGND VGND VPWR VPWR _0797_/A sky130_fd_sc_hd__or4_1
X_1345_ _1294_/X _1343_/Y _1344_/X VGND VGND VPWR VPWR _1684_/D sky130_fd_sc_hd__a21oi_1
X_1414_ _1414_/A VGND VGND VPWR VPWR _1707_/D sky130_fd_sc_hd__clkbuf_1
X_1276_ _1276_/A VGND VGND VPWR VPWR _1608_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1130_ _1502_/A VGND VGND VPWR VPWR _1161_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1061_ _1617_/Q _1063_/B VGND VGND VPWR VPWR _1062_/A sky130_fd_sc_hd__or2_1
X_0845_ _0833_/X _0834_/X _0835_/X _0844_/X _0847_/A VGND VGND VPWR VPWR _0845_/X
+ sky130_fd_sc_hd__o221a_1
X_0914_ _1034_/C VGND VGND VPWR VPWR _0948_/A sky130_fd_sc_hd__clkbuf_1
X_1328_ _1333_/A _1333_/B _1298_/X VGND VGND VPWR VPWR _1328_/X sky130_fd_sc_hd__a21o_1
X_1259_ _1259_/A VGND VGND VPWR VPWR _1668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1113_ _1256_/A VGND VGND VPWR VPWR _1144_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1044_ _1375_/A _1276_/A VGND VGND VPWR VPWR _1067_/B sky130_fd_sc_hd__nand2_1
X_0828_ _0828_/A VGND VGND VPWR VPWR _0942_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1662_ _1662_/CLK _1662_/D VGND VGND VPWR VPWR _1662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1731_ _1732_/CLK _1731_/D VGND VGND VPWR VPWR _1731_/Q sky130_fd_sc_hd__dfxtp_1
X_1593_ _1603_/A _1593_/B VGND VGND VPWR VPWR _1594_/A sky130_fd_sc_hd__and2_1
X_1027_ _1729_/Q _1029_/B _1029_/C VGND VGND VPWR VPWR _1028_/A sky130_fd_sc_hd__and3_1
XFILLER_39_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1576_ _1576_/A VGND VGND VPWR VPWR _1576_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1714_ _1734_/CLK _1714_/D VGND VGND VPWR VPWR _1714_/Q sky130_fd_sc_hd__dfxtp_1
X_1645_ _1650_/CLK _1645_/D VGND VGND VPWR VPWR _1645_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1430_ _1430_/A VGND VGND VPWR VPWR _1716_/D sky130_fd_sc_hd__clkbuf_1
X_1292_ _1486_/A VGND VGND VPWR VPWR _1338_/S sky130_fd_sc_hd__clkbuf_2
X_1361_ _1375_/A VGND VGND VPWR VPWR _1361_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xoutput80 _0945_/X VGND VGND VPWR VPWR slave_dat_o[3] sky130_fd_sc_hd__buf_2
XFILLER_31_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1559_ _1757_/Q _1542_/X _1558_/X _1546_/X VGND VGND VPWR VPWR _1560_/B sky130_fd_sc_hd__a22o_1
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1628_ _1717_/CLK _1628_/D VGND VGND VPWR VPWR _1628_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_36_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0861_ _1580_/B VGND VGND VPWR VPWR _1568_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_0930_ _0948_/A _1400_/A VGND VGND VPWR VPWR _0931_/A sky130_fd_sc_hd__and2_1
X_0792_ _1656_/Q _1655_/Q _0792_/C _0792_/D VGND VGND VPWR VPWR _1353_/B sky130_fd_sc_hd__or4_2
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1413_ _1413_/A _1439_/C VGND VGND VPWR VPWR _1414_/A sky130_fd_sc_hd__and2_1
X_1344_ _0847_/A _1298_/X _1502_/A VGND VGND VPWR VPWR _1344_/X sky130_fd_sc_hd__a21o_1
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1275_ _1674_/Q _1080_/X _1274_/X _1083_/X VGND VGND VPWR VPWR _1674_/D sky130_fd_sc_hd__o211a_1
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1060_ _1060_/A VGND VGND VPWR VPWR _1616_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0844_ _1676_/Q VGND VGND VPWR VPWR _0844_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_0913_ _1020_/A VGND VGND VPWR VPWR _1034_/C sky130_fd_sc_hd__clkbuf_2
X_1327_ _1333_/A _1333_/B VGND VGND VPWR VPWR _1327_/Y sky130_fd_sc_hd__nor2_1
X_1258_ _1521_/A _1258_/B VGND VGND VPWR VPWR _1259_/A sky130_fd_sc_hd__and2_1
X_1189_ input32/X _1159_/X _1175_/X _1649_/Q VGND VGND VPWR VPWR _1190_/B sky130_fd_sc_hd__o22a_1
XFILLER_24_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1043_ _1043_/A VGND VGND VPWR VPWR _1610_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1112_ _1375_/A VGND VGND VPWR VPWR _1256_/A sky130_fd_sc_hd__clkbuf_2
X_0827_ _1679_/Q VGND VGND VPWR VPWR _0830_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1592_ _1763_/Q _1573_/X _1591_/X _1576_/X VGND VGND VPWR VPWR _1593_/B sky130_fd_sc_hd__a22o_1
X_1661_ _1662_/CLK _1661_/D VGND VGND VPWR VPWR _1661_/Q sky130_fd_sc_hd__dfxtp_1
X_1730_ _1730_/CLK _1730_/D VGND VGND VPWR VPWR _1730_/Q sky130_fd_sc_hd__dfxtp_1
X_1026_ _1026_/A VGND VGND VPWR VPWR _1026_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1713_ _1730_/CLK _1713_/D VGND VGND VPWR VPWR _1713_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_0 slave_adr_i[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1575_ _1760_/Q _1524_/X _1575_/S VGND VGND VPWR VPWR _1575_/X sky130_fd_sc_hd__mux2_1
X_1644_ _1650_/CLK _1644_/D VGND VGND VPWR VPWR _1644_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1009_ _1721_/Q _1017_/B _1017_/C VGND VGND VPWR VPWR _1010_/A sky130_fd_sc_hd__and3_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_9_0_CLK clkbuf_4_9_0_CLK/A VGND VGND VPWR VPWR _1734_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1360_ _1687_/Q _1351_/X _1359_/X VGND VGND VPWR VPWR _1687_/D sky130_fd_sc_hd__o21a_1
Xoutput70 _1016_/X VGND VGND VPWR VPWR slave_dat_o[23] sky130_fd_sc_hd__buf_2
X_1291_ _1314_/S VGND VGND VPWR VPWR _1486_/A sky130_fd_sc_hd__clkbuf_2
Xoutput81 _0949_/X VGND VGND VPWR VPWR slave_dat_o[4] sky130_fd_sc_hd__buf_2
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1489_ _1491_/A _1745_/Q _1488_/X VGND VGND VPWR VPWR _1489_/Y sky130_fd_sc_hd__o21ai_1
X_1558_ _1508_/X _1757_/Q _1558_/S VGND VGND VPWR VPWR _1558_/X sky130_fd_sc_hd__mux2_1
X_1627_ _1717_/CLK _1627_/D VGND VGND VPWR VPWR _1627_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0860_ _1498_/A _0879_/B VGND VGND VPWR VPWR _1580_/B sky130_fd_sc_hd__xnor2_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0791_ _1654_/Q _1653_/Q _1652_/Q _1651_/Q VGND VGND VPWR VPWR _0792_/D sky130_fd_sc_hd__or4_1
X_1343_ _1684_/Q _1342_/B _1339_/A _1339_/B _1342_/Y VGND VGND VPWR VPWR _1343_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1412_ _1443_/A VGND VGND VPWR VPWR _1439_/C sky130_fd_sc_hd__clkbuf_2
X_1274_ _1624_/Q _1274_/B VGND VGND VPWR VPWR _1274_/X sky130_fd_sc_hd__or2_1
XFILLER_22_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0989_ _1623_/Q _0993_/B _0989_/C VGND VGND VPWR VPWR _0989_/X sky130_fd_sc_hd__and3_1
XFILLER_27_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0912_ _1395_/A _1459_/A VGND VGND VPWR VPWR _1020_/A sky130_fd_sc_hd__nor2_2
X_0843_ _0846_/A _0840_/X _0842_/X VGND VGND VPWR VPWR _0847_/C sky130_fd_sc_hd__o21ai_1
X_1326_ _1681_/Q _1325_/Y _1486_/A VGND VGND VPWR VPWR _1333_/B sky130_fd_sc_hd__mux2_1
X_1257_ input21/X _1242_/X _1243_/X _1668_/Q VGND VGND VPWR VPWR _1258_/B sky130_fd_sc_hd__a22o_1
XFILLER_17_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1188_ _1188_/A VGND VGND VPWR VPWR _1648_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1042_ _1048_/A _1610_/Q _1477_/B VGND VGND VPWR VPWR _1043_/A sky130_fd_sc_hd__and3_1
X_1111_ _1111_/A VGND VGND VPWR VPWR _1627_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0826_ _0826_/A _0828_/A _1741_/Q VGND VGND VPWR VPWR _1313_/A sky130_fd_sc_hd__or3b_1
X_1309_ _1300_/X _1308_/X _1298_/X VGND VGND VPWR VPWR _1309_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1591_ _1562_/X _1763_/Q _1591_/S VGND VGND VPWR VPWR _1591_/X sky130_fd_sc_hd__mux2_1
X_1660_ _1662_/CLK _1660_/D VGND VGND VPWR VPWR _1660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1025_ _1728_/Q _1029_/B _1029_/C VGND VGND VPWR VPWR _1026_/A sky130_fd_sc_hd__and3_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0809_ _1742_/Q VGND VGND VPWR VPWR _1477_/A sky130_fd_sc_hd__inv_2
XFILLER_29_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1 slave_adr_i[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1643_ _1650_/CLK _1643_/D VGND VGND VPWR VPWR _1643_/Q sky130_fd_sc_hd__dfxtp_1
X_1712_ _1712_/CLK _1712_/D VGND VGND VPWR VPWR _1712_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1574_ _1595_/A _1574_/B VGND VGND VPWR VPWR _1575_/S sky130_fd_sc_hd__nor2_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1008_ _1020_/A VGND VGND VPWR VPWR _1017_/C sky130_fd_sc_hd__clkbuf_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput82 _0954_/X VGND VGND VPWR VPWR slave_dat_o[5] sky130_fd_sc_hd__buf_2
Xoutput60 _0992_/X VGND VGND VPWR VPWR slave_dat_o[14] sky130_fd_sc_hd__buf_2
Xoutput71 _1018_/X VGND VGND VPWR VPWR slave_dat_o[24] sky130_fd_sc_hd__buf_2
XFILLER_48_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1290_ _1348_/B _1288_/X _1289_/X VGND VGND VPWR VPWR _1314_/S sky130_fd_sc_hd__o21ai_1
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1626_ _1717_/CLK _1626_/D VGND VGND VPWR VPWR _1626_/Q sky130_fd_sc_hd__dfxtp_1
X_1488_ _1488_/A VGND VGND VPWR VPWR _1488_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1557_ _1590_/A _1590_/B _1580_/C _1557_/D VGND VGND VPWR VPWR _1558_/S sky130_fd_sc_hd__or4_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0790_ _1650_/Q _1649_/Q _1642_/Q _1641_/Q VGND VGND VPWR VPWR _0792_/C sky130_fd_sc_hd__or4_1
X_1342_ _1342_/A _1342_/B VGND VGND VPWR VPWR _1342_/Y sky130_fd_sc_hd__nand2_1
X_1411_ _1411_/A _1411_/B VGND VGND VPWR VPWR _1443_/A sky130_fd_sc_hd__nor2_1
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1273_ _1074_/X _1272_/X _1305_/A VGND VGND VPWR VPWR _1673_/D sky130_fd_sc_hd__a21oi_1
XFILLER_36_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0988_ _0988_/A VGND VGND VPWR VPWR _0988_/X sky130_fd_sc_hd__clkbuf_1
X_1609_ _1767_/Q _1080_/A _1608_/X _1329_/X VGND VGND VPWR VPWR _1767_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_4_8_0_CLK clkbuf_4_9_0_CLK/A VGND VGND VPWR VPWR _1717_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0842_ _0808_/X _1342_/A _0824_/A _0841_/X VGND VGND VPWR VPWR _0842_/X sky130_fd_sc_hd__a22o_1
X_0911_ _1079_/B _0798_/X _0907_/X _1347_/D _0910_/Y VGND VGND VPWR VPWR _1459_/A
+ sky130_fd_sc_hd__a32o_1
X_1325_ _1325_/A VGND VGND VPWR VPWR _1325_/Y sky130_fd_sc_hd__inv_2
X_1256_ _1256_/A VGND VGND VPWR VPWR _1521_/A sky130_fd_sc_hd__buf_2
XFILLER_33_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1187_ _1216_/A _1187_/B VGND VGND VPWR VPWR _1188_/A sky130_fd_sc_hd__and2_1
XFILLER_24_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1110_ _1504_/A _1110_/B VGND VGND VPWR VPWR _1111_/A sky130_fd_sc_hd__or2_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1041_ _1276_/A VGND VGND VPWR VPWR _1477_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0825_ _1678_/Q VGND VGND VPWR VPWR _0825_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1308_ _1477_/A _1475_/A _0942_/A _1342_/B _1306_/X VGND VGND VPWR VPWR _1308_/X
+ sky130_fd_sc_hd__a41o_1
X_1239_ input16/X _1231_/X _1211_/X _1663_/Q VGND VGND VPWR VPWR _1240_/B sky130_fd_sc_hd__o22a_1
XFILLER_44_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1590_ _1590_/A _1590_/B _1590_/C _1600_/D VGND VGND VPWR VPWR _1591_/S sky130_fd_sc_hd__or4_1
XFILLER_38_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1024_ _1024_/A VGND VGND VPWR VPWR _1024_/X sky130_fd_sc_hd__clkbuf_1
X_0808_ _1683_/Q VGND VGND VPWR VPWR _0808_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_2 slave_adr_i[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1642_ _1650_/CLK _1642_/D VGND VGND VPWR VPWR _1642_/Q sky130_fd_sc_hd__dfxtp_1
X_1711_ _1730_/CLK _1711_/D VGND VGND VPWR VPWR _1711_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1573_ _1573_/A VGND VGND VPWR VPWR _1573_/X sky130_fd_sc_hd__clkbuf_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1007_ _1069_/A VGND VGND VPWR VPWR _1017_/B sky130_fd_sc_hd__clkbuf_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput83 _0960_/X VGND VGND VPWR VPWR slave_dat_o[6] sky130_fd_sc_hd__buf_2
Xoutput72 _1022_/X VGND VGND VPWR VPWR slave_dat_o[25] sky130_fd_sc_hd__buf_2
Xoutput61 _0996_/X VGND VGND VPWR VPWR slave_dat_o[15] sky130_fd_sc_hd__buf_2
XFILLER_48_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1556_ _1556_/A VGND VGND VPWR VPWR _1583_/A sky130_fd_sc_hd__clkbuf_1
X_1768__90 VGND VGND VPWR VPWR _1768__90/HI slave_err_o sky130_fd_sc_hd__conb_1
X_1625_ _1671_/CLK _1625_/D VGND VGND VPWR VPWR _1625_/Q sky130_fd_sc_hd__dfxtp_1
X_1487_ _1504_/B _1606_/B VGND VGND VPWR VPWR _1488_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1410_ _1410_/A VGND VGND VPWR VPWR _1706_/D sky130_fd_sc_hd__clkbuf_1
X_1341_ _0808_/X _1323_/A _1339_/Y _1340_/X _1329_/X VGND VGND VPWR VPWR _1683_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1272_ _1734_/Q _1272_/B _1673_/Q VGND VGND VPWR VPWR _1272_/X sky130_fd_sc_hd__or3b_1
XFILLER_36_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0987_ _0995_/A _1425_/A VGND VGND VPWR VPWR _0988_/A sky130_fd_sc_hd__and2_1
XFILLER_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1539_ _1754_/Q _1507_/X _1538_/X _1514_/X VGND VGND VPWR VPWR _1540_/B sky130_fd_sc_hd__a22o_1
X_1608_ _1630_/Q _1608_/B VGND VGND VPWR VPWR _1608_/X sky130_fd_sc_hd__or2_1
XFILLER_27_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0841_ _0841_/A _0841_/B VGND VGND VPWR VPWR _0841_/X sky130_fd_sc_hd__or2_1
X_0910_ _1733_/Q VGND VGND VPWR VPWR _0910_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1324_ _1680_/Q _1294_/X _1323_/Y _1279_/X VGND VGND VPWR VPWR _1680_/D sky130_fd_sc_hd__o211a_1
X_1186_ input31/X _1170_/X _1171_/X _1648_/Q VGND VGND VPWR VPWR _1187_/B sky130_fd_sc_hd__a22o_1
X_1255_ _1255_/A VGND VGND VPWR VPWR _1667_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1040_ _1644_/Q _1040_/B _1353_/D VGND VGND VPWR VPWR _1276_/A sky130_fd_sc_hd__or3_2
Xclkbuf_4_7_0_CLK clkbuf_4_7_0_CLK/A VGND VGND VPWR VPWR _1766_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0824_ _0824_/A _0841_/A _0824_/C VGND VGND VPWR VPWR _0846_/A sky130_fd_sc_hd__nand3_1
XFILLER_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1307_ _1477_/A _1475_/A _1314_/S _1299_/X _1306_/X VGND VGND VPWR VPWR _1321_/A
+ sky130_fd_sc_hd__a311o_1
X_1238_ _1411_/A VGND VGND VPWR VPWR _1267_/A sky130_fd_sc_hd__clkbuf_1
X_1169_ _1169_/A VGND VGND VPWR VPWR _1643_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1023_ _1727_/Q _1029_/B _1029_/C VGND VGND VPWR VPWR _1024_/A sky130_fd_sc_hd__and3_1
X_0807_ _1684_/Q VGND VGND VPWR VPWR _0847_/A sky130_fd_sc_hd__inv_2
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_3 slave_adr_i[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1572_ _1572_/A VGND VGND VPWR VPWR _1759_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1641_ _1662_/CLK _1641_/D VGND VGND VPWR VPWR _1641_/Q sky130_fd_sc_hd__dfxtp_1
X_1710_ _1730_/CLK _1710_/D VGND VGND VPWR VPWR _1710_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1006_ _1006_/A VGND VGND VPWR VPWR _1006_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput84 _0965_/X VGND VGND VPWR VPWR slave_dat_o[7] sky130_fd_sc_hd__buf_2
Xoutput62 _1000_/X VGND VGND VPWR VPWR slave_dat_o[16] sky130_fd_sc_hd__buf_2
Xoutput73 _1024_/X VGND VGND VPWR VPWR slave_dat_o[26] sky130_fd_sc_hd__buf_2
XFILLER_48_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1555_ _1555_/A VGND VGND VPWR VPWR _1756_/D sky130_fd_sc_hd__clkbuf_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1624_ _1733_/CLK _1624_/D VGND VGND VPWR VPWR _1624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1486_ _1486_/A VGND VGND VPWR VPWR _1504_/B sky130_fd_sc_hd__inv_2
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1340_ _1339_/A _1339_/B _1298_/X VGND VGND VPWR VPWR _1340_/X sky130_fd_sc_hd__a21o_1
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1271_ _1271_/A VGND VGND VPWR VPWR _1672_/D sky130_fd_sc_hd__clkbuf_1
X_0986_ _1714_/Q _0940_/X _0967_/X _1698_/Q VGND VGND VPWR VPWR _1425_/A sky130_fd_sc_hd__a22o_1
X_1538_ _1754_/Q _1524_/X _1538_/S VGND VGND VPWR VPWR _1538_/X sky130_fd_sc_hd__mux2_1
X_1607_ _1607_/A VGND VGND VPWR VPWR _1766_/D sky130_fd_sc_hd__clkbuf_1
X_1469_ _1469_/A VGND VGND VPWR VPWR _1469_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0840_ _0846_/B _0837_/X _0839_/X VGND VGND VPWR VPWR _0840_/X sky130_fd_sc_hd__o21a_1
X_1323_ _1323_/A _1333_/A _1323_/C VGND VGND VPWR VPWR _1323_/Y sky130_fd_sc_hd__nand3_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1254_ _1267_/A _1254_/B VGND VGND VPWR VPWR _1255_/A sky130_fd_sc_hd__or2_1
X_1185_ _1256_/A VGND VGND VPWR VPWR _1216_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_0969_ _1034_/C VGND VGND VPWR VPWR _0995_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_9_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0823_ _0808_/X _1342_/A _1325_/A _1680_/Q _0841_/B VGND VGND VPWR VPWR _0824_/C
+ sky130_fd_sc_hd__a221oi_1
X_1306_ _1348_/B _1288_/X _1289_/X _0825_/X VGND VGND VPWR VPWR _1306_/X sky130_fd_sc_hd__o211a_1
X_1237_ _1237_/A VGND VGND VPWR VPWR _1662_/D sky130_fd_sc_hd__clkbuf_1
X_1099_ _1411_/A VGND VGND VPWR VPWR _1504_/A sky130_fd_sc_hd__clkbuf_2
X_1168_ _1197_/A _1168_/B VGND VGND VPWR VPWR _1169_/A sky130_fd_sc_hd__or2_1
XFILLER_20_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1022_ _1022_/A VGND VGND VPWR VPWR _1022_/X sky130_fd_sc_hd__clkbuf_1
X_0806_ _1509_/A VGND VGND VPWR VPWR _0806_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_6_0_CLK clkbuf_4_7_0_CLK/A VGND VGND VPWR VPWR _1767_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_4 slave_adr_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1571_ _1583_/A _1571_/B VGND VGND VPWR VPWR _1572_/A sky130_fd_sc_hd__and2_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1640_ _1650_/CLK _1640_/D VGND VGND VPWR VPWR _1640_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1005_ _1720_/Q _1433_/A _1005_/C VGND VGND VPWR VPWR _1006_/A sky130_fd_sc_hd__and3_1
XFILLER_41_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput85 _0971_/X VGND VGND VPWR VPWR slave_dat_o[8] sky130_fd_sc_hd__buf_2
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput63 _1002_/X VGND VGND VPWR VPWR slave_dat_o[17] sky130_fd_sc_hd__buf_2
Xoutput74 _1026_/X VGND VGND VPWR VPWR slave_dat_o[27] sky130_fd_sc_hd__buf_2
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1554_ _1554_/A _1554_/B VGND VGND VPWR VPWR _1555_/A sky130_fd_sc_hd__and2_1
X_1623_ _1767_/CLK _1623_/D VGND VGND VPWR VPWR _1623_/Q sky130_fd_sc_hd__dfxtp_1
X_1485_ _0921_/A _1070_/B _0961_/B _1484_/X _1329_/X VGND VGND VPWR VPWR _1744_/D
+ sky130_fd_sc_hd__o311a_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

