magic
tech sky130A
magscale 1 2
timestamp 1647793929
<< obsli1 >>
rect 1104 2159 53360 54417
<< obsm1 >>
rect 106 8 54450 55820
<< metal2 >>
rect 110 55850 166 56650
rect 294 55850 350 56650
rect 570 55850 626 56650
rect 846 55850 902 56650
rect 1122 55850 1178 56650
rect 1398 55850 1454 56650
rect 1674 55850 1730 56650
rect 1950 55850 2006 56650
rect 2226 55850 2282 56650
rect 2502 55850 2558 56650
rect 2778 55850 2834 56650
rect 2962 55850 3018 56650
rect 3238 55850 3294 56650
rect 3514 55850 3570 56650
rect 3790 55850 3846 56650
rect 4066 55850 4122 56650
rect 4342 55850 4398 56650
rect 4618 55850 4674 56650
rect 4894 55850 4950 56650
rect 5170 55850 5226 56650
rect 5446 55850 5502 56650
rect 5630 55850 5686 56650
rect 5906 55850 5962 56650
rect 6182 55850 6238 56650
rect 6458 55850 6514 56650
rect 6734 55850 6790 56650
rect 7010 55850 7066 56650
rect 7286 55850 7342 56650
rect 7562 55850 7618 56650
rect 7838 55850 7894 56650
rect 8114 55850 8170 56650
rect 8298 55850 8354 56650
rect 8574 55850 8630 56650
rect 8850 55850 8906 56650
rect 9126 55850 9182 56650
rect 9402 55850 9458 56650
rect 9678 55850 9734 56650
rect 9954 55850 10010 56650
rect 10230 55850 10286 56650
rect 10506 55850 10562 56650
rect 10782 55850 10838 56650
rect 10966 55850 11022 56650
rect 11242 55850 11298 56650
rect 11518 55850 11574 56650
rect 11794 55850 11850 56650
rect 12070 55850 12126 56650
rect 12346 55850 12402 56650
rect 12622 55850 12678 56650
rect 12898 55850 12954 56650
rect 13174 55850 13230 56650
rect 13450 55850 13506 56650
rect 13726 55850 13782 56650
rect 13910 55850 13966 56650
rect 14186 55850 14242 56650
rect 14462 55850 14518 56650
rect 14738 55850 14794 56650
rect 15014 55850 15070 56650
rect 15290 55850 15346 56650
rect 15566 55850 15622 56650
rect 15842 55850 15898 56650
rect 16118 55850 16174 56650
rect 16394 55850 16450 56650
rect 16578 55850 16634 56650
rect 16854 55850 16910 56650
rect 17130 55850 17186 56650
rect 17406 55850 17462 56650
rect 17682 55850 17738 56650
rect 17958 55850 18014 56650
rect 18234 55850 18290 56650
rect 18510 55850 18566 56650
rect 18786 55850 18842 56650
rect 19062 55850 19118 56650
rect 19246 55850 19302 56650
rect 19522 55850 19578 56650
rect 19798 55850 19854 56650
rect 20074 55850 20130 56650
rect 20350 55850 20406 56650
rect 20626 55850 20682 56650
rect 20902 55850 20958 56650
rect 21178 55850 21234 56650
rect 21454 55850 21510 56650
rect 21730 55850 21786 56650
rect 21914 55850 21970 56650
rect 22190 55850 22246 56650
rect 22466 55850 22522 56650
rect 22742 55850 22798 56650
rect 23018 55850 23074 56650
rect 23294 55850 23350 56650
rect 23570 55850 23626 56650
rect 23846 55850 23902 56650
rect 24122 55850 24178 56650
rect 24398 55850 24454 56650
rect 24582 55850 24638 56650
rect 24858 55850 24914 56650
rect 25134 55850 25190 56650
rect 25410 55850 25466 56650
rect 25686 55850 25742 56650
rect 25962 55850 26018 56650
rect 26238 55850 26294 56650
rect 26514 55850 26570 56650
rect 26790 55850 26846 56650
rect 27066 55850 27122 56650
rect 27342 55850 27398 56650
rect 27526 55850 27582 56650
rect 27802 55850 27858 56650
rect 28078 55850 28134 56650
rect 28354 55850 28410 56650
rect 28630 55850 28686 56650
rect 28906 55850 28962 56650
rect 29182 55850 29238 56650
rect 29458 55850 29514 56650
rect 29734 55850 29790 56650
rect 30010 55850 30066 56650
rect 30194 55850 30250 56650
rect 30470 55850 30526 56650
rect 30746 55850 30802 56650
rect 31022 55850 31078 56650
rect 31298 55850 31354 56650
rect 31574 55850 31630 56650
rect 31850 55850 31906 56650
rect 32126 55850 32182 56650
rect 32402 55850 32458 56650
rect 32678 55850 32734 56650
rect 32862 55850 32918 56650
rect 33138 55850 33194 56650
rect 33414 55850 33470 56650
rect 33690 55850 33746 56650
rect 33966 55850 34022 56650
rect 34242 55850 34298 56650
rect 34518 55850 34574 56650
rect 34794 55850 34850 56650
rect 35070 55850 35126 56650
rect 35346 55850 35402 56650
rect 35530 55850 35586 56650
rect 35806 55850 35862 56650
rect 36082 55850 36138 56650
rect 36358 55850 36414 56650
rect 36634 55850 36690 56650
rect 36910 55850 36966 56650
rect 37186 55850 37242 56650
rect 37462 55850 37518 56650
rect 37738 55850 37794 56650
rect 38014 55850 38070 56650
rect 38198 55850 38254 56650
rect 38474 55850 38530 56650
rect 38750 55850 38806 56650
rect 39026 55850 39082 56650
rect 39302 55850 39358 56650
rect 39578 55850 39634 56650
rect 39854 55850 39910 56650
rect 40130 55850 40186 56650
rect 40406 55850 40462 56650
rect 40682 55850 40738 56650
rect 40958 55850 41014 56650
rect 41142 55850 41198 56650
rect 41418 55850 41474 56650
rect 41694 55850 41750 56650
rect 41970 55850 42026 56650
rect 42246 55850 42302 56650
rect 42522 55850 42578 56650
rect 42798 55850 42854 56650
rect 43074 55850 43130 56650
rect 43350 55850 43406 56650
rect 43626 55850 43682 56650
rect 43810 55850 43866 56650
rect 44086 55850 44142 56650
rect 44362 55850 44418 56650
rect 44638 55850 44694 56650
rect 44914 55850 44970 56650
rect 45190 55850 45246 56650
rect 45466 55850 45522 56650
rect 45742 55850 45798 56650
rect 46018 55850 46074 56650
rect 46294 55850 46350 56650
rect 46478 55850 46534 56650
rect 46754 55850 46810 56650
rect 47030 55850 47086 56650
rect 47306 55850 47362 56650
rect 47582 55850 47638 56650
rect 47858 55850 47914 56650
rect 48134 55850 48190 56650
rect 48410 55850 48466 56650
rect 48686 55850 48742 56650
rect 48962 55850 49018 56650
rect 49146 55850 49202 56650
rect 49422 55850 49478 56650
rect 49698 55850 49754 56650
rect 49974 55850 50030 56650
rect 50250 55850 50306 56650
rect 50526 55850 50582 56650
rect 50802 55850 50858 56650
rect 51078 55850 51134 56650
rect 51354 55850 51410 56650
rect 51630 55850 51686 56650
rect 51814 55850 51870 56650
rect 52090 55850 52146 56650
rect 52366 55850 52422 56650
rect 52642 55850 52698 56650
rect 52918 55850 52974 56650
rect 53194 55850 53250 56650
rect 53470 55850 53526 56650
rect 53746 55850 53802 56650
rect 54022 55850 54078 56650
rect 54298 55850 54354 56650
rect 110 0 166 800
rect 294 0 350 800
rect 570 0 626 800
rect 846 0 902 800
rect 1122 0 1178 800
rect 1398 0 1454 800
rect 1674 0 1730 800
rect 1950 0 2006 800
rect 2226 0 2282 800
rect 2502 0 2558 800
rect 2778 0 2834 800
rect 2962 0 3018 800
rect 3238 0 3294 800
rect 3514 0 3570 800
rect 3790 0 3846 800
rect 4066 0 4122 800
rect 4342 0 4398 800
rect 4618 0 4674 800
rect 4894 0 4950 800
rect 5170 0 5226 800
rect 5446 0 5502 800
rect 5630 0 5686 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6458 0 6514 800
rect 6734 0 6790 800
rect 7010 0 7066 800
rect 7286 0 7342 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8298 0 8354 800
rect 8574 0 8630 800
rect 8850 0 8906 800
rect 9126 0 9182 800
rect 9402 0 9458 800
rect 9678 0 9734 800
rect 9954 0 10010 800
rect 10230 0 10286 800
rect 10506 0 10562 800
rect 10782 0 10838 800
rect 10966 0 11022 800
rect 11242 0 11298 800
rect 11518 0 11574 800
rect 11794 0 11850 800
rect 12070 0 12126 800
rect 12346 0 12402 800
rect 12622 0 12678 800
rect 12898 0 12954 800
rect 13174 0 13230 800
rect 13450 0 13506 800
rect 13726 0 13782 800
rect 13910 0 13966 800
rect 14186 0 14242 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15290 0 15346 800
rect 15566 0 15622 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16394 0 16450 800
rect 16578 0 16634 800
rect 16854 0 16910 800
rect 17130 0 17186 800
rect 17406 0 17462 800
rect 17682 0 17738 800
rect 17958 0 18014 800
rect 18234 0 18290 800
rect 18510 0 18566 800
rect 18786 0 18842 800
rect 19062 0 19118 800
rect 19246 0 19302 800
rect 19522 0 19578 800
rect 19798 0 19854 800
rect 20074 0 20130 800
rect 20350 0 20406 800
rect 20626 0 20682 800
rect 20902 0 20958 800
rect 21178 0 21234 800
rect 21454 0 21510 800
rect 21730 0 21786 800
rect 21914 0 21970 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23294 0 23350 800
rect 23570 0 23626 800
rect 23846 0 23902 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24582 0 24638 800
rect 24858 0 24914 800
rect 25134 0 25190 800
rect 25410 0 25466 800
rect 25686 0 25742 800
rect 25962 0 26018 800
rect 26238 0 26294 800
rect 26514 0 26570 800
rect 26790 0 26846 800
rect 27066 0 27122 800
rect 27342 0 27398 800
rect 27526 0 27582 800
rect 27802 0 27858 800
rect 28078 0 28134 800
rect 28354 0 28410 800
rect 28630 0 28686 800
rect 28906 0 28962 800
rect 29182 0 29238 800
rect 29458 0 29514 800
rect 29734 0 29790 800
rect 30010 0 30066 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32678 0 32734 800
rect 32862 0 32918 800
rect 33138 0 33194 800
rect 33414 0 33470 800
rect 33690 0 33746 800
rect 33966 0 34022 800
rect 34242 0 34298 800
rect 34518 0 34574 800
rect 34794 0 34850 800
rect 35070 0 35126 800
rect 35346 0 35402 800
rect 35530 0 35586 800
rect 35806 0 35862 800
rect 36082 0 36138 800
rect 36358 0 36414 800
rect 36634 0 36690 800
rect 36910 0 36966 800
rect 37186 0 37242 800
rect 37462 0 37518 800
rect 37738 0 37794 800
rect 38014 0 38070 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38750 0 38806 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39578 0 39634 800
rect 39854 0 39910 800
rect 40130 0 40186 800
rect 40406 0 40462 800
rect 40682 0 40738 800
rect 40958 0 41014 800
rect 41142 0 41198 800
rect 41418 0 41474 800
rect 41694 0 41750 800
rect 41970 0 42026 800
rect 42246 0 42302 800
rect 42522 0 42578 800
rect 42798 0 42854 800
rect 43074 0 43130 800
rect 43350 0 43406 800
rect 43626 0 43682 800
rect 43810 0 43866 800
rect 44086 0 44142 800
rect 44362 0 44418 800
rect 44638 0 44694 800
rect 44914 0 44970 800
rect 45190 0 45246 800
rect 45466 0 45522 800
rect 45742 0 45798 800
rect 46018 0 46074 800
rect 46294 0 46350 800
rect 46478 0 46534 800
rect 46754 0 46810 800
rect 47030 0 47086 800
rect 47306 0 47362 800
rect 47582 0 47638 800
rect 47858 0 47914 800
rect 48134 0 48190 800
rect 48410 0 48466 800
rect 48686 0 48742 800
rect 48962 0 49018 800
rect 49146 0 49202 800
rect 49422 0 49478 800
rect 49698 0 49754 800
rect 49974 0 50030 800
rect 50250 0 50306 800
rect 50526 0 50582 800
rect 50802 0 50858 800
rect 51078 0 51134 800
rect 51354 0 51410 800
rect 51630 0 51686 800
rect 51814 0 51870 800
rect 52090 0 52146 800
rect 52366 0 52422 800
rect 52642 0 52698 800
rect 52918 0 52974 800
rect 53194 0 53250 800
rect 53470 0 53526 800
rect 53746 0 53802 800
rect 54022 0 54078 800
rect 54298 0 54354 800
<< obsm2 >>
rect 222 55794 238 56545
rect 406 55794 514 56545
rect 682 55794 790 56545
rect 958 55794 1066 56545
rect 1234 55794 1342 56545
rect 1510 55794 1618 56545
rect 1786 55794 1894 56545
rect 2062 55794 2170 56545
rect 2338 55794 2446 56545
rect 2614 55794 2722 56545
rect 2890 55794 2906 56545
rect 3074 55794 3182 56545
rect 3350 55794 3458 56545
rect 3626 55794 3734 56545
rect 3902 55794 4010 56545
rect 4178 55794 4286 56545
rect 4454 55794 4562 56545
rect 4730 55794 4838 56545
rect 5006 55794 5114 56545
rect 5282 55794 5390 56545
rect 5558 55794 5574 56545
rect 5742 55794 5850 56545
rect 6018 55794 6126 56545
rect 6294 55794 6402 56545
rect 6570 55794 6678 56545
rect 6846 55794 6954 56545
rect 7122 55794 7230 56545
rect 7398 55794 7506 56545
rect 7674 55794 7782 56545
rect 7950 55794 8058 56545
rect 8226 55794 8242 56545
rect 8410 55794 8518 56545
rect 8686 55794 8794 56545
rect 8962 55794 9070 56545
rect 9238 55794 9346 56545
rect 9514 55794 9622 56545
rect 9790 55794 9898 56545
rect 10066 55794 10174 56545
rect 10342 55794 10450 56545
rect 10618 55794 10726 56545
rect 10894 55794 10910 56545
rect 11078 55794 11186 56545
rect 11354 55794 11462 56545
rect 11630 55794 11738 56545
rect 11906 55794 12014 56545
rect 12182 55794 12290 56545
rect 12458 55794 12566 56545
rect 12734 55794 12842 56545
rect 13010 55794 13118 56545
rect 13286 55794 13394 56545
rect 13562 55794 13670 56545
rect 13838 55794 13854 56545
rect 14022 55794 14130 56545
rect 14298 55794 14406 56545
rect 14574 55794 14682 56545
rect 14850 55794 14958 56545
rect 15126 55794 15234 56545
rect 15402 55794 15510 56545
rect 15678 55794 15786 56545
rect 15954 55794 16062 56545
rect 16230 55794 16338 56545
rect 16506 55794 16522 56545
rect 16690 55794 16798 56545
rect 16966 55794 17074 56545
rect 17242 55794 17350 56545
rect 17518 55794 17626 56545
rect 17794 55794 17902 56545
rect 18070 55794 18178 56545
rect 18346 55794 18454 56545
rect 18622 55794 18730 56545
rect 18898 55794 19006 56545
rect 19174 55794 19190 56545
rect 19358 55794 19466 56545
rect 19634 55794 19742 56545
rect 19910 55794 20018 56545
rect 20186 55794 20294 56545
rect 20462 55794 20570 56545
rect 20738 55794 20846 56545
rect 21014 55794 21122 56545
rect 21290 55794 21398 56545
rect 21566 55794 21674 56545
rect 21842 55794 21858 56545
rect 22026 55794 22134 56545
rect 22302 55794 22410 56545
rect 22578 55794 22686 56545
rect 22854 55794 22962 56545
rect 23130 55794 23238 56545
rect 23406 55794 23514 56545
rect 23682 55794 23790 56545
rect 23958 55794 24066 56545
rect 24234 55794 24342 56545
rect 24510 55794 24526 56545
rect 24694 55794 24802 56545
rect 24970 55794 25078 56545
rect 25246 55794 25354 56545
rect 25522 55794 25630 56545
rect 25798 55794 25906 56545
rect 26074 55794 26182 56545
rect 26350 55794 26458 56545
rect 26626 55794 26734 56545
rect 26902 55794 27010 56545
rect 27178 55794 27286 56545
rect 27454 55794 27470 56545
rect 27638 55794 27746 56545
rect 27914 55794 28022 56545
rect 28190 55794 28298 56545
rect 28466 55794 28574 56545
rect 28742 55794 28850 56545
rect 29018 55794 29126 56545
rect 29294 55794 29402 56545
rect 29570 55794 29678 56545
rect 29846 55794 29954 56545
rect 30122 55794 30138 56545
rect 30306 55794 30414 56545
rect 30582 55794 30690 56545
rect 30858 55794 30966 56545
rect 31134 55794 31242 56545
rect 31410 55794 31518 56545
rect 31686 55794 31794 56545
rect 31962 55794 32070 56545
rect 32238 55794 32346 56545
rect 32514 55794 32622 56545
rect 32790 55794 32806 56545
rect 32974 55794 33082 56545
rect 33250 55794 33358 56545
rect 33526 55794 33634 56545
rect 33802 55794 33910 56545
rect 34078 55794 34186 56545
rect 34354 55794 34462 56545
rect 34630 55794 34738 56545
rect 34906 55794 35014 56545
rect 35182 55794 35290 56545
rect 35458 55794 35474 56545
rect 35642 55794 35750 56545
rect 35918 55794 36026 56545
rect 36194 55794 36302 56545
rect 36470 55794 36578 56545
rect 36746 55794 36854 56545
rect 37022 55794 37130 56545
rect 37298 55794 37406 56545
rect 37574 55794 37682 56545
rect 37850 55794 37958 56545
rect 38126 55794 38142 56545
rect 38310 55794 38418 56545
rect 38586 55794 38694 56545
rect 38862 55794 38970 56545
rect 39138 55794 39246 56545
rect 39414 55794 39522 56545
rect 39690 55794 39798 56545
rect 39966 55794 40074 56545
rect 40242 55794 40350 56545
rect 40518 55794 40626 56545
rect 40794 55794 40902 56545
rect 41070 55794 41086 56545
rect 41254 55794 41362 56545
rect 41530 55794 41638 56545
rect 41806 55794 41914 56545
rect 42082 55794 42190 56545
rect 42358 55794 42466 56545
rect 42634 55794 42742 56545
rect 42910 55794 43018 56545
rect 43186 55794 43294 56545
rect 43462 55794 43570 56545
rect 43738 55794 43754 56545
rect 43922 55794 44030 56545
rect 44198 55794 44306 56545
rect 44474 55794 44582 56545
rect 44750 55794 44858 56545
rect 45026 55794 45134 56545
rect 45302 55794 45410 56545
rect 45578 55794 45686 56545
rect 45854 55794 45962 56545
rect 46130 55794 46238 56545
rect 46406 55794 46422 56545
rect 46590 55794 46698 56545
rect 46866 55794 46974 56545
rect 47142 55794 47250 56545
rect 47418 55794 47526 56545
rect 47694 55794 47802 56545
rect 47970 55794 48078 56545
rect 48246 55794 48354 56545
rect 48522 55794 48630 56545
rect 48798 55794 48906 56545
rect 49074 55794 49090 56545
rect 49258 55794 49366 56545
rect 49534 55794 49642 56545
rect 49810 55794 49918 56545
rect 50086 55794 50194 56545
rect 50362 55794 50470 56545
rect 50638 55794 50746 56545
rect 50914 55794 51022 56545
rect 51190 55794 51298 56545
rect 51466 55794 51574 56545
rect 51742 55794 51758 56545
rect 51926 55794 52034 56545
rect 52202 55794 52310 56545
rect 52478 55794 52586 56545
rect 52754 55794 52862 56545
rect 53030 55794 53138 56545
rect 53306 55794 53414 56545
rect 53582 55794 53690 56545
rect 53858 55794 53966 56545
rect 54134 55794 54242 56545
rect 54410 55794 54444 56545
rect 112 856 54444 55794
rect 222 2 238 856
rect 406 2 514 856
rect 682 2 790 856
rect 958 2 1066 856
rect 1234 2 1342 856
rect 1510 2 1618 856
rect 1786 2 1894 856
rect 2062 2 2170 856
rect 2338 2 2446 856
rect 2614 2 2722 856
rect 2890 2 2906 856
rect 3074 2 3182 856
rect 3350 2 3458 856
rect 3626 2 3734 856
rect 3902 2 4010 856
rect 4178 2 4286 856
rect 4454 2 4562 856
rect 4730 2 4838 856
rect 5006 2 5114 856
rect 5282 2 5390 856
rect 5558 2 5574 856
rect 5742 2 5850 856
rect 6018 2 6126 856
rect 6294 2 6402 856
rect 6570 2 6678 856
rect 6846 2 6954 856
rect 7122 2 7230 856
rect 7398 2 7506 856
rect 7674 2 7782 856
rect 7950 2 8058 856
rect 8226 2 8242 856
rect 8410 2 8518 856
rect 8686 2 8794 856
rect 8962 2 9070 856
rect 9238 2 9346 856
rect 9514 2 9622 856
rect 9790 2 9898 856
rect 10066 2 10174 856
rect 10342 2 10450 856
rect 10618 2 10726 856
rect 10894 2 10910 856
rect 11078 2 11186 856
rect 11354 2 11462 856
rect 11630 2 11738 856
rect 11906 2 12014 856
rect 12182 2 12290 856
rect 12458 2 12566 856
rect 12734 2 12842 856
rect 13010 2 13118 856
rect 13286 2 13394 856
rect 13562 2 13670 856
rect 13838 2 13854 856
rect 14022 2 14130 856
rect 14298 2 14406 856
rect 14574 2 14682 856
rect 14850 2 14958 856
rect 15126 2 15234 856
rect 15402 2 15510 856
rect 15678 2 15786 856
rect 15954 2 16062 856
rect 16230 2 16338 856
rect 16506 2 16522 856
rect 16690 2 16798 856
rect 16966 2 17074 856
rect 17242 2 17350 856
rect 17518 2 17626 856
rect 17794 2 17902 856
rect 18070 2 18178 856
rect 18346 2 18454 856
rect 18622 2 18730 856
rect 18898 2 19006 856
rect 19174 2 19190 856
rect 19358 2 19466 856
rect 19634 2 19742 856
rect 19910 2 20018 856
rect 20186 2 20294 856
rect 20462 2 20570 856
rect 20738 2 20846 856
rect 21014 2 21122 856
rect 21290 2 21398 856
rect 21566 2 21674 856
rect 21842 2 21858 856
rect 22026 2 22134 856
rect 22302 2 22410 856
rect 22578 2 22686 856
rect 22854 2 22962 856
rect 23130 2 23238 856
rect 23406 2 23514 856
rect 23682 2 23790 856
rect 23958 2 24066 856
rect 24234 2 24342 856
rect 24510 2 24526 856
rect 24694 2 24802 856
rect 24970 2 25078 856
rect 25246 2 25354 856
rect 25522 2 25630 856
rect 25798 2 25906 856
rect 26074 2 26182 856
rect 26350 2 26458 856
rect 26626 2 26734 856
rect 26902 2 27010 856
rect 27178 2 27286 856
rect 27454 2 27470 856
rect 27638 2 27746 856
rect 27914 2 28022 856
rect 28190 2 28298 856
rect 28466 2 28574 856
rect 28742 2 28850 856
rect 29018 2 29126 856
rect 29294 2 29402 856
rect 29570 2 29678 856
rect 29846 2 29954 856
rect 30122 2 30138 856
rect 30306 2 30414 856
rect 30582 2 30690 856
rect 30858 2 30966 856
rect 31134 2 31242 856
rect 31410 2 31518 856
rect 31686 2 31794 856
rect 31962 2 32070 856
rect 32238 2 32346 856
rect 32514 2 32622 856
rect 32790 2 32806 856
rect 32974 2 33082 856
rect 33250 2 33358 856
rect 33526 2 33634 856
rect 33802 2 33910 856
rect 34078 2 34186 856
rect 34354 2 34462 856
rect 34630 2 34738 856
rect 34906 2 35014 856
rect 35182 2 35290 856
rect 35458 2 35474 856
rect 35642 2 35750 856
rect 35918 2 36026 856
rect 36194 2 36302 856
rect 36470 2 36578 856
rect 36746 2 36854 856
rect 37022 2 37130 856
rect 37298 2 37406 856
rect 37574 2 37682 856
rect 37850 2 37958 856
rect 38126 2 38142 856
rect 38310 2 38418 856
rect 38586 2 38694 856
rect 38862 2 38970 856
rect 39138 2 39246 856
rect 39414 2 39522 856
rect 39690 2 39798 856
rect 39966 2 40074 856
rect 40242 2 40350 856
rect 40518 2 40626 856
rect 40794 2 40902 856
rect 41070 2 41086 856
rect 41254 2 41362 856
rect 41530 2 41638 856
rect 41806 2 41914 856
rect 42082 2 42190 856
rect 42358 2 42466 856
rect 42634 2 42742 856
rect 42910 2 43018 856
rect 43186 2 43294 856
rect 43462 2 43570 856
rect 43738 2 43754 856
rect 43922 2 44030 856
rect 44198 2 44306 856
rect 44474 2 44582 856
rect 44750 2 44858 856
rect 45026 2 45134 856
rect 45302 2 45410 856
rect 45578 2 45686 856
rect 45854 2 45962 856
rect 46130 2 46238 856
rect 46406 2 46422 856
rect 46590 2 46698 856
rect 46866 2 46974 856
rect 47142 2 47250 856
rect 47418 2 47526 856
rect 47694 2 47802 856
rect 47970 2 48078 856
rect 48246 2 48354 856
rect 48522 2 48630 856
rect 48798 2 48906 856
rect 49074 2 49090 856
rect 49258 2 49366 856
rect 49534 2 49642 856
rect 49810 2 49918 856
rect 50086 2 50194 856
rect 50362 2 50470 856
rect 50638 2 50746 856
rect 50914 2 51022 856
rect 51190 2 51298 856
rect 51466 2 51574 856
rect 51742 2 51758 856
rect 51926 2 52034 856
rect 52202 2 52310 856
rect 52478 2 52586 856
rect 52754 2 52862 856
rect 53030 2 53138 856
rect 53306 2 53414 856
rect 53582 2 53690 856
rect 53858 2 53966 856
rect 54134 2 54242 856
rect 54410 2 54444 856
<< metal3 >>
rect 53706 56448 54506 56568
rect 53706 56176 54506 56296
rect 53706 55904 54506 56024
rect 53706 55632 54506 55752
rect 53706 55360 54506 55480
rect 53706 55088 54506 55208
rect 53706 54816 54506 54936
rect 53706 54544 54506 54664
rect 53706 54272 54506 54392
rect 53706 54000 54506 54120
rect 53706 53728 54506 53848
rect 53706 53456 54506 53576
rect 53706 53184 54506 53304
rect 53706 52912 54506 53032
rect 53706 52640 54506 52760
rect 53706 52368 54506 52488
rect 53706 52096 54506 52216
rect 53706 51824 54506 51944
rect 53706 51552 54506 51672
rect 53706 51280 54506 51400
rect 53706 51008 54506 51128
rect 53706 50736 54506 50856
rect 53706 50328 54506 50448
rect 53706 50056 54506 50176
rect 53706 49784 54506 49904
rect 53706 49512 54506 49632
rect 53706 49240 54506 49360
rect 53706 48968 54506 49088
rect 53706 48696 54506 48816
rect 53706 48424 54506 48544
rect 53706 48152 54506 48272
rect 53706 47880 54506 48000
rect 53706 47608 54506 47728
rect 53706 47336 54506 47456
rect 53706 47064 54506 47184
rect 53706 46792 54506 46912
rect 53706 46520 54506 46640
rect 53706 46248 54506 46368
rect 53706 45976 54506 46096
rect 53706 45704 54506 45824
rect 53706 45432 54506 45552
rect 53706 45160 54506 45280
rect 53706 44888 54506 45008
rect 53706 44616 54506 44736
rect 53706 44344 54506 44464
rect 53706 43936 54506 44056
rect 53706 43664 54506 43784
rect 53706 43392 54506 43512
rect 53706 43120 54506 43240
rect 53706 42848 54506 42968
rect 0 42440 800 42560
rect 53706 42576 54506 42696
rect 53706 42304 54506 42424
rect 53706 42032 54506 42152
rect 53706 41760 54506 41880
rect 53706 41488 54506 41608
rect 53706 41216 54506 41336
rect 53706 40944 54506 41064
rect 53706 40672 54506 40792
rect 53706 40400 54506 40520
rect 53706 40128 54506 40248
rect 53706 39856 54506 39976
rect 53706 39584 54506 39704
rect 53706 39312 54506 39432
rect 53706 39040 54506 39160
rect 53706 38768 54506 38888
rect 53706 38496 54506 38616
rect 53706 38224 54506 38344
rect 53706 37952 54506 38072
rect 53706 37544 54506 37664
rect 53706 37272 54506 37392
rect 53706 37000 54506 37120
rect 53706 36728 54506 36848
rect 53706 36456 54506 36576
rect 53706 36184 54506 36304
rect 53706 35912 54506 36032
rect 53706 35640 54506 35760
rect 53706 35368 54506 35488
rect 53706 35096 54506 35216
rect 53706 34824 54506 34944
rect 53706 34552 54506 34672
rect 53706 34280 54506 34400
rect 53706 34008 54506 34128
rect 53706 33736 54506 33856
rect 53706 33464 54506 33584
rect 53706 33192 54506 33312
rect 53706 32920 54506 33040
rect 53706 32648 54506 32768
rect 53706 32376 54506 32496
rect 53706 32104 54506 32224
rect 53706 31832 54506 31952
rect 53706 31424 54506 31544
rect 53706 31152 54506 31272
rect 53706 30880 54506 31000
rect 53706 30608 54506 30728
rect 53706 30336 54506 30456
rect 53706 30064 54506 30184
rect 53706 29792 54506 29912
rect 53706 29520 54506 29640
rect 53706 29248 54506 29368
rect 53706 28976 54506 29096
rect 53706 28704 54506 28824
rect 53706 28432 54506 28552
rect 53706 28160 54506 28280
rect 53706 27888 54506 28008
rect 53706 27616 54506 27736
rect 53706 27344 54506 27464
rect 53706 27072 54506 27192
rect 53706 26800 54506 26920
rect 53706 26528 54506 26648
rect 53706 26256 54506 26376
rect 53706 25984 54506 26104
rect 53706 25712 54506 25832
rect 53706 25440 54506 25560
rect 53706 25032 54506 25152
rect 53706 24760 54506 24880
rect 53706 24488 54506 24608
rect 53706 24216 54506 24336
rect 53706 23944 54506 24064
rect 53706 23672 54506 23792
rect 53706 23400 54506 23520
rect 53706 23128 54506 23248
rect 53706 22856 54506 22976
rect 53706 22584 54506 22704
rect 53706 22312 54506 22432
rect 53706 22040 54506 22160
rect 53706 21768 54506 21888
rect 53706 21496 54506 21616
rect 53706 21224 54506 21344
rect 53706 20952 54506 21072
rect 53706 20680 54506 20800
rect 53706 20408 54506 20528
rect 53706 20136 54506 20256
rect 53706 19864 54506 19984
rect 53706 19592 54506 19712
rect 53706 19320 54506 19440
rect 53706 19048 54506 19168
rect 53706 18640 54506 18760
rect 53706 18368 54506 18488
rect 53706 18096 54506 18216
rect 53706 17824 54506 17944
rect 53706 17552 54506 17672
rect 53706 17280 54506 17400
rect 53706 17008 54506 17128
rect 53706 16736 54506 16856
rect 53706 16464 54506 16584
rect 53706 16192 54506 16312
rect 53706 15920 54506 16040
rect 53706 15648 54506 15768
rect 53706 15376 54506 15496
rect 53706 15104 54506 15224
rect 53706 14832 54506 14952
rect 53706 14560 54506 14680
rect 0 14152 800 14272
rect 53706 14288 54506 14408
rect 53706 14016 54506 14136
rect 53706 13744 54506 13864
rect 53706 13472 54506 13592
rect 53706 13200 54506 13320
rect 53706 12928 54506 13048
rect 53706 12520 54506 12640
rect 53706 12248 54506 12368
rect 53706 11976 54506 12096
rect 53706 11704 54506 11824
rect 53706 11432 54506 11552
rect 53706 11160 54506 11280
rect 53706 10888 54506 11008
rect 53706 10616 54506 10736
rect 53706 10344 54506 10464
rect 53706 10072 54506 10192
rect 53706 9800 54506 9920
rect 53706 9528 54506 9648
rect 53706 9256 54506 9376
rect 53706 8984 54506 9104
rect 53706 8712 54506 8832
rect 53706 8440 54506 8560
rect 53706 8168 54506 8288
rect 53706 7896 54506 8016
rect 53706 7624 54506 7744
rect 53706 7352 54506 7472
rect 53706 7080 54506 7200
rect 53706 6808 54506 6928
rect 53706 6536 54506 6656
rect 53706 6128 54506 6248
rect 53706 5856 54506 5976
rect 53706 5584 54506 5704
rect 53706 5312 54506 5432
rect 53706 5040 54506 5160
rect 53706 4768 54506 4888
rect 53706 4496 54506 4616
rect 53706 4224 54506 4344
rect 53706 3952 54506 4072
rect 53706 3680 54506 3800
rect 53706 3408 54506 3528
rect 53706 3136 54506 3256
rect 53706 2864 54506 2984
rect 53706 2592 54506 2712
rect 53706 2320 54506 2440
rect 53706 2048 54506 2168
rect 53706 1776 54506 1896
rect 53706 1504 54506 1624
rect 53706 1232 54506 1352
rect 53706 960 54506 1080
rect 53706 688 54506 808
rect 53706 416 54506 536
rect 53706 144 54506 264
<< obsm3 >>
rect 790 50656 53626 56541
rect 790 50528 53706 50656
rect 790 44264 53626 50528
rect 790 44136 53706 44264
rect 790 42640 53626 44136
rect 880 42360 53626 42640
rect 790 37872 53626 42360
rect 790 37744 53706 37872
rect 790 31752 53626 37744
rect 790 31624 53706 31752
rect 790 25360 53626 31624
rect 790 25232 53706 25360
rect 790 18968 53626 25232
rect 790 18840 53706 18968
rect 790 14352 53626 18840
rect 880 14072 53626 14352
rect 790 12848 53626 14072
rect 790 12720 53706 12848
rect 790 6456 53626 12720
rect 790 6328 53706 6456
rect 790 64 53626 6328
rect 790 35 53706 64
<< metal4 >>
rect 4208 2128 4528 54448
rect 19568 2128 19888 54448
rect 34928 2128 35248 54448
rect 50288 2128 50608 54448
<< obsm4 >>
rect 795 54528 52749 56269
rect 795 2048 4128 54528
rect 4608 2048 19488 54528
rect 19968 2048 34848 54528
rect 35328 2048 50208 54528
rect 50688 2048 52749 54528
rect 795 35 52749 2048
<< labels >>
rlabel metal3 s 0 14152 800 14272 6 CLK
port 1 nsew signal input
rlabel metal2 s 110 0 166 800 6 EN_core_dmem_request_put
port 2 nsew signal input
rlabel metal2 s 294 0 350 800 6 EN_core_dmem_response_get
port 3 nsew signal input
rlabel metal2 s 570 0 626 800 6 EN_core_imem_request_put
port 4 nsew signal input
rlabel metal2 s 846 0 902 800 6 EN_core_imem_response_get
port 5 nsew signal input
rlabel metal3 s 53706 144 54506 264 6 EN_fmc_dmem_request_get
port 6 nsew signal input
rlabel metal3 s 53706 416 54506 536 6 EN_fmc_dmem_response_put
port 7 nsew signal input
rlabel metal3 s 53706 688 54506 808 6 EN_fmc_imem_request_get
port 8 nsew signal input
rlabel metal3 s 53706 960 54506 1080 6 EN_fmc_imem_response_put
port 9 nsew signal input
rlabel metal2 s 110 55850 166 56650 6 EN_ram_dmem_request_get
port 10 nsew signal input
rlabel metal2 s 294 55850 350 56650 6 EN_ram_dmem_response_put
port 11 nsew signal input
rlabel metal2 s 570 55850 626 56650 6 EN_ram_imem_request_get
port 12 nsew signal input
rlabel metal2 s 846 55850 902 56650 6 EN_ram_imem_response_put
port 13 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 RDY_core_dmem_request_put
port 14 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 RDY_core_dmem_response_get
port 15 nsew signal output
rlabel metal2 s 1674 0 1730 800 6 RDY_core_imem_request_put
port 16 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 RDY_core_imem_response_get
port 17 nsew signal output
rlabel metal3 s 53706 1232 54506 1352 6 RDY_fmc_dmem_request_get
port 18 nsew signal output
rlabel metal3 s 53706 1504 54506 1624 6 RDY_fmc_dmem_response_put
port 19 nsew signal output
rlabel metal3 s 53706 1776 54506 1896 6 RDY_fmc_imem_request_get
port 20 nsew signal output
rlabel metal3 s 53706 2048 54506 2168 6 RDY_fmc_imem_response_put
port 21 nsew signal output
rlabel metal2 s 1122 55850 1178 56650 6 RDY_ram_dmem_request_get
port 22 nsew signal output
rlabel metal2 s 1398 55850 1454 56650 6 RDY_ram_dmem_response_put
port 23 nsew signal output
rlabel metal2 s 1674 55850 1730 56650 6 RDY_ram_imem_request_get
port 24 nsew signal output
rlabel metal2 s 1950 55850 2006 56650 6 RDY_ram_imem_response_put
port 25 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 RST_N
port 26 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 core_dmem_request_put[0]
port 27 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 core_dmem_request_put[10]
port 28 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 core_dmem_request_put[11]
port 29 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 core_dmem_request_put[12]
port 30 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 core_dmem_request_put[13]
port 31 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 core_dmem_request_put[14]
port 32 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 core_dmem_request_put[15]
port 33 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 core_dmem_request_put[16]
port 34 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 core_dmem_request_put[17]
port 35 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 core_dmem_request_put[18]
port 36 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 core_dmem_request_put[19]
port 37 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 core_dmem_request_put[1]
port 38 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 core_dmem_request_put[20]
port 39 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 core_dmem_request_put[21]
port 40 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 core_dmem_request_put[22]
port 41 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 core_dmem_request_put[23]
port 42 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 core_dmem_request_put[24]
port 43 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 core_dmem_request_put[25]
port 44 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 core_dmem_request_put[26]
port 45 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 core_dmem_request_put[27]
port 46 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 core_dmem_request_put[28]
port 47 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 core_dmem_request_put[29]
port 48 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 core_dmem_request_put[2]
port 49 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 core_dmem_request_put[30]
port 50 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 core_dmem_request_put[31]
port 51 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 core_dmem_request_put[32]
port 52 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 core_dmem_request_put[33]
port 53 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 core_dmem_request_put[34]
port 54 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 core_dmem_request_put[35]
port 55 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 core_dmem_request_put[36]
port 56 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 core_dmem_request_put[37]
port 57 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 core_dmem_request_put[38]
port 58 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 core_dmem_request_put[39]
port 59 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 core_dmem_request_put[3]
port 60 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 core_dmem_request_put[40]
port 61 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 core_dmem_request_put[41]
port 62 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 core_dmem_request_put[42]
port 63 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 core_dmem_request_put[43]
port 64 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 core_dmem_request_put[44]
port 65 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 core_dmem_request_put[45]
port 66 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 core_dmem_request_put[46]
port 67 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 core_dmem_request_put[47]
port 68 nsew signal input
rlabel metal2 s 40682 0 40738 800 6 core_dmem_request_put[48]
port 69 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 core_dmem_request_put[49]
port 70 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 core_dmem_request_put[4]
port 71 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 core_dmem_request_put[50]
port 72 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 core_dmem_request_put[51]
port 73 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 core_dmem_request_put[52]
port 74 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 core_dmem_request_put[53]
port 75 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 core_dmem_request_put[54]
port 76 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 core_dmem_request_put[55]
port 77 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 core_dmem_request_put[56]
port 78 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 core_dmem_request_put[57]
port 79 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 core_dmem_request_put[58]
port 80 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 core_dmem_request_put[59]
port 81 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 core_dmem_request_put[5]
port 82 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 core_dmem_request_put[60]
port 83 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 core_dmem_request_put[61]
port 84 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 core_dmem_request_put[62]
port 85 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 core_dmem_request_put[63]
port 86 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 core_dmem_request_put[64]
port 87 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 core_dmem_request_put[65]
port 88 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 core_dmem_request_put[66]
port 89 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 core_dmem_request_put[67]
port 90 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 core_dmem_request_put[68]
port 91 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 core_dmem_request_put[69]
port 92 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 core_dmem_request_put[6]
port 93 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 core_dmem_request_put[70]
port 94 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 core_dmem_request_put[71]
port 95 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 core_dmem_request_put[72]
port 96 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 core_dmem_request_put[73]
port 97 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 core_dmem_request_put[74]
port 98 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 core_dmem_request_put[75]
port 99 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 core_dmem_request_put[76]
port 100 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 core_dmem_request_put[77]
port 101 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 core_dmem_request_put[78]
port 102 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 core_dmem_request_put[79]
port 103 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 core_dmem_request_put[7]
port 104 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 core_dmem_request_put[80]
port 105 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 core_dmem_request_put[81]
port 106 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 core_dmem_request_put[82]
port 107 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 core_dmem_request_put[83]
port 108 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 core_dmem_request_put[84]
port 109 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 core_dmem_request_put[85]
port 110 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 core_dmem_request_put[86]
port 111 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 core_dmem_request_put[87]
port 112 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 core_dmem_request_put[88]
port 113 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 core_dmem_request_put[89]
port 114 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 core_dmem_request_put[8]
port 115 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 core_dmem_request_put[90]
port 116 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 core_dmem_request_put[91]
port 117 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 core_dmem_request_put[92]
port 118 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 core_dmem_request_put[93]
port 119 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 core_dmem_request_put[94]
port 120 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 core_dmem_request_put[95]
port 121 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 core_dmem_request_put[96]
port 122 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 core_dmem_request_put[97]
port 123 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 core_dmem_request_put[98]
port 124 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 core_dmem_request_put[99]
port 125 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 core_dmem_request_put[9]
port 126 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 core_dmem_response_get[0]
port 127 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 core_dmem_response_get[10]
port 128 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 core_dmem_response_get[11]
port 129 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 core_dmem_response_get[12]
port 130 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 core_dmem_response_get[13]
port 131 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 core_dmem_response_get[14]
port 132 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 core_dmem_response_get[15]
port 133 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 core_dmem_response_get[16]
port 134 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 core_dmem_response_get[17]
port 135 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 core_dmem_response_get[18]
port 136 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 core_dmem_response_get[19]
port 137 nsew signal output
rlabel metal2 s 3514 0 3570 800 6 core_dmem_response_get[1]
port 138 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 core_dmem_response_get[20]
port 139 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 core_dmem_response_get[21]
port 140 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 core_dmem_response_get[22]
port 141 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 core_dmem_response_get[23]
port 142 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 core_dmem_response_get[24]
port 143 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 core_dmem_response_get[25]
port 144 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 core_dmem_response_get[26]
port 145 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 core_dmem_response_get[27]
port 146 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 core_dmem_response_get[28]
port 147 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 core_dmem_response_get[29]
port 148 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 core_dmem_response_get[2]
port 149 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 core_dmem_response_get[30]
port 150 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 core_dmem_response_get[31]
port 151 nsew signal output
rlabel metal2 s 5630 0 5686 800 6 core_dmem_response_get[3]
port 152 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 core_dmem_response_get[4]
port 153 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 core_dmem_response_get[5]
port 154 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 core_dmem_response_get[6]
port 155 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 core_dmem_response_get[7]
port 156 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 core_dmem_response_get[8]
port 157 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 core_dmem_response_get[9]
port 158 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 core_imem_request_put[0]
port 159 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 core_imem_request_put[10]
port 160 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 core_imem_request_put[11]
port 161 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 core_imem_request_put[12]
port 162 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 core_imem_request_put[13]
port 163 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 core_imem_request_put[14]
port 164 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 core_imem_request_put[15]
port 165 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 core_imem_request_put[16]
port 166 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 core_imem_request_put[17]
port 167 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 core_imem_request_put[18]
port 168 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 core_imem_request_put[19]
port 169 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 core_imem_request_put[1]
port 170 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 core_imem_request_put[20]
port 171 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 core_imem_request_put[21]
port 172 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 core_imem_request_put[22]
port 173 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 core_imem_request_put[23]
port 174 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 core_imem_request_put[24]
port 175 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 core_imem_request_put[25]
port 176 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 core_imem_request_put[26]
port 177 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 core_imem_request_put[27]
port 178 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 core_imem_request_put[28]
port 179 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 core_imem_request_put[29]
port 180 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 core_imem_request_put[2]
port 181 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 core_imem_request_put[30]
port 182 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 core_imem_request_put[31]
port 183 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 core_imem_request_put[3]
port 184 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 core_imem_request_put[4]
port 185 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 core_imem_request_put[5]
port 186 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 core_imem_request_put[6]
port 187 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 core_imem_request_put[7]
port 188 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 core_imem_request_put[8]
port 189 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 core_imem_request_put[9]
port 190 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 core_imem_response_get[0]
port 191 nsew signal output
rlabel metal2 s 13726 0 13782 800 6 core_imem_response_get[10]
port 192 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 core_imem_response_get[11]
port 193 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 core_imem_response_get[12]
port 194 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 core_imem_response_get[13]
port 195 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 core_imem_response_get[14]
port 196 nsew signal output
rlabel metal2 s 19062 0 19118 800 6 core_imem_response_get[15]
port 197 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 core_imem_response_get[16]
port 198 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 core_imem_response_get[17]
port 199 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 core_imem_response_get[18]
port 200 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 core_imem_response_get[19]
port 201 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 core_imem_response_get[1]
port 202 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 core_imem_response_get[20]
port 203 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 core_imem_response_get[21]
port 204 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 core_imem_response_get[22]
port 205 nsew signal output
rlabel metal2 s 27526 0 27582 800 6 core_imem_response_get[23]
port 206 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 core_imem_response_get[24]
port 207 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 core_imem_response_get[25]
port 208 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 core_imem_response_get[26]
port 209 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 core_imem_response_get[27]
port 210 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 core_imem_response_get[28]
port 211 nsew signal output
rlabel metal2 s 33966 0 34022 800 6 core_imem_response_get[29]
port 212 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 core_imem_response_get[2]
port 213 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 core_imem_response_get[30]
port 214 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 core_imem_response_get[31]
port 215 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 core_imem_response_get[3]
port 216 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 core_imem_response_get[4]
port 217 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 core_imem_response_get[5]
port 218 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 core_imem_response_get[6]
port 219 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 core_imem_response_get[7]
port 220 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 core_imem_response_get[8]
port 221 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 core_imem_response_get[9]
port 222 nsew signal output
rlabel metal3 s 53706 2320 54506 2440 6 fmc_dmem_request_get[0]
port 223 nsew signal output
rlabel metal3 s 53706 13472 54506 13592 6 fmc_dmem_request_get[10]
port 224 nsew signal output
rlabel metal3 s 53706 14560 54506 14680 6 fmc_dmem_request_get[11]
port 225 nsew signal output
rlabel metal3 s 53706 15648 54506 15768 6 fmc_dmem_request_get[12]
port 226 nsew signal output
rlabel metal3 s 53706 16736 54506 16856 6 fmc_dmem_request_get[13]
port 227 nsew signal output
rlabel metal3 s 53706 17824 54506 17944 6 fmc_dmem_request_get[14]
port 228 nsew signal output
rlabel metal3 s 53706 19048 54506 19168 6 fmc_dmem_request_get[15]
port 229 nsew signal output
rlabel metal3 s 53706 20136 54506 20256 6 fmc_dmem_request_get[16]
port 230 nsew signal output
rlabel metal3 s 53706 21224 54506 21344 6 fmc_dmem_request_get[17]
port 231 nsew signal output
rlabel metal3 s 53706 22312 54506 22432 6 fmc_dmem_request_get[18]
port 232 nsew signal output
rlabel metal3 s 53706 23400 54506 23520 6 fmc_dmem_request_get[19]
port 233 nsew signal output
rlabel metal3 s 53706 3408 54506 3528 6 fmc_dmem_request_get[1]
port 234 nsew signal output
rlabel metal3 s 53706 24488 54506 24608 6 fmc_dmem_request_get[20]
port 235 nsew signal output
rlabel metal3 s 53706 25712 54506 25832 6 fmc_dmem_request_get[21]
port 236 nsew signal output
rlabel metal3 s 53706 26800 54506 26920 6 fmc_dmem_request_get[22]
port 237 nsew signal output
rlabel metal3 s 53706 27888 54506 28008 6 fmc_dmem_request_get[23]
port 238 nsew signal output
rlabel metal3 s 53706 28976 54506 29096 6 fmc_dmem_request_get[24]
port 239 nsew signal output
rlabel metal3 s 53706 30064 54506 30184 6 fmc_dmem_request_get[25]
port 240 nsew signal output
rlabel metal3 s 53706 31152 54506 31272 6 fmc_dmem_request_get[26]
port 241 nsew signal output
rlabel metal3 s 53706 32376 54506 32496 6 fmc_dmem_request_get[27]
port 242 nsew signal output
rlabel metal3 s 53706 33464 54506 33584 6 fmc_dmem_request_get[28]
port 243 nsew signal output
rlabel metal3 s 53706 34552 54506 34672 6 fmc_dmem_request_get[29]
port 244 nsew signal output
rlabel metal3 s 53706 4496 54506 4616 6 fmc_dmem_request_get[2]
port 245 nsew signal output
rlabel metal3 s 53706 35640 54506 35760 6 fmc_dmem_request_get[30]
port 246 nsew signal output
rlabel metal3 s 53706 36728 54506 36848 6 fmc_dmem_request_get[31]
port 247 nsew signal output
rlabel metal3 s 53706 37952 54506 38072 6 fmc_dmem_request_get[32]
port 248 nsew signal output
rlabel metal3 s 53706 38224 54506 38344 6 fmc_dmem_request_get[33]
port 249 nsew signal output
rlabel metal3 s 53706 38496 54506 38616 6 fmc_dmem_request_get[34]
port 250 nsew signal output
rlabel metal3 s 53706 38768 54506 38888 6 fmc_dmem_request_get[35]
port 251 nsew signal output
rlabel metal3 s 53706 39040 54506 39160 6 fmc_dmem_request_get[36]
port 252 nsew signal output
rlabel metal3 s 53706 39312 54506 39432 6 fmc_dmem_request_get[37]
port 253 nsew signal output
rlabel metal3 s 53706 39584 54506 39704 6 fmc_dmem_request_get[38]
port 254 nsew signal output
rlabel metal3 s 53706 39856 54506 39976 6 fmc_dmem_request_get[39]
port 255 nsew signal output
rlabel metal3 s 53706 5584 54506 5704 6 fmc_dmem_request_get[3]
port 256 nsew signal output
rlabel metal3 s 53706 40128 54506 40248 6 fmc_dmem_request_get[40]
port 257 nsew signal output
rlabel metal3 s 53706 40400 54506 40520 6 fmc_dmem_request_get[41]
port 258 nsew signal output
rlabel metal3 s 53706 40672 54506 40792 6 fmc_dmem_request_get[42]
port 259 nsew signal output
rlabel metal3 s 53706 40944 54506 41064 6 fmc_dmem_request_get[43]
port 260 nsew signal output
rlabel metal3 s 53706 41216 54506 41336 6 fmc_dmem_request_get[44]
port 261 nsew signal output
rlabel metal3 s 53706 41488 54506 41608 6 fmc_dmem_request_get[45]
port 262 nsew signal output
rlabel metal3 s 53706 41760 54506 41880 6 fmc_dmem_request_get[46]
port 263 nsew signal output
rlabel metal3 s 53706 42032 54506 42152 6 fmc_dmem_request_get[47]
port 264 nsew signal output
rlabel metal3 s 53706 42304 54506 42424 6 fmc_dmem_request_get[48]
port 265 nsew signal output
rlabel metal3 s 53706 42576 54506 42696 6 fmc_dmem_request_get[49]
port 266 nsew signal output
rlabel metal3 s 53706 6808 54506 6928 6 fmc_dmem_request_get[4]
port 267 nsew signal output
rlabel metal3 s 53706 42848 54506 42968 6 fmc_dmem_request_get[50]
port 268 nsew signal output
rlabel metal3 s 53706 43120 54506 43240 6 fmc_dmem_request_get[51]
port 269 nsew signal output
rlabel metal3 s 53706 43392 54506 43512 6 fmc_dmem_request_get[52]
port 270 nsew signal output
rlabel metal3 s 53706 43664 54506 43784 6 fmc_dmem_request_get[53]
port 271 nsew signal output
rlabel metal3 s 53706 43936 54506 44056 6 fmc_dmem_request_get[54]
port 272 nsew signal output
rlabel metal3 s 53706 44344 54506 44464 6 fmc_dmem_request_get[55]
port 273 nsew signal output
rlabel metal3 s 53706 44616 54506 44736 6 fmc_dmem_request_get[56]
port 274 nsew signal output
rlabel metal3 s 53706 44888 54506 45008 6 fmc_dmem_request_get[57]
port 275 nsew signal output
rlabel metal3 s 53706 45160 54506 45280 6 fmc_dmem_request_get[58]
port 276 nsew signal output
rlabel metal3 s 53706 45432 54506 45552 6 fmc_dmem_request_get[59]
port 277 nsew signal output
rlabel metal3 s 53706 7896 54506 8016 6 fmc_dmem_request_get[5]
port 278 nsew signal output
rlabel metal3 s 53706 45704 54506 45824 6 fmc_dmem_request_get[60]
port 279 nsew signal output
rlabel metal3 s 53706 45976 54506 46096 6 fmc_dmem_request_get[61]
port 280 nsew signal output
rlabel metal3 s 53706 46248 54506 46368 6 fmc_dmem_request_get[62]
port 281 nsew signal output
rlabel metal3 s 53706 46520 54506 46640 6 fmc_dmem_request_get[63]
port 282 nsew signal output
rlabel metal3 s 53706 46792 54506 46912 6 fmc_dmem_request_get[64]
port 283 nsew signal output
rlabel metal3 s 53706 47064 54506 47184 6 fmc_dmem_request_get[65]
port 284 nsew signal output
rlabel metal3 s 53706 47336 54506 47456 6 fmc_dmem_request_get[66]
port 285 nsew signal output
rlabel metal3 s 53706 47608 54506 47728 6 fmc_dmem_request_get[67]
port 286 nsew signal output
rlabel metal3 s 53706 47880 54506 48000 6 fmc_dmem_request_get[68]
port 287 nsew signal output
rlabel metal3 s 53706 48152 54506 48272 6 fmc_dmem_request_get[69]
port 288 nsew signal output
rlabel metal3 s 53706 8984 54506 9104 6 fmc_dmem_request_get[6]
port 289 nsew signal output
rlabel metal3 s 53706 48424 54506 48544 6 fmc_dmem_request_get[70]
port 290 nsew signal output
rlabel metal3 s 53706 48696 54506 48816 6 fmc_dmem_request_get[71]
port 291 nsew signal output
rlabel metal3 s 53706 48968 54506 49088 6 fmc_dmem_request_get[72]
port 292 nsew signal output
rlabel metal3 s 53706 49240 54506 49360 6 fmc_dmem_request_get[73]
port 293 nsew signal output
rlabel metal3 s 53706 49512 54506 49632 6 fmc_dmem_request_get[74]
port 294 nsew signal output
rlabel metal3 s 53706 49784 54506 49904 6 fmc_dmem_request_get[75]
port 295 nsew signal output
rlabel metal3 s 53706 50056 54506 50176 6 fmc_dmem_request_get[76]
port 296 nsew signal output
rlabel metal3 s 53706 50328 54506 50448 6 fmc_dmem_request_get[77]
port 297 nsew signal output
rlabel metal3 s 53706 50736 54506 50856 6 fmc_dmem_request_get[78]
port 298 nsew signal output
rlabel metal3 s 53706 51008 54506 51128 6 fmc_dmem_request_get[79]
port 299 nsew signal output
rlabel metal3 s 53706 10072 54506 10192 6 fmc_dmem_request_get[7]
port 300 nsew signal output
rlabel metal3 s 53706 51280 54506 51400 6 fmc_dmem_request_get[80]
port 301 nsew signal output
rlabel metal3 s 53706 51552 54506 51672 6 fmc_dmem_request_get[81]
port 302 nsew signal output
rlabel metal3 s 53706 51824 54506 51944 6 fmc_dmem_request_get[82]
port 303 nsew signal output
rlabel metal3 s 53706 52096 54506 52216 6 fmc_dmem_request_get[83]
port 304 nsew signal output
rlabel metal3 s 53706 52368 54506 52488 6 fmc_dmem_request_get[84]
port 305 nsew signal output
rlabel metal3 s 53706 52640 54506 52760 6 fmc_dmem_request_get[85]
port 306 nsew signal output
rlabel metal3 s 53706 52912 54506 53032 6 fmc_dmem_request_get[86]
port 307 nsew signal output
rlabel metal3 s 53706 53184 54506 53304 6 fmc_dmem_request_get[87]
port 308 nsew signal output
rlabel metal3 s 53706 53456 54506 53576 6 fmc_dmem_request_get[88]
port 309 nsew signal output
rlabel metal3 s 53706 53728 54506 53848 6 fmc_dmem_request_get[89]
port 310 nsew signal output
rlabel metal3 s 53706 11160 54506 11280 6 fmc_dmem_request_get[8]
port 311 nsew signal output
rlabel metal3 s 53706 54000 54506 54120 6 fmc_dmem_request_get[90]
port 312 nsew signal output
rlabel metal3 s 53706 54272 54506 54392 6 fmc_dmem_request_get[91]
port 313 nsew signal output
rlabel metal3 s 53706 54544 54506 54664 6 fmc_dmem_request_get[92]
port 314 nsew signal output
rlabel metal3 s 53706 54816 54506 54936 6 fmc_dmem_request_get[93]
port 315 nsew signal output
rlabel metal3 s 53706 55088 54506 55208 6 fmc_dmem_request_get[94]
port 316 nsew signal output
rlabel metal3 s 53706 55360 54506 55480 6 fmc_dmem_request_get[95]
port 317 nsew signal output
rlabel metal3 s 53706 55632 54506 55752 6 fmc_dmem_request_get[96]
port 318 nsew signal output
rlabel metal3 s 53706 55904 54506 56024 6 fmc_dmem_request_get[97]
port 319 nsew signal output
rlabel metal3 s 53706 56176 54506 56296 6 fmc_dmem_request_get[98]
port 320 nsew signal output
rlabel metal3 s 53706 56448 54506 56568 6 fmc_dmem_request_get[99]
port 321 nsew signal output
rlabel metal3 s 53706 12248 54506 12368 6 fmc_dmem_request_get[9]
port 322 nsew signal output
rlabel metal3 s 53706 2592 54506 2712 6 fmc_dmem_response_put[0]
port 323 nsew signal input
rlabel metal3 s 53706 13744 54506 13864 6 fmc_dmem_response_put[10]
port 324 nsew signal input
rlabel metal3 s 53706 14832 54506 14952 6 fmc_dmem_response_put[11]
port 325 nsew signal input
rlabel metal3 s 53706 15920 54506 16040 6 fmc_dmem_response_put[12]
port 326 nsew signal input
rlabel metal3 s 53706 17008 54506 17128 6 fmc_dmem_response_put[13]
port 327 nsew signal input
rlabel metal3 s 53706 18096 54506 18216 6 fmc_dmem_response_put[14]
port 328 nsew signal input
rlabel metal3 s 53706 19320 54506 19440 6 fmc_dmem_response_put[15]
port 329 nsew signal input
rlabel metal3 s 53706 20408 54506 20528 6 fmc_dmem_response_put[16]
port 330 nsew signal input
rlabel metal3 s 53706 21496 54506 21616 6 fmc_dmem_response_put[17]
port 331 nsew signal input
rlabel metal3 s 53706 22584 54506 22704 6 fmc_dmem_response_put[18]
port 332 nsew signal input
rlabel metal3 s 53706 23672 54506 23792 6 fmc_dmem_response_put[19]
port 333 nsew signal input
rlabel metal3 s 53706 3680 54506 3800 6 fmc_dmem_response_put[1]
port 334 nsew signal input
rlabel metal3 s 53706 24760 54506 24880 6 fmc_dmem_response_put[20]
port 335 nsew signal input
rlabel metal3 s 53706 25984 54506 26104 6 fmc_dmem_response_put[21]
port 336 nsew signal input
rlabel metal3 s 53706 27072 54506 27192 6 fmc_dmem_response_put[22]
port 337 nsew signal input
rlabel metal3 s 53706 28160 54506 28280 6 fmc_dmem_response_put[23]
port 338 nsew signal input
rlabel metal3 s 53706 29248 54506 29368 6 fmc_dmem_response_put[24]
port 339 nsew signal input
rlabel metal3 s 53706 30336 54506 30456 6 fmc_dmem_response_put[25]
port 340 nsew signal input
rlabel metal3 s 53706 31424 54506 31544 6 fmc_dmem_response_put[26]
port 341 nsew signal input
rlabel metal3 s 53706 32648 54506 32768 6 fmc_dmem_response_put[27]
port 342 nsew signal input
rlabel metal3 s 53706 33736 54506 33856 6 fmc_dmem_response_put[28]
port 343 nsew signal input
rlabel metal3 s 53706 34824 54506 34944 6 fmc_dmem_response_put[29]
port 344 nsew signal input
rlabel metal3 s 53706 4768 54506 4888 6 fmc_dmem_response_put[2]
port 345 nsew signal input
rlabel metal3 s 53706 35912 54506 36032 6 fmc_dmem_response_put[30]
port 346 nsew signal input
rlabel metal3 s 53706 37000 54506 37120 6 fmc_dmem_response_put[31]
port 347 nsew signal input
rlabel metal3 s 53706 5856 54506 5976 6 fmc_dmem_response_put[3]
port 348 nsew signal input
rlabel metal3 s 53706 7080 54506 7200 6 fmc_dmem_response_put[4]
port 349 nsew signal input
rlabel metal3 s 53706 8168 54506 8288 6 fmc_dmem_response_put[5]
port 350 nsew signal input
rlabel metal3 s 53706 9256 54506 9376 6 fmc_dmem_response_put[6]
port 351 nsew signal input
rlabel metal3 s 53706 10344 54506 10464 6 fmc_dmem_response_put[7]
port 352 nsew signal input
rlabel metal3 s 53706 11432 54506 11552 6 fmc_dmem_response_put[8]
port 353 nsew signal input
rlabel metal3 s 53706 12520 54506 12640 6 fmc_dmem_response_put[9]
port 354 nsew signal input
rlabel metal3 s 53706 2864 54506 2984 6 fmc_imem_request_get[0]
port 355 nsew signal output
rlabel metal3 s 53706 14016 54506 14136 6 fmc_imem_request_get[10]
port 356 nsew signal output
rlabel metal3 s 53706 15104 54506 15224 6 fmc_imem_request_get[11]
port 357 nsew signal output
rlabel metal3 s 53706 16192 54506 16312 6 fmc_imem_request_get[12]
port 358 nsew signal output
rlabel metal3 s 53706 17280 54506 17400 6 fmc_imem_request_get[13]
port 359 nsew signal output
rlabel metal3 s 53706 18368 54506 18488 6 fmc_imem_request_get[14]
port 360 nsew signal output
rlabel metal3 s 53706 19592 54506 19712 6 fmc_imem_request_get[15]
port 361 nsew signal output
rlabel metal3 s 53706 20680 54506 20800 6 fmc_imem_request_get[16]
port 362 nsew signal output
rlabel metal3 s 53706 21768 54506 21888 6 fmc_imem_request_get[17]
port 363 nsew signal output
rlabel metal3 s 53706 22856 54506 22976 6 fmc_imem_request_get[18]
port 364 nsew signal output
rlabel metal3 s 53706 23944 54506 24064 6 fmc_imem_request_get[19]
port 365 nsew signal output
rlabel metal3 s 53706 3952 54506 4072 6 fmc_imem_request_get[1]
port 366 nsew signal output
rlabel metal3 s 53706 25032 54506 25152 6 fmc_imem_request_get[20]
port 367 nsew signal output
rlabel metal3 s 53706 26256 54506 26376 6 fmc_imem_request_get[21]
port 368 nsew signal output
rlabel metal3 s 53706 27344 54506 27464 6 fmc_imem_request_get[22]
port 369 nsew signal output
rlabel metal3 s 53706 28432 54506 28552 6 fmc_imem_request_get[23]
port 370 nsew signal output
rlabel metal3 s 53706 29520 54506 29640 6 fmc_imem_request_get[24]
port 371 nsew signal output
rlabel metal3 s 53706 30608 54506 30728 6 fmc_imem_request_get[25]
port 372 nsew signal output
rlabel metal3 s 53706 31832 54506 31952 6 fmc_imem_request_get[26]
port 373 nsew signal output
rlabel metal3 s 53706 32920 54506 33040 6 fmc_imem_request_get[27]
port 374 nsew signal output
rlabel metal3 s 53706 34008 54506 34128 6 fmc_imem_request_get[28]
port 375 nsew signal output
rlabel metal3 s 53706 35096 54506 35216 6 fmc_imem_request_get[29]
port 376 nsew signal output
rlabel metal3 s 53706 5040 54506 5160 6 fmc_imem_request_get[2]
port 377 nsew signal output
rlabel metal3 s 53706 36184 54506 36304 6 fmc_imem_request_get[30]
port 378 nsew signal output
rlabel metal3 s 53706 37272 54506 37392 6 fmc_imem_request_get[31]
port 379 nsew signal output
rlabel metal3 s 53706 6128 54506 6248 6 fmc_imem_request_get[3]
port 380 nsew signal output
rlabel metal3 s 53706 7352 54506 7472 6 fmc_imem_request_get[4]
port 381 nsew signal output
rlabel metal3 s 53706 8440 54506 8560 6 fmc_imem_request_get[5]
port 382 nsew signal output
rlabel metal3 s 53706 9528 54506 9648 6 fmc_imem_request_get[6]
port 383 nsew signal output
rlabel metal3 s 53706 10616 54506 10736 6 fmc_imem_request_get[7]
port 384 nsew signal output
rlabel metal3 s 53706 11704 54506 11824 6 fmc_imem_request_get[8]
port 385 nsew signal output
rlabel metal3 s 53706 12928 54506 13048 6 fmc_imem_request_get[9]
port 386 nsew signal output
rlabel metal3 s 53706 3136 54506 3256 6 fmc_imem_response_put[0]
port 387 nsew signal input
rlabel metal3 s 53706 14288 54506 14408 6 fmc_imem_response_put[10]
port 388 nsew signal input
rlabel metal3 s 53706 15376 54506 15496 6 fmc_imem_response_put[11]
port 389 nsew signal input
rlabel metal3 s 53706 16464 54506 16584 6 fmc_imem_response_put[12]
port 390 nsew signal input
rlabel metal3 s 53706 17552 54506 17672 6 fmc_imem_response_put[13]
port 391 nsew signal input
rlabel metal3 s 53706 18640 54506 18760 6 fmc_imem_response_put[14]
port 392 nsew signal input
rlabel metal3 s 53706 19864 54506 19984 6 fmc_imem_response_put[15]
port 393 nsew signal input
rlabel metal3 s 53706 20952 54506 21072 6 fmc_imem_response_put[16]
port 394 nsew signal input
rlabel metal3 s 53706 22040 54506 22160 6 fmc_imem_response_put[17]
port 395 nsew signal input
rlabel metal3 s 53706 23128 54506 23248 6 fmc_imem_response_put[18]
port 396 nsew signal input
rlabel metal3 s 53706 24216 54506 24336 6 fmc_imem_response_put[19]
port 397 nsew signal input
rlabel metal3 s 53706 4224 54506 4344 6 fmc_imem_response_put[1]
port 398 nsew signal input
rlabel metal3 s 53706 25440 54506 25560 6 fmc_imem_response_put[20]
port 399 nsew signal input
rlabel metal3 s 53706 26528 54506 26648 6 fmc_imem_response_put[21]
port 400 nsew signal input
rlabel metal3 s 53706 27616 54506 27736 6 fmc_imem_response_put[22]
port 401 nsew signal input
rlabel metal3 s 53706 28704 54506 28824 6 fmc_imem_response_put[23]
port 402 nsew signal input
rlabel metal3 s 53706 29792 54506 29912 6 fmc_imem_response_put[24]
port 403 nsew signal input
rlabel metal3 s 53706 30880 54506 31000 6 fmc_imem_response_put[25]
port 404 nsew signal input
rlabel metal3 s 53706 32104 54506 32224 6 fmc_imem_response_put[26]
port 405 nsew signal input
rlabel metal3 s 53706 33192 54506 33312 6 fmc_imem_response_put[27]
port 406 nsew signal input
rlabel metal3 s 53706 34280 54506 34400 6 fmc_imem_response_put[28]
port 407 nsew signal input
rlabel metal3 s 53706 35368 54506 35488 6 fmc_imem_response_put[29]
port 408 nsew signal input
rlabel metal3 s 53706 5312 54506 5432 6 fmc_imem_response_put[2]
port 409 nsew signal input
rlabel metal3 s 53706 36456 54506 36576 6 fmc_imem_response_put[30]
port 410 nsew signal input
rlabel metal3 s 53706 37544 54506 37664 6 fmc_imem_response_put[31]
port 411 nsew signal input
rlabel metal3 s 53706 6536 54506 6656 6 fmc_imem_response_put[3]
port 412 nsew signal input
rlabel metal3 s 53706 7624 54506 7744 6 fmc_imem_response_put[4]
port 413 nsew signal input
rlabel metal3 s 53706 8712 54506 8832 6 fmc_imem_response_put[5]
port 414 nsew signal input
rlabel metal3 s 53706 9800 54506 9920 6 fmc_imem_response_put[6]
port 415 nsew signal input
rlabel metal3 s 53706 10888 54506 11008 6 fmc_imem_response_put[7]
port 416 nsew signal input
rlabel metal3 s 53706 11976 54506 12096 6 fmc_imem_response_put[8]
port 417 nsew signal input
rlabel metal3 s 53706 13200 54506 13320 6 fmc_imem_response_put[9]
port 418 nsew signal input
rlabel metal2 s 2226 55850 2282 56650 6 ram_dmem_request_get[0]
port 419 nsew signal output
rlabel metal2 s 12898 55850 12954 56650 6 ram_dmem_request_get[10]
port 420 nsew signal output
rlabel metal2 s 13910 55850 13966 56650 6 ram_dmem_request_get[11]
port 421 nsew signal output
rlabel metal2 s 15014 55850 15070 56650 6 ram_dmem_request_get[12]
port 422 nsew signal output
rlabel metal2 s 16118 55850 16174 56650 6 ram_dmem_request_get[13]
port 423 nsew signal output
rlabel metal2 s 17130 55850 17186 56650 6 ram_dmem_request_get[14]
port 424 nsew signal output
rlabel metal2 s 18234 55850 18290 56650 6 ram_dmem_request_get[15]
port 425 nsew signal output
rlabel metal2 s 19246 55850 19302 56650 6 ram_dmem_request_get[16]
port 426 nsew signal output
rlabel metal2 s 20350 55850 20406 56650 6 ram_dmem_request_get[17]
port 427 nsew signal output
rlabel metal2 s 21454 55850 21510 56650 6 ram_dmem_request_get[18]
port 428 nsew signal output
rlabel metal2 s 22466 55850 22522 56650 6 ram_dmem_request_get[19]
port 429 nsew signal output
rlabel metal2 s 3238 55850 3294 56650 6 ram_dmem_request_get[1]
port 430 nsew signal output
rlabel metal2 s 23570 55850 23626 56650 6 ram_dmem_request_get[20]
port 431 nsew signal output
rlabel metal2 s 24582 55850 24638 56650 6 ram_dmem_request_get[21]
port 432 nsew signal output
rlabel metal2 s 25686 55850 25742 56650 6 ram_dmem_request_get[22]
port 433 nsew signal output
rlabel metal2 s 26790 55850 26846 56650 6 ram_dmem_request_get[23]
port 434 nsew signal output
rlabel metal2 s 27802 55850 27858 56650 6 ram_dmem_request_get[24]
port 435 nsew signal output
rlabel metal2 s 28906 55850 28962 56650 6 ram_dmem_request_get[25]
port 436 nsew signal output
rlabel metal2 s 30010 55850 30066 56650 6 ram_dmem_request_get[26]
port 437 nsew signal output
rlabel metal2 s 31022 55850 31078 56650 6 ram_dmem_request_get[27]
port 438 nsew signal output
rlabel metal2 s 32126 55850 32182 56650 6 ram_dmem_request_get[28]
port 439 nsew signal output
rlabel metal2 s 33138 55850 33194 56650 6 ram_dmem_request_get[29]
port 440 nsew signal output
rlabel metal2 s 4342 55850 4398 56650 6 ram_dmem_request_get[2]
port 441 nsew signal output
rlabel metal2 s 34242 55850 34298 56650 6 ram_dmem_request_get[30]
port 442 nsew signal output
rlabel metal2 s 35346 55850 35402 56650 6 ram_dmem_request_get[31]
port 443 nsew signal output
rlabel metal2 s 36358 55850 36414 56650 6 ram_dmem_request_get[32]
port 444 nsew signal output
rlabel metal2 s 36634 55850 36690 56650 6 ram_dmem_request_get[33]
port 445 nsew signal output
rlabel metal2 s 36910 55850 36966 56650 6 ram_dmem_request_get[34]
port 446 nsew signal output
rlabel metal2 s 37186 55850 37242 56650 6 ram_dmem_request_get[35]
port 447 nsew signal output
rlabel metal2 s 37462 55850 37518 56650 6 ram_dmem_request_get[36]
port 448 nsew signal output
rlabel metal2 s 37738 55850 37794 56650 6 ram_dmem_request_get[37]
port 449 nsew signal output
rlabel metal2 s 38014 55850 38070 56650 6 ram_dmem_request_get[38]
port 450 nsew signal output
rlabel metal2 s 38198 55850 38254 56650 6 ram_dmem_request_get[39]
port 451 nsew signal output
rlabel metal2 s 5446 55850 5502 56650 6 ram_dmem_request_get[3]
port 452 nsew signal output
rlabel metal2 s 38474 55850 38530 56650 6 ram_dmem_request_get[40]
port 453 nsew signal output
rlabel metal2 s 38750 55850 38806 56650 6 ram_dmem_request_get[41]
port 454 nsew signal output
rlabel metal2 s 39026 55850 39082 56650 6 ram_dmem_request_get[42]
port 455 nsew signal output
rlabel metal2 s 39302 55850 39358 56650 6 ram_dmem_request_get[43]
port 456 nsew signal output
rlabel metal2 s 39578 55850 39634 56650 6 ram_dmem_request_get[44]
port 457 nsew signal output
rlabel metal2 s 39854 55850 39910 56650 6 ram_dmem_request_get[45]
port 458 nsew signal output
rlabel metal2 s 40130 55850 40186 56650 6 ram_dmem_request_get[46]
port 459 nsew signal output
rlabel metal2 s 40406 55850 40462 56650 6 ram_dmem_request_get[47]
port 460 nsew signal output
rlabel metal2 s 40682 55850 40738 56650 6 ram_dmem_request_get[48]
port 461 nsew signal output
rlabel metal2 s 40958 55850 41014 56650 6 ram_dmem_request_get[49]
port 462 nsew signal output
rlabel metal2 s 6458 55850 6514 56650 6 ram_dmem_request_get[4]
port 463 nsew signal output
rlabel metal2 s 41142 55850 41198 56650 6 ram_dmem_request_get[50]
port 464 nsew signal output
rlabel metal2 s 41418 55850 41474 56650 6 ram_dmem_request_get[51]
port 465 nsew signal output
rlabel metal2 s 41694 55850 41750 56650 6 ram_dmem_request_get[52]
port 466 nsew signal output
rlabel metal2 s 41970 55850 42026 56650 6 ram_dmem_request_get[53]
port 467 nsew signal output
rlabel metal2 s 42246 55850 42302 56650 6 ram_dmem_request_get[54]
port 468 nsew signal output
rlabel metal2 s 42522 55850 42578 56650 6 ram_dmem_request_get[55]
port 469 nsew signal output
rlabel metal2 s 42798 55850 42854 56650 6 ram_dmem_request_get[56]
port 470 nsew signal output
rlabel metal2 s 43074 55850 43130 56650 6 ram_dmem_request_get[57]
port 471 nsew signal output
rlabel metal2 s 43350 55850 43406 56650 6 ram_dmem_request_get[58]
port 472 nsew signal output
rlabel metal2 s 43626 55850 43682 56650 6 ram_dmem_request_get[59]
port 473 nsew signal output
rlabel metal2 s 7562 55850 7618 56650 6 ram_dmem_request_get[5]
port 474 nsew signal output
rlabel metal2 s 43810 55850 43866 56650 6 ram_dmem_request_get[60]
port 475 nsew signal output
rlabel metal2 s 44086 55850 44142 56650 6 ram_dmem_request_get[61]
port 476 nsew signal output
rlabel metal2 s 44362 55850 44418 56650 6 ram_dmem_request_get[62]
port 477 nsew signal output
rlabel metal2 s 44638 55850 44694 56650 6 ram_dmem_request_get[63]
port 478 nsew signal output
rlabel metal2 s 44914 55850 44970 56650 6 ram_dmem_request_get[64]
port 479 nsew signal output
rlabel metal2 s 45190 55850 45246 56650 6 ram_dmem_request_get[65]
port 480 nsew signal output
rlabel metal2 s 45466 55850 45522 56650 6 ram_dmem_request_get[66]
port 481 nsew signal output
rlabel metal2 s 45742 55850 45798 56650 6 ram_dmem_request_get[67]
port 482 nsew signal output
rlabel metal2 s 46018 55850 46074 56650 6 ram_dmem_request_get[68]
port 483 nsew signal output
rlabel metal2 s 46294 55850 46350 56650 6 ram_dmem_request_get[69]
port 484 nsew signal output
rlabel metal2 s 8574 55850 8630 56650 6 ram_dmem_request_get[6]
port 485 nsew signal output
rlabel metal2 s 46478 55850 46534 56650 6 ram_dmem_request_get[70]
port 486 nsew signal output
rlabel metal2 s 46754 55850 46810 56650 6 ram_dmem_request_get[71]
port 487 nsew signal output
rlabel metal2 s 47030 55850 47086 56650 6 ram_dmem_request_get[72]
port 488 nsew signal output
rlabel metal2 s 47306 55850 47362 56650 6 ram_dmem_request_get[73]
port 489 nsew signal output
rlabel metal2 s 47582 55850 47638 56650 6 ram_dmem_request_get[74]
port 490 nsew signal output
rlabel metal2 s 47858 55850 47914 56650 6 ram_dmem_request_get[75]
port 491 nsew signal output
rlabel metal2 s 48134 55850 48190 56650 6 ram_dmem_request_get[76]
port 492 nsew signal output
rlabel metal2 s 48410 55850 48466 56650 6 ram_dmem_request_get[77]
port 493 nsew signal output
rlabel metal2 s 48686 55850 48742 56650 6 ram_dmem_request_get[78]
port 494 nsew signal output
rlabel metal2 s 48962 55850 49018 56650 6 ram_dmem_request_get[79]
port 495 nsew signal output
rlabel metal2 s 9678 55850 9734 56650 6 ram_dmem_request_get[7]
port 496 nsew signal output
rlabel metal2 s 49146 55850 49202 56650 6 ram_dmem_request_get[80]
port 497 nsew signal output
rlabel metal2 s 49422 55850 49478 56650 6 ram_dmem_request_get[81]
port 498 nsew signal output
rlabel metal2 s 49698 55850 49754 56650 6 ram_dmem_request_get[82]
port 499 nsew signal output
rlabel metal2 s 49974 55850 50030 56650 6 ram_dmem_request_get[83]
port 500 nsew signal output
rlabel metal2 s 50250 55850 50306 56650 6 ram_dmem_request_get[84]
port 501 nsew signal output
rlabel metal2 s 50526 55850 50582 56650 6 ram_dmem_request_get[85]
port 502 nsew signal output
rlabel metal2 s 50802 55850 50858 56650 6 ram_dmem_request_get[86]
port 503 nsew signal output
rlabel metal2 s 51078 55850 51134 56650 6 ram_dmem_request_get[87]
port 504 nsew signal output
rlabel metal2 s 51354 55850 51410 56650 6 ram_dmem_request_get[88]
port 505 nsew signal output
rlabel metal2 s 51630 55850 51686 56650 6 ram_dmem_request_get[89]
port 506 nsew signal output
rlabel metal2 s 10782 55850 10838 56650 6 ram_dmem_request_get[8]
port 507 nsew signal output
rlabel metal2 s 51814 55850 51870 56650 6 ram_dmem_request_get[90]
port 508 nsew signal output
rlabel metal2 s 52090 55850 52146 56650 6 ram_dmem_request_get[91]
port 509 nsew signal output
rlabel metal2 s 52366 55850 52422 56650 6 ram_dmem_request_get[92]
port 510 nsew signal output
rlabel metal2 s 52642 55850 52698 56650 6 ram_dmem_request_get[93]
port 511 nsew signal output
rlabel metal2 s 52918 55850 52974 56650 6 ram_dmem_request_get[94]
port 512 nsew signal output
rlabel metal2 s 53194 55850 53250 56650 6 ram_dmem_request_get[95]
port 513 nsew signal output
rlabel metal2 s 53470 55850 53526 56650 6 ram_dmem_request_get[96]
port 514 nsew signal output
rlabel metal2 s 53746 55850 53802 56650 6 ram_dmem_request_get[97]
port 515 nsew signal output
rlabel metal2 s 54022 55850 54078 56650 6 ram_dmem_request_get[98]
port 516 nsew signal output
rlabel metal2 s 54298 55850 54354 56650 6 ram_dmem_request_get[99]
port 517 nsew signal output
rlabel metal2 s 11794 55850 11850 56650 6 ram_dmem_request_get[9]
port 518 nsew signal output
rlabel metal2 s 2502 55850 2558 56650 6 ram_dmem_response_put[0]
port 519 nsew signal input
rlabel metal2 s 13174 55850 13230 56650 6 ram_dmem_response_put[10]
port 520 nsew signal input
rlabel metal2 s 14186 55850 14242 56650 6 ram_dmem_response_put[11]
port 521 nsew signal input
rlabel metal2 s 15290 55850 15346 56650 6 ram_dmem_response_put[12]
port 522 nsew signal input
rlabel metal2 s 16394 55850 16450 56650 6 ram_dmem_response_put[13]
port 523 nsew signal input
rlabel metal2 s 17406 55850 17462 56650 6 ram_dmem_response_put[14]
port 524 nsew signal input
rlabel metal2 s 18510 55850 18566 56650 6 ram_dmem_response_put[15]
port 525 nsew signal input
rlabel metal2 s 19522 55850 19578 56650 6 ram_dmem_response_put[16]
port 526 nsew signal input
rlabel metal2 s 20626 55850 20682 56650 6 ram_dmem_response_put[17]
port 527 nsew signal input
rlabel metal2 s 21730 55850 21786 56650 6 ram_dmem_response_put[18]
port 528 nsew signal input
rlabel metal2 s 22742 55850 22798 56650 6 ram_dmem_response_put[19]
port 529 nsew signal input
rlabel metal2 s 3514 55850 3570 56650 6 ram_dmem_response_put[1]
port 530 nsew signal input
rlabel metal2 s 23846 55850 23902 56650 6 ram_dmem_response_put[20]
port 531 nsew signal input
rlabel metal2 s 24858 55850 24914 56650 6 ram_dmem_response_put[21]
port 532 nsew signal input
rlabel metal2 s 25962 55850 26018 56650 6 ram_dmem_response_put[22]
port 533 nsew signal input
rlabel metal2 s 27066 55850 27122 56650 6 ram_dmem_response_put[23]
port 534 nsew signal input
rlabel metal2 s 28078 55850 28134 56650 6 ram_dmem_response_put[24]
port 535 nsew signal input
rlabel metal2 s 29182 55850 29238 56650 6 ram_dmem_response_put[25]
port 536 nsew signal input
rlabel metal2 s 30194 55850 30250 56650 6 ram_dmem_response_put[26]
port 537 nsew signal input
rlabel metal2 s 31298 55850 31354 56650 6 ram_dmem_response_put[27]
port 538 nsew signal input
rlabel metal2 s 32402 55850 32458 56650 6 ram_dmem_response_put[28]
port 539 nsew signal input
rlabel metal2 s 33414 55850 33470 56650 6 ram_dmem_response_put[29]
port 540 nsew signal input
rlabel metal2 s 4618 55850 4674 56650 6 ram_dmem_response_put[2]
port 541 nsew signal input
rlabel metal2 s 34518 55850 34574 56650 6 ram_dmem_response_put[30]
port 542 nsew signal input
rlabel metal2 s 35530 55850 35586 56650 6 ram_dmem_response_put[31]
port 543 nsew signal input
rlabel metal2 s 5630 55850 5686 56650 6 ram_dmem_response_put[3]
port 544 nsew signal input
rlabel metal2 s 6734 55850 6790 56650 6 ram_dmem_response_put[4]
port 545 nsew signal input
rlabel metal2 s 7838 55850 7894 56650 6 ram_dmem_response_put[5]
port 546 nsew signal input
rlabel metal2 s 8850 55850 8906 56650 6 ram_dmem_response_put[6]
port 547 nsew signal input
rlabel metal2 s 9954 55850 10010 56650 6 ram_dmem_response_put[7]
port 548 nsew signal input
rlabel metal2 s 10966 55850 11022 56650 6 ram_dmem_response_put[8]
port 549 nsew signal input
rlabel metal2 s 12070 55850 12126 56650 6 ram_dmem_response_put[9]
port 550 nsew signal input
rlabel metal2 s 2778 55850 2834 56650 6 ram_imem_request_get[0]
port 551 nsew signal output
rlabel metal2 s 13450 55850 13506 56650 6 ram_imem_request_get[10]
port 552 nsew signal output
rlabel metal2 s 14462 55850 14518 56650 6 ram_imem_request_get[11]
port 553 nsew signal output
rlabel metal2 s 15566 55850 15622 56650 6 ram_imem_request_get[12]
port 554 nsew signal output
rlabel metal2 s 16578 55850 16634 56650 6 ram_imem_request_get[13]
port 555 nsew signal output
rlabel metal2 s 17682 55850 17738 56650 6 ram_imem_request_get[14]
port 556 nsew signal output
rlabel metal2 s 18786 55850 18842 56650 6 ram_imem_request_get[15]
port 557 nsew signal output
rlabel metal2 s 19798 55850 19854 56650 6 ram_imem_request_get[16]
port 558 nsew signal output
rlabel metal2 s 20902 55850 20958 56650 6 ram_imem_request_get[17]
port 559 nsew signal output
rlabel metal2 s 21914 55850 21970 56650 6 ram_imem_request_get[18]
port 560 nsew signal output
rlabel metal2 s 23018 55850 23074 56650 6 ram_imem_request_get[19]
port 561 nsew signal output
rlabel metal2 s 3790 55850 3846 56650 6 ram_imem_request_get[1]
port 562 nsew signal output
rlabel metal2 s 24122 55850 24178 56650 6 ram_imem_request_get[20]
port 563 nsew signal output
rlabel metal2 s 25134 55850 25190 56650 6 ram_imem_request_get[21]
port 564 nsew signal output
rlabel metal2 s 26238 55850 26294 56650 6 ram_imem_request_get[22]
port 565 nsew signal output
rlabel metal2 s 27342 55850 27398 56650 6 ram_imem_request_get[23]
port 566 nsew signal output
rlabel metal2 s 28354 55850 28410 56650 6 ram_imem_request_get[24]
port 567 nsew signal output
rlabel metal2 s 29458 55850 29514 56650 6 ram_imem_request_get[25]
port 568 nsew signal output
rlabel metal2 s 30470 55850 30526 56650 6 ram_imem_request_get[26]
port 569 nsew signal output
rlabel metal2 s 31574 55850 31630 56650 6 ram_imem_request_get[27]
port 570 nsew signal output
rlabel metal2 s 32678 55850 32734 56650 6 ram_imem_request_get[28]
port 571 nsew signal output
rlabel metal2 s 33690 55850 33746 56650 6 ram_imem_request_get[29]
port 572 nsew signal output
rlabel metal2 s 4894 55850 4950 56650 6 ram_imem_request_get[2]
port 573 nsew signal output
rlabel metal2 s 34794 55850 34850 56650 6 ram_imem_request_get[30]
port 574 nsew signal output
rlabel metal2 s 35806 55850 35862 56650 6 ram_imem_request_get[31]
port 575 nsew signal output
rlabel metal2 s 5906 55850 5962 56650 6 ram_imem_request_get[3]
port 576 nsew signal output
rlabel metal2 s 7010 55850 7066 56650 6 ram_imem_request_get[4]
port 577 nsew signal output
rlabel metal2 s 8114 55850 8170 56650 6 ram_imem_request_get[5]
port 578 nsew signal output
rlabel metal2 s 9126 55850 9182 56650 6 ram_imem_request_get[6]
port 579 nsew signal output
rlabel metal2 s 10230 55850 10286 56650 6 ram_imem_request_get[7]
port 580 nsew signal output
rlabel metal2 s 11242 55850 11298 56650 6 ram_imem_request_get[8]
port 581 nsew signal output
rlabel metal2 s 12346 55850 12402 56650 6 ram_imem_request_get[9]
port 582 nsew signal output
rlabel metal2 s 2962 55850 3018 56650 6 ram_imem_response_put[0]
port 583 nsew signal input
rlabel metal2 s 13726 55850 13782 56650 6 ram_imem_response_put[10]
port 584 nsew signal input
rlabel metal2 s 14738 55850 14794 56650 6 ram_imem_response_put[11]
port 585 nsew signal input
rlabel metal2 s 15842 55850 15898 56650 6 ram_imem_response_put[12]
port 586 nsew signal input
rlabel metal2 s 16854 55850 16910 56650 6 ram_imem_response_put[13]
port 587 nsew signal input
rlabel metal2 s 17958 55850 18014 56650 6 ram_imem_response_put[14]
port 588 nsew signal input
rlabel metal2 s 19062 55850 19118 56650 6 ram_imem_response_put[15]
port 589 nsew signal input
rlabel metal2 s 20074 55850 20130 56650 6 ram_imem_response_put[16]
port 590 nsew signal input
rlabel metal2 s 21178 55850 21234 56650 6 ram_imem_response_put[17]
port 591 nsew signal input
rlabel metal2 s 22190 55850 22246 56650 6 ram_imem_response_put[18]
port 592 nsew signal input
rlabel metal2 s 23294 55850 23350 56650 6 ram_imem_response_put[19]
port 593 nsew signal input
rlabel metal2 s 4066 55850 4122 56650 6 ram_imem_response_put[1]
port 594 nsew signal input
rlabel metal2 s 24398 55850 24454 56650 6 ram_imem_response_put[20]
port 595 nsew signal input
rlabel metal2 s 25410 55850 25466 56650 6 ram_imem_response_put[21]
port 596 nsew signal input
rlabel metal2 s 26514 55850 26570 56650 6 ram_imem_response_put[22]
port 597 nsew signal input
rlabel metal2 s 27526 55850 27582 56650 6 ram_imem_response_put[23]
port 598 nsew signal input
rlabel metal2 s 28630 55850 28686 56650 6 ram_imem_response_put[24]
port 599 nsew signal input
rlabel metal2 s 29734 55850 29790 56650 6 ram_imem_response_put[25]
port 600 nsew signal input
rlabel metal2 s 30746 55850 30802 56650 6 ram_imem_response_put[26]
port 601 nsew signal input
rlabel metal2 s 31850 55850 31906 56650 6 ram_imem_response_put[27]
port 602 nsew signal input
rlabel metal2 s 32862 55850 32918 56650 6 ram_imem_response_put[28]
port 603 nsew signal input
rlabel metal2 s 33966 55850 34022 56650 6 ram_imem_response_put[29]
port 604 nsew signal input
rlabel metal2 s 5170 55850 5226 56650 6 ram_imem_response_put[2]
port 605 nsew signal input
rlabel metal2 s 35070 55850 35126 56650 6 ram_imem_response_put[30]
port 606 nsew signal input
rlabel metal2 s 36082 55850 36138 56650 6 ram_imem_response_put[31]
port 607 nsew signal input
rlabel metal2 s 6182 55850 6238 56650 6 ram_imem_response_put[3]
port 608 nsew signal input
rlabel metal2 s 7286 55850 7342 56650 6 ram_imem_response_put[4]
port 609 nsew signal input
rlabel metal2 s 8298 55850 8354 56650 6 ram_imem_response_put[5]
port 610 nsew signal input
rlabel metal2 s 9402 55850 9458 56650 6 ram_imem_response_put[6]
port 611 nsew signal input
rlabel metal2 s 10506 55850 10562 56650 6 ram_imem_response_put[7]
port 612 nsew signal input
rlabel metal2 s 11518 55850 11574 56650 6 ram_imem_response_put[8]
port 613 nsew signal input
rlabel metal2 s 12622 55850 12678 56650 6 ram_imem_response_put[9]
port 614 nsew signal input
rlabel metal4 s 4208 2128 4528 54448 6 vccd1
port 615 nsew power input
rlabel metal4 s 34928 2128 35248 54448 6 vccd1
port 615 nsew power input
rlabel metal4 s 19568 2128 19888 54448 6 vssd1
port 616 nsew ground input
rlabel metal4 s 50288 2128 50608 54448 6 vssd1
port 616 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 54506 56650
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9336382
string GDS_FILE /home/q3k/sky130/qf105/openlane/mkLanaiFrontend/runs/mkLanaiFrontend/results/finishing/mkLanaiFrontend.magic.gds
string GDS_START 448676
<< end >>

