* NGSPICE file created from mkQF100Memory.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__fakediode_2 abstract view
.subckt sky130_ef_sc_hd__fakediode_2 DIODE VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_2 abstract view
.subckt sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_1 abstract view
.subckt sky130_fd_sc_hd__o311ai_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_1 abstract view
.subckt sky130_fd_sc_hd__o41ai_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

.subckt mkQF100Memory CLK EN_memory_dmem_request_put EN_memory_dmem_response_get EN_memory_imem_request_put
+ EN_memory_imem_response_get RDY_memory_dmem_request_put RDY_memory_dmem_response_get
+ RDY_memory_imem_request_put RDY_memory_imem_response_get RST_N VGND VPWR memory_dmem_request_put[0]
+ memory_dmem_request_put[10] memory_dmem_request_put[11] memory_dmem_request_put[12]
+ memory_dmem_request_put[13] memory_dmem_request_put[14] memory_dmem_request_put[15]
+ memory_dmem_request_put[16] memory_dmem_request_put[17] memory_dmem_request_put[18]
+ memory_dmem_request_put[19] memory_dmem_request_put[1] memory_dmem_request_put[20]
+ memory_dmem_request_put[21] memory_dmem_request_put[22] memory_dmem_request_put[23]
+ memory_dmem_request_put[24] memory_dmem_request_put[25] memory_dmem_request_put[26]
+ memory_dmem_request_put[27] memory_dmem_request_put[28] memory_dmem_request_put[29]
+ memory_dmem_request_put[2] memory_dmem_request_put[30] memory_dmem_request_put[31]
+ memory_dmem_request_put[32] memory_dmem_request_put[33] memory_dmem_request_put[34]
+ memory_dmem_request_put[35] memory_dmem_request_put[36] memory_dmem_request_put[37]
+ memory_dmem_request_put[38] memory_dmem_request_put[39] memory_dmem_request_put[3]
+ memory_dmem_request_put[40] memory_dmem_request_put[41] memory_dmem_request_put[42]
+ memory_dmem_request_put[43] memory_dmem_request_put[44] memory_dmem_request_put[45]
+ memory_dmem_request_put[46] memory_dmem_request_put[47] memory_dmem_request_put[48]
+ memory_dmem_request_put[49] memory_dmem_request_put[4] memory_dmem_request_put[50]
+ memory_dmem_request_put[51] memory_dmem_request_put[52] memory_dmem_request_put[53]
+ memory_dmem_request_put[54] memory_dmem_request_put[55] memory_dmem_request_put[56]
+ memory_dmem_request_put[57] memory_dmem_request_put[58] memory_dmem_request_put[59]
+ memory_dmem_request_put[5] memory_dmem_request_put[60] memory_dmem_request_put[61]
+ memory_dmem_request_put[62] memory_dmem_request_put[63] memory_dmem_request_put[64]
+ memory_dmem_request_put[65] memory_dmem_request_put[66] memory_dmem_request_put[67]
+ memory_dmem_request_put[68] memory_dmem_request_put[69] memory_dmem_request_put[6]
+ memory_dmem_request_put[70] memory_dmem_request_put[71] memory_dmem_request_put[72]
+ memory_dmem_request_put[73] memory_dmem_request_put[74] memory_dmem_request_put[75]
+ memory_dmem_request_put[76] memory_dmem_request_put[77] memory_dmem_request_put[78]
+ memory_dmem_request_put[79] memory_dmem_request_put[7] memory_dmem_request_put[80]
+ memory_dmem_request_put[81] memory_dmem_request_put[82] memory_dmem_request_put[83]
+ memory_dmem_request_put[84] memory_dmem_request_put[85] memory_dmem_request_put[86]
+ memory_dmem_request_put[87] memory_dmem_request_put[88] memory_dmem_request_put[89]
+ memory_dmem_request_put[8] memory_dmem_request_put[90] memory_dmem_request_put[91]
+ memory_dmem_request_put[92] memory_dmem_request_put[93] memory_dmem_request_put[94]
+ memory_dmem_request_put[95] memory_dmem_request_put[96] memory_dmem_request_put[97]
+ memory_dmem_request_put[98] memory_dmem_request_put[99] memory_dmem_request_put[9]
+ memory_dmem_response_get[0] memory_dmem_response_get[10] memory_dmem_response_get[11]
+ memory_dmem_response_get[12] memory_dmem_response_get[13] memory_dmem_response_get[14]
+ memory_dmem_response_get[15] memory_dmem_response_get[16] memory_dmem_response_get[17]
+ memory_dmem_response_get[18] memory_dmem_response_get[19] memory_dmem_response_get[1]
+ memory_dmem_response_get[20] memory_dmem_response_get[21] memory_dmem_response_get[22]
+ memory_dmem_response_get[23] memory_dmem_response_get[24] memory_dmem_response_get[25]
+ memory_dmem_response_get[26] memory_dmem_response_get[27] memory_dmem_response_get[28]
+ memory_dmem_response_get[29] memory_dmem_response_get[2] memory_dmem_response_get[30]
+ memory_dmem_response_get[31] memory_dmem_response_get[3] memory_dmem_response_get[4]
+ memory_dmem_response_get[5] memory_dmem_response_get[6] memory_dmem_response_get[7]
+ memory_dmem_response_get[8] memory_dmem_response_get[9] memory_imem_request_put[0]
+ memory_imem_request_put[10] memory_imem_request_put[11] memory_imem_request_put[12]
+ memory_imem_request_put[13] memory_imem_request_put[14] memory_imem_request_put[15]
+ memory_imem_request_put[16] memory_imem_request_put[17] memory_imem_request_put[18]
+ memory_imem_request_put[19] memory_imem_request_put[1] memory_imem_request_put[20]
+ memory_imem_request_put[21] memory_imem_request_put[22] memory_imem_request_put[23]
+ memory_imem_request_put[24] memory_imem_request_put[25] memory_imem_request_put[26]
+ memory_imem_request_put[27] memory_imem_request_put[28] memory_imem_request_put[29]
+ memory_imem_request_put[2] memory_imem_request_put[30] memory_imem_request_put[31]
+ memory_imem_request_put[3] memory_imem_request_put[4] memory_imem_request_put[5]
+ memory_imem_request_put[6] memory_imem_request_put[7] memory_imem_request_put[8]
+ memory_imem_request_put[9] memory_imem_response_get[0] memory_imem_response_get[10]
+ memory_imem_response_get[11] memory_imem_response_get[12] memory_imem_response_get[13]
+ memory_imem_response_get[14] memory_imem_response_get[15] memory_imem_response_get[16]
+ memory_imem_response_get[17] memory_imem_response_get[18] memory_imem_response_get[19]
+ memory_imem_response_get[1] memory_imem_response_get[20] memory_imem_response_get[21]
+ memory_imem_response_get[22] memory_imem_response_get[23] memory_imem_response_get[24]
+ memory_imem_response_get[25] memory_imem_response_get[26] memory_imem_response_get[27]
+ memory_imem_response_get[28] memory_imem_response_get[29] memory_imem_response_get[2]
+ memory_imem_response_get[30] memory_imem_response_get[31] memory_imem_response_get[3]
+ memory_imem_response_get[4] memory_imem_response_get[5] memory_imem_response_get[6]
+ memory_imem_response_get[7] memory_imem_response_get[8] memory_imem_response_get[9]
XANTENNA__4935__A _5118_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3155_ _3162_/A VGND VGND VPWR VPWR _3603_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__3691__A2 _3690_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3086_ _6185_/Q _6077_/Q _3094_/S VGND VGND VPWR VPWR _3087_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3979__B1 _3495_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3050__S _3054_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5188__D _5188_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4092__D _4092_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3994__A3 _3525_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4670__A _4955_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5196__A2 _5189_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3988_ _3553_/X _3347_/X _3537_/A _3583_/X VGND VGND VPWR VPWR _3988_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_50_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4943__A2 _5118_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5727_ _5045_/A _5455_/X _5403_/X _5163_/X VGND VGND VPWR VPWR _5727_/X sky130_fd_sc_hd__a211o_1
XFILLER_109_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3286__A _3828_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5658_ _4783_/X _4398_/X _4665_/A _4672_/X _4965_/Y VGND VGND VPWR VPWR _5658_/Y
+ sky130_fd_sc_hd__o2111ai_1
XANTENNA__4156__B1 _3508_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4609_ _4243_/X _4362_/X _4910_/A _4864_/B _4364_/X VGND VGND VPWR VPWR _5746_/D
+ sky130_fd_sc_hd__o311a_2
X_5589_ _5589_/A VGND VGND VPWR VPWR _6154_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3903__B1 _3488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5105__C1 _5068_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5656__B1 _5655_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5006__A _5006_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5120__A2 _5078_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4474__A4 _4865_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5959__A1 _5680_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3682__A2 _3666_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3419__C1 _3308_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4631__A1 input11/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4631__B2 input19/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5676__A _5676_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4580__A _4580_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4919__C1 _4744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5187__A2 _5976_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4147__B1 _3218_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4698__A1 _4673_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5895__B1 _4771_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6159__CLK _6197_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4458__C _5009_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5111__A2 _4735_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5350__S _5350_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4960_ _4960_/A VGND VGND VPWR VPWR _4960_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__4622__A1 _4617_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4622__B2 _5755_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4193__C _4193_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4891_ _4891_/A VGND VGND VPWR VPWR _4891_/X sky130_fd_sc_hd__clkbuf_2
X_3911_ _3911_/A _3911_/B _3911_/C VGND VGND VPWR VPWR _4036_/C sky130_fd_sc_hd__and3_2
XANTENNA__3976__A3 _4128_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4490__A _4929_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5178__A2 _4788_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3842_ _3814_/A _3573_/X _3807_/A _4105_/A _3841_/X VGND VGND VPWR VPWR _3842_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_32_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4925__A2 _4735_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3773_ _3773_/A _3773_/B _3773_/C VGND VGND VPWR VPWR _3881_/B sky130_fd_sc_hd__and3_4
X_5512_ _6128_/Q _5504_/X _5447_/X _5511_/X VGND VGND VPWR VPWR _6128_/D sky130_fd_sc_hd__a211o_1
XFILLER_118_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4138__B1 _3709_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5443_ _5443_/A VGND VGND VPWR VPWR _6109_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4153__A3 _3515_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3834__A _4135_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5886__B1 _5237_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5374_ _5373_/Y _5371_/A _6097_/Q VGND VGND VPWR VPWR _5374_/X sky130_fd_sc_hd__a21o_1
X_4325_ _4747_/A VGND VGND VPWR VPWR _5687_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3897__C1 _3975_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3361__A1 _3254_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5638__A0 _6177_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4256_ _4307_/A _4317_/A _4246_/B _4309_/A _4255_/Y VGND VGND VPWR VPWR _4700_/A
+ sky130_fd_sc_hd__o41ai_4
XFILLER_101_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3207_ _3754_/A VGND VGND VPWR VPWR _3509_/A sky130_fd_sc_hd__buf_2
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4665__A _4665_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4310__B1 _6137_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4187_ _4520_/A _4405_/C _4859_/C _4238_/A VGND VGND VPWR VPWR _4188_/A sky130_fd_sc_hd__a31o_1
X_3138_ _4044_/B VGND VGND VPWR VPWR _3748_/A sky130_fd_sc_hd__buf_2
XANTENNA__3664__A2 _3636_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4815__D _4815_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4613__A1 _5746_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3069_ _3069_/A VGND VGND VPWR VPWR _3069_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5810__B1 _5676_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5169__A2 _5102_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4916__A2 _6138_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3447__C _3447_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4129__B1 _3762_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5877__B1 _4360_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3744__A _3744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3352__A1 _3327_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3888__C1 _3887_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4575__A _4878_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5644__A3 _5490_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3910__C _3910_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3655__A2 _3653_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5796__A2_N _4859_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5801__B1 _5145_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3407__A2 _3767_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3958__A3 _3205_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3919__A _3919_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4080__A2 _3919_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4907__A2 _4718_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6014__B _6014_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5868__B1 _4765_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3654__A _4083_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3879__C1 _3878_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3894__A2 _3183_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5291__D _6202_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4110_ _3260_/A _3708_/A _3847_/A _3509_/A VGND VGND VPWR VPWR _4110_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_68_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5090_ input27/X _4804_/X _5042_/X input11/X VGND VGND VPWR VPWR _5090_/X sky130_fd_sc_hd__a22o_2
XANTENNA__4485__A _4485_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4041_ _3679_/X _3347_/X _3533_/X _4040_/X VGND VGND VPWR VPWR _4041_/X sky130_fd_sc_hd__a31o_1
XFILLER_110_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3646__A2 _4135_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3711__C_N _3746_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4056__C1 _3302_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5399__A2 _5445_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5992_ _6200_/Q _5286_/B _5985_/B VGND VGND VPWR VPWR _5998_/A sky130_fd_sc_hd__a21boi_1
X_4943_ _5755_/D _5118_/C _4956_/D _5878_/A VGND VGND VPWR VPWR _4943_/Y sky130_fd_sc_hd__a31oi_4
XANTENNA__3803__C1 _3802_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4071__A2 _3546_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3829__A _4074_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4874_ _5240_/A _4581_/C _5903_/A _4686_/X VGND VGND VPWR VPWR _4874_/X sky130_fd_sc_hd__a31o_2
XFILLER_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3825_ _3775_/Y _3824_/Y _3562_/X VGND VGND VPWR VPWR _3825_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3756_ _3756_/A _3799_/A _3756_/C VGND VGND VPWR VPWR _3756_/X sky130_fd_sc_hd__and3_1
XANTENNA__5571__A2 _5985_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5859__B1 _4890_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3687_ _3687_/A _3687_/B VGND VGND VPWR VPWR _3687_/Y sky130_fd_sc_hd__nor2_4
X_5426_ _5424_/Y _5425_/Y _5528_/B VGND VGND VPWR VPWR _6106_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__3283__B _3815_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4531__B1 _5107_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3885__A2 _3756_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5357_ _6061_/Q _6092_/Q _5361_/S VGND VGND VPWR VPWR _5358_/A sky130_fd_sc_hd__mux2_1
X_4308_ _4308_/A VGND VGND VPWR VPWR _4308_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5288_ _5508_/A VGND VGND VPWR VPWR _5288_/X sky130_fd_sc_hd__buf_4
XANTENNA__4395__A _4395_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4239_ _5643_/B VGND VGND VPWR VPWR _4239_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4834__A1 _5102_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3637__A2 _3342_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5003__B _5003_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4047__C1 _3744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3739__A _3904_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4062__A2 _3524_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5011__A1 _4644_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4770__B1 _5188_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3474__A _4092_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5392__C _5392_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4117__A3 _3849_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input55_A memory_dmem_request_put[81] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4825__A1 _4750_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6009__B _6013_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5786__C1 _5029_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5250__A1 _5096_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4053__A2 _3362_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3800__A2 _3522_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5002__A1 _4997_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4590_ _4673_/A _4996_/A _5680_/B _4574_/A VGND VGND VPWR VPWR _4590_/X sky130_fd_sc_hd__a22o_1
X_3610_ _4105_/B _3607_/X _3608_/X _3938_/B VGND VGND VPWR VPWR _3613_/B sky130_fd_sc_hd__a22o_1
XANTENNA__3013__A0 _6025_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3564__A1 _3499_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3541_ _3891_/A VGND VGND VPWR VPWR _3541_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3384__A _3956_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3472_ _3647_/A VGND VGND VPWR VPWR _3911_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3815__C _3815_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4199__B _4718_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5211_ _5211_/A VGND VGND VPWR VPWR _5211_/X sky130_fd_sc_hd__clkbuf_4
X_6191_ _6196_/CLK _6191_/D VGND VGND VPWR VPWR _6191_/Q sky130_fd_sc_hd__dfxtp_1
X_5142_ _5136_/X _5138_/Y _4494_/X _4568_/X VGND VGND VPWR VPWR _5142_/X sky130_fd_sc_hd__a31o_1
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5069__A1 _4931_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5073_ _5073_/A VGND VGND VPWR VPWR _5078_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_84_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4816__A1 _4814_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3619__A2 _3616_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4024_ _4021_/X _4023_/Y _3508_/X _3302_/X _3866_/X VGND VGND VPWR VPWR _4024_/Y
+ sky130_fd_sc_hd__a311oi_1
XFILLER_80_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_7_0_CLK_A clkbuf_4_7_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5241__A1 _4610_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5777__C1 _4572_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5975_ _5715_/X _4390_/X _5735_/X _5974_/Y VGND VGND VPWR VPWR _5982_/A sky130_fd_sc_hd__o22ai_1
X_4926_ _4926_/A _4926_/B _4926_/C VGND VGND VPWR VPWR _4927_/A sky130_fd_sc_hd__and3_2
XANTENNA__5792__A2 _5712_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4857_ _4581_/Y _4852_/Y _4855_/Y _5732_/B VGND VGND VPWR VPWR _4857_/Y sky130_fd_sc_hd__a31oi_4
XANTENNA__3278__B _4073_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3808_ _3807_/X _3748_/C _3724_/B VGND VGND VPWR VPWR _3808_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3004__A0 _6021_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4788_ _4926_/A _4788_/B _5744_/A _5016_/A VGND VGND VPWR VPWR _5836_/A sky130_fd_sc_hd__and4_2
XANTENNA__4752__B1 _4316_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5493__B _5501_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3294__A _3802_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3739_ _3904_/A VGND VGND VPWR VPWR _4149_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_121_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5409_ _6102_/Q _5425_/B VGND VGND VPWR VPWR _5409_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5232__A1 _5230_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3469__A _3609_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5783__A2 _5176_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3243__B1 _3239_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3794__A1 _3699_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4991__B1 _5924_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5535__A2 _4333_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4743__B1 _4931_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5940__C1 _5125_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6011__C _6011_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3849__A2 _3711_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3932__A _3967_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5623__S _5627_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5471__A1 _6116_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5471__B2 _5260_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3379__A _3606_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4026__A2 _4048_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4482__B _4482_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5223__A1 _4716_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5760_ _5754_/Y _5755_/X _5759_/Y VGND VGND VPWR VPWR _5760_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5774__A2 _5773_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4711_ _4345_/X _4691_/X _4694_/X _4698_/X _4710_/Y VGND VGND VPWR VPWR _4711_/X
+ sky130_fd_sc_hd__o311a_1
X_5691_ _4570_/Y _4571_/X _5684_/Y _5690_/Y VGND VGND VPWR VPWR _5691_/Y sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__3785__A1 _3139_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4982__B1 _4981_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4642_ _4642_/A VGND VGND VPWR VPWR _4642_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4573_ _5148_/D _4332_/X _4572_/X _4378_/Y VGND VGND VPWR VPWR _4573_/X sky130_fd_sc_hd__o211a_1
XFILLER_116_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3545__C _3967_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3524_ _3583_/C VGND VGND VPWR VPWR _3524_/X sky130_fd_sc_hd__clkbuf_4
X_3455_ _3802_/D VGND VGND VPWR VPWR _3966_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_103_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3386_ _3386_/A VGND VGND VPWR VPWR _3657_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_69_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6174_ _6201_/CLK _6174_/D VGND VGND VPWR VPWR _6174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5125_ _5125_/A VGND VGND VPWR VPWR _5175_/A sky130_fd_sc_hd__buf_4
X_5056_ _4461_/X _4576_/X _4771_/X _5020_/X _5055_/X VGND VGND VPWR VPWR _5056_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_29_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4673__A _4673_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4007_ _4083_/A _3720_/A _3660_/B _3876_/X _3860_/A VGND VGND VPWR VPWR _4007_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_72_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5769__A _5924_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5462__A1 input22/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5462__B2 input14/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5214__A1 _5211_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3569__A1_N _3564_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4017__A2 _4016_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3289__A _3786_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5765__A2 _5764_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5958_ _4629_/A _4975_/X _5955_/Y _5957_/Y VGND VGND VPWR VPWR _5958_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_25_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4909_ _5757_/A VGND VGND VPWR VPWR _4984_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3776__A1 _3673_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5889_ _4823_/X _5887_/Y _5888_/X _5006_/X VGND VGND VPWR VPWR _5889_/X sky130_fd_sc_hd__o211a_2
XFILLER_21_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5517__A2 _5504_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6042__CLK _6045_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5922__C1 _4984_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5009__A _5009_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4740__A3 _4707_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6192__CLK _6196_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4256__A2 _4317_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input18_A memory_dmem_request_put[44] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3909__A_N _3286_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4008__A2 _3534_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3199__A _3891_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5205__A1 _6122_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3927__A _4048_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4731__A3 _4524_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output86_A _3129_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4758__A _4955_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5353__S _5361_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _3687_/B VGND VGND VPWR VPWR _3476_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__5141__B1 _5140_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4495__A2 _4492_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5692__A1 _4771_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3171_ _3353_/A VGND VGND VPWR VPWR _3282_/A sky130_fd_sc_hd__buf_2
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5589__A _5589_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4493__A _4623_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5995__A2 _5985_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5812_ _5097_/X _5944_/A _4671_/X _5944_/C _4657_/A VGND VGND VPWR VPWR _5813_/C
+ sky130_fd_sc_hd__a41o_1
XFILLER_34_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5743_ _5743_/A _5743_/B VGND VGND VPWR VPWR _5746_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5747__A2 _5708_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3758__A1 _3959_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6065__CLK _6203_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5755__C _5755_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5674_ _5674_/A _5674_/B _5725_/C VGND VGND VPWR VPWR _5674_/Y sky130_fd_sc_hd__nand3_1
XFILLER_30_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4625_ _4606_/Y _4607_/X _4613_/X _4622_/Y _5734_/A VGND VGND VPWR VPWR _4625_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__5904__C1 _5125_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3048__S _3054_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4556_ _4556_/A VGND VGND VPWR VPWR _4556_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5380__B1 _6098_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3930__A1 _4039_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3507_ _3478_/Y _3505_/X _4088_/C VGND VGND VPWR VPWR _3507_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4487_ _4483_/X _4485_/X _4864_/A VGND VGND VPWR VPWR _4487_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4668__A _4668_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3572__A _3572_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3438_ _3756_/A _3438_/B _4152_/C _3983_/A VGND VGND VPWR VPWR _3438_/X sky130_fd_sc_hd__or4_4
XANTENNA__5132__B1 _4241_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3369_ _4042_/A _3686_/A _3756_/C VGND VGND VPWR VPWR _3369_/X sky130_fd_sc_hd__and3_2
XANTENNA__5683__A1 _4422_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5683__B2 _5033_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ _6197_/CLK _6157_/D VGND VGND VPWR VPWR _6157_/Q sky130_fd_sc_hd__dfxtp_1
X_5108_ _5106_/X _5680_/A _4666_/A _4305_/Y VGND VGND VPWR VPWR _5108_/X sky130_fd_sc_hd__o211a_1
XFILLER_57_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3694__B1 _3208_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5499__A _5499_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6088_ _6176_/CLK _6088_/D VGND VGND VPWR VPWR _6088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5039_ _4799_/X _6053_/Q _4995_/X _5038_/Y VGND VGND VPWR VPWR _6053_/D sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__3997__A1 _3781_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5199__B1 _5198_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5738__A2 _5170_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_4_0_CLK_A clkbuf_3_5_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4410__A2 _5944_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4850__B _4974_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5910__A2 _4378_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4713__A3 _4952_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3921__A1 _3508_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4578__A _4578_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3482__A _3482_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput86 _3129_/Y VGND VGND VPWR VPWR RDY_memory_imem_request_put sky130_fd_sc_hd__buf_2
Xoutput97 _3100_/X VGND VGND VPWR VPWR memory_dmem_response_get[18] sky130_fd_sc_hd__buf_2
XFILLER_0_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_15_0_CLK_A clkbuf_3_7_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5426__A1 _5424_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4229__A2 _4513_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5977__A2 _5680_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output124_A _3022_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3988__A1 _3553_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6088__CLK _6176_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4401__A2 _4330_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3657__A _3657_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5348__S _5350_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4410_ _4398_/X _5944_/A _4403_/X _4409_/X VGND VGND VPWR VPWR _4410_/Y sky130_fd_sc_hd__a211oi_2
XANTENNA__5901__A2 _5897_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5390_ _5432_/A VGND VGND VPWR VPWR _5445_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4488__A _4878_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3912__A1 _3708_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3912__B2 _3515_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4341_ _4405_/A _4341_/B _4405_/C _4405_/D VGND VGND VPWR VPWR _4341_/Y sky130_fd_sc_hd__nand4_2
XFILLER_98_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5114__B1 _4393_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4272_ _4301_/A _4285_/B VGND VGND VPWR VPWR _4272_/X sky130_fd_sc_hd__and2_2
XFILLER_101_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5665__A1 _4873_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4468__A2 _4461_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3223_ _4065_/B VGND VGND VPWR VPWR _3223_/X sky130_fd_sc_hd__clkbuf_4
X_6011_ _6011_/A _6011_/B _6011_/C VGND VGND VPWR VPWR _6206_/D sky130_fd_sc_hd__nand3_1
XFILLER_100_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3676__B1 _3675_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3154_ _3233_/A VGND VGND VPWR VPWR _3162_/A sky130_fd_sc_hd__inv_2
XANTENNA__4625__C1 _5734_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3085_ _3096_/A VGND VGND VPWR VPWR _3094_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__3979__A1 _3660_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_5_0_CLK clkbuf_4_5_0_CLK/A VGND VGND VPWR VPWR _6155_/CLK sky130_fd_sc_hd__clkbuf_2
XANTENNA__5050__C1 _4937_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3567__A _3998_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3987_ _3357_/X _6037_/Q _3982_/X _3986_/X VGND VGND VPWR VPWR _6037_/D sky130_fd_sc_hd__a211o_1
X_5726_ _6183_/Q _5646_/X _5703_/Y _5725_/Y VGND VGND VPWR VPWR _6183_/D sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__4943__A3 _4956_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5657_ _4732_/B _4822_/X _5652_/Y _5656_/X VGND VGND VPWR VPWR _5657_/Y sky130_fd_sc_hd__o31ai_1
XANTENNA__5782__A _5782_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4156__A1 _4151_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5353__A0 _6047_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4608_ _4832_/A VGND VGND VPWR VPWR _4864_/B sky130_fd_sc_hd__buf_4
XFILLER_2_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5588_ _6154_/Q _6022_/Q _5594_/S VGND VGND VPWR VPWR _5589_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4398__A _5240_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4539_ _5079_/A _4534_/X _4538_/X VGND VGND VPWR VPWR _4539_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3903__A1 _3830_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5105__B1 _5755_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5656__A1 _4924_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5959__A2 _4891_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3682__A3 _3631_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3419__B1 _4004_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5022__A _5022_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4631__A2 _4717_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4861__A _4936_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4919__B1 _4675_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5041__C1 _4987_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3477__A _4102_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5592__A0 _6156_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4147__A1 _3533_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5396__A2_N _2986_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5344__A0 _6058_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5895__A1 _4692_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4698__A2 _4563_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3658__B1 _3657_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4607__C1 _4369_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3656__B1_N _4102_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5867__A _5899_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4622__A2 _4618_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4890_ _4890_/A _4890_/B _4890_/C _5028_/A VGND VGND VPWR VPWR _4890_/X sky130_fd_sc_hd__and4_1
XFILLER_83_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4771__A _5721_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3910_ _3910_/A _3910_/B _3910_/C VGND VGND VPWR VPWR _3910_/X sky130_fd_sc_hd__and3_1
XFILLER_51_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5032__C1 _4472_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3841_ _3841_/A _3841_/B _3593_/D VGND VGND VPWR VPWR _3841_/X sky130_fd_sc_hd__or3b_1
XFILLER_32_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3772_ _3781_/D _3966_/B VGND VGND VPWR VPWR _3773_/C sky130_fd_sc_hd__nand2_4
XANTENNA__5583__A0 _6152_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5511_ _5093_/X _4802_/X _5262_/X _5425_/B VGND VGND VPWR VPWR _5511_/X sky130_fd_sc_hd__o31a_1
XANTENNA__4138__A1 _3926_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5335__A0 _6054_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5442_ _5442_/A _5468_/B VGND VGND VPWR VPWR _5443_/A sky130_fd_sc_hd__and2_1
XANTENNA__6103__CLK _6145_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5886__A1 _4665_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5373_ _4238_/A _5805_/A _5381_/B _5369_/X VGND VGND VPWR VPWR _5373_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_99_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4324_ _4527_/A _4536_/A _4527_/C _4527_/D VGND VGND VPWR VPWR _4747_/A sky130_fd_sc_hd__a22o_2
XANTENNA__3897__B1 _3470_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5107__A _5107_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3361__A2 _4135_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5638__A1 _6045_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4946__A _4946_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3649__B1 _3749_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4255_ _4268_/A _4244_/A _4264_/C _4245_/A _4254_/Y VGND VGND VPWR VPWR _4255_/Y
+ sky130_fd_sc_hd__o41ai_4
XFILLER_47_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3206_ _3275_/B VGND VGND VPWR VPWR _3754_/A sky130_fd_sc_hd__buf_2
XANTENNA__4310__A1 _4482_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4186_ _4186_/A _6178_/Q VGND VGND VPWR VPWR _4238_/A sky130_fd_sc_hd__and2_1
X_3137_ _3687_/B VGND VGND VPWR VPWR _4044_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_55_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3664__A3 _3594_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4613__A2 _4610_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5810__A1 _6116_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3068_ _6193_/Q _6069_/Q _3072_/S VGND VGND VPWR VPWR _3069_/A sky130_fd_sc_hd__mux2_2
XANTENNA__5169__A3 _4457_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3297__A _3864_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5709_ _4838_/X _5029_/X _4385_/A _4387_/X VGND VGND VPWR VPWR _5709_/Y sky130_fd_sc_hd__a31oi_2
XANTENNA__4129__A1 _3835_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4129__B2 _3876_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5326__A0 _6186_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5877__A1 _5976_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3744__B _3744_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3352__A2 _3335_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3888__B1 _3635_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4837__C1 _4836_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4856__A _4856_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3760__A _3881_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5687__A _5687_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5801__A1 _5800_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3407__A3 _3882_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5262__C1 _5261_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3958__A4 _3543_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3812__B1 _3862_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_1_0_CLK_A clkbuf_2_1_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3000__A _5985_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6014__C _6014_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6126__CLK _6207_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6002__A2_N _5291_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5317__A0 _6182_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5868__A1 _5867_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3879__B1 _3685_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5361__S _5361_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4040_ _4073_/D _4149_/D _3998_/D _4042_/D _3543_/B VGND VGND VPWR VPWR _4040_/X
+ sky130_fd_sc_hd__o32a_2
XFILLER_68_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3646__A3 _3938_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5253__C1 _5252_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4056__B1 _3580_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5399__A3 _5395_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5991_ _6198_/Q _5570_/X _5990_/Y VGND VGND VPWR VPWR _6198_/D sky130_fd_sc_hd__a21oi_1
X_4942_ _4942_/A VGND VGND VPWR VPWR _5878_/A sky130_fd_sc_hd__buf_2
XANTENNA__3803__B1 _3962_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3200__A1_N _3134_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4873_ _4873_/A VGND VGND VPWR VPWR _5903_/A sky130_fd_sc_hd__clkbuf_4
X_3824_ _3628_/C _3674_/X _3479_/X VGND VGND VPWR VPWR _3824_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5556__B1 _5388_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3755_ _3962_/A VGND VGND VPWR VPWR _3815_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_118_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3686_ _3686_/A _3746_/B _3773_/B _3802_/A VGND VGND VPWR VPWR _3686_/X sky130_fd_sc_hd__and4_1
XFILLER_118_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5859__A1 _4777_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5425_ _6106_/Q _5425_/B VGND VGND VPWR VPWR _5425_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4531__A1 _5878_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3056__S _3056_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_4_3_0_CLK_A clkbuf_4_3_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5356_ _5356_/A VGND VGND VPWR VPWR _6091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3885__A3 _3841_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4307_ _4307_/A VGND VGND VPWR VPWR _4482_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3580__A _3580_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5287_ input5/X VGND VGND VPWR VPWR _5508_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4238_ _4238_/A VGND VGND VPWR VPWR _5643_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__4834__A2 _4831_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3637__A3 _4124_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_67_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4169_ _4169_/A _4169_/B VGND VGND VPWR VPWR _4205_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5003__C _5003_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4047__B1 _4046_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5795__B1 _5060_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6149__CLK _6197_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5011__A2 _4642_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4770__A1 _4788_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3755__A _3962_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5392__D _5438_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4586__A _4879_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input48_A memory_dmem_request_put[74] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4825__A2 _4917_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4286__B1 _6133_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4038__B1 _3990_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5786__B1 _4541_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5250__A2 _4414_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4053__A3 _3571_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5002__A2 _4789_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3013__A1 _6157_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3564__A2 _4065_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3540_ _3508_/X _3531_/X _3539_/X VGND VGND VPWR VPWR _3540_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3384__B _3956_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3471_ _3571_/C _3468_/X _3470_/X VGND VGND VPWR VPWR _3476_/C sky130_fd_sc_hd__o21a_1
XANTENNA__5880__A _5880_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5210_ _5011_/X _5209_/X _4498_/X VGND VGND VPWR VPWR _5220_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__3815__D _3975_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4199__C _4804_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6190_ _6205_/CLK _6190_/D VGND VGND VPWR VPWR _6190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5141_ _5136_/X _5138_/Y _5140_/X VGND VGND VPWR VPWR _5141_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_69_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4496__A _4520_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3721__C1 _3327_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5069__A2 _4871_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5072_ _5069_/X _5071_/X _4494_/X VGND VGND VPWR VPWR _5072_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_96_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4816__A2 _4815_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4023_ _3536_/X _3524_/X _3975_/C _3612_/D _4022_/X VGND VGND VPWR VPWR _4023_/Y
+ sky130_fd_sc_hd__a41oi_2
XFILLER_65_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4029__B1 _3476_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5777__B1 _4574_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5241__A2 _5048_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5974_ _5756_/X _5757_/X _5929_/Y _5973_/Y VGND VGND VPWR VPWR _5974_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__3788__C1 _3787_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4925_ _5123_/B _4735_/Y _4924_/X VGND VGND VPWR VPWR _4925_/Y sky130_fd_sc_hd__a21oi_1
X_4856_ _4856_/A VGND VGND VPWR VPWR _5732_/B sky130_fd_sc_hd__buf_4
X_3807_ _3807_/A _3814_/A _4044_/A VGND VGND VPWR VPWR _3807_/X sky130_fd_sc_hd__and3_1
XANTENNA__3004__A1 _6153_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4752__A1 _4750_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4787_ _4787_/A VGND VGND VPWR VPWR _5062_/A sky130_fd_sc_hd__buf_2
XFILLER_118_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3738_ _3736_/Y _3737_/X _3815_/A VGND VGND VPWR VPWR _3738_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3669_ _3447_/C _3527_/C _3278_/A _4092_/A VGND VGND VPWR VPWR _3673_/B sky130_fd_sc_hd__a31o_4
XANTENNA__3960__C1 _4002_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5408_ _5482_/A VGND VGND VPWR VPWR _5425_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__6101__D _6101_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5339_ _6056_/Q _6084_/Q _5339_/S VGND VGND VPWR VPWR _5340_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5465__C1 _5464_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5217__C1 _4556_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5768__B1 _5767_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5232__A2 _5231_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3243__A1 _3211_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3243__B2 _3241_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3794__A2 _3793_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4991__A1 _5715_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3485__A _3873_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4743__A1 _4739_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5535__A3 _5529_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5940__B1 _5905_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3849__A3 _3719_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3932__B _3932_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5471__A2 _5222_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3379__B _3432_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4026__A3 _3882_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4482__C _4985_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5759__B1 _5758_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5223__A2 _4513_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _4422_/A _4699_/X _4708_/Y _4709_/X VGND VGND VPWR VPWR _4710_/Y sky130_fd_sc_hd__o211ai_2
X_5690_ _5690_/A _5746_/A _5690_/C _5690_/D VGND VGND VPWR VPWR _5690_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__3785__A2 _3577_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4982__A1 _4975_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4982__B2 _4189_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4641_ _4855_/D _5745_/A _4843_/C _5710_/A VGND VGND VPWR VPWR _5004_/D sky130_fd_sc_hd__a31o_2
XFILLER_116_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4572_ _4643_/A VGND VGND VPWR VPWR _4572_/X sky130_fd_sc_hd__buf_2
XANTENNA__5931__B1 _5955_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3523_ _3588_/C VGND VGND VPWR VPWR _3583_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__3545__D _3700_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3454_ _3396_/X _3452_/X _3453_/X _6018_/Q _3357_/X VGND VGND VPWR VPWR _6018_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_103_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3385_ _3686_/A VGND VGND VPWR VPWR _3893_/C sky130_fd_sc_hd__clkbuf_4
X_6173_ _6176_/CLK _6173_/D VGND VGND VPWR VPWR _6173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5124_ _5124_/A _5124_/B VGND VGND VPWR VPWR _5124_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5055_ _5720_/A _5720_/B _4541_/A _4793_/X VGND VGND VPWR VPWR _5055_/X sky130_fd_sc_hd__a31o_1
XFILLER_38_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4006_ _4135_/A _3814_/A _3574_/X VGND VGND VPWR VPWR _4006_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_55_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5462__A2 _5437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4673__B _4673_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5214__A2 _4754_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5957_ _6107_/Q _4241_/X _5905_/X _5956_/X VGND VGND VPWR VPWR _5957_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_52_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3776__A2 _3674_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4908_ _4716_/X _4513_/A input39/X _5805_/B _4907_/X VGND VGND VPWR VPWR _4908_/X
+ sky130_fd_sc_hd__o311a_2
X_5888_ _5211_/X _5761_/B _4839_/Y _5020_/A VGND VGND VPWR VPWR _5888_/X sky130_fd_sc_hd__a31o_1
X_4839_ _4754_/A _4437_/A _4697_/A VGND VGND VPWR VPWR _4839_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_119_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5922__B1 _5163_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3933__C1 _3893_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_0_0_CLK_A clkbuf_3_1_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4864__A _4864_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4110__C1 _3509_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4256__A3 _4246_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4008__A3 _4006_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5205__A2 _4807_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_11_0_CLK_A clkbuf_3_5_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5913__B1 _5098_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5634__S _5638_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5141__A1 _5136_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3170_ _4004_/A _3648_/A _4065_/A VGND VGND VPWR VPWR _3170_/X sky130_fd_sc_hd__and3_1
XFILLER_67_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5692__A2 _4773_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4774__A _5073_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4404__B1 _6134_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5811_ _5811_/A _5811_/B VGND VGND VPWR VPWR _5811_/Y sky130_fd_sc_hd__nor2_1
X_5742_ _4999_/A _4378_/A _4353_/A _5741_/Y VGND VGND VPWR VPWR _5743_/A sky130_fd_sc_hd__o2bb2ai_4
XFILLER_62_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3758__A2 _3815_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5755__D _5755_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5673_ _5673_/A VGND VGND VPWR VPWR _5725_/C sky130_fd_sc_hd__buf_2
XFILLER_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4624_ _4819_/A VGND VGND VPWR VPWR _5734_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5904__B1 _5982_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5750__A1_N _6184_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4555_ _5061_/A _4555_/B _4787_/A VGND VGND VPWR VPWR _4556_/A sky130_fd_sc_hd__or3_2
XANTENNA__5380__B2 _5382_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3506_ _3828_/A VGND VGND VPWR VPWR _4088_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4668__B _4668_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4486_ _4738_/B VGND VGND VPWR VPWR _4864_/A sky130_fd_sc_hd__buf_2
XANTENNA__3930__A2 _3923_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3437_ _3437_/A _3437_/B _3437_/C VGND VGND VPWR VPWR _3438_/B sky130_fd_sc_hd__and3_2
XANTENNA__5132__B2 _5131_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3064__S _3072_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3368_ _3631_/A VGND VGND VPWR VPWR _3756_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__5683__A2 _4699_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3694__A1 _3195_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6156_ _6197_/CLK _6156_/D VGND VGND VPWR VPWR _6156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5107_ _5107_/A VGND VGND VPWR VPWR _5680_/A sky130_fd_sc_hd__buf_2
XANTENNA__4684__A _4685_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3299_ _3299_/A _3299_/B _3537_/B _3491_/A VGND VGND VPWR VPWR _3881_/A sky130_fd_sc_hd__or4b_4
X_6087_ _6176_/CLK _6087_/D VGND VGND VPWR VPWR _6087_/Q sky130_fd_sc_hd__dfxtp_1
X_5038_ _4952_/B _5012_/Y _5220_/C _5037_/Y VGND VGND VPWR VPWR _5038_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__5840__C1 _5839_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3997__A2 _3781_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5199__A1 _5174_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4159__C1 _3717_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3906__C1 _4105_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5910__A3 _4852_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3763__A _3828_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5659__C1 _4699_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3921__A2 _3917_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput87 _2979_/X VGND VGND VPWR VPWR RDY_memory_imem_response_get sky130_fd_sc_hd__buf_2
Xoutput98 _3102_/X VGND VGND VPWR VPWR memory_dmem_response_get[19] sky130_fd_sc_hd__buf_2
XFILLER_88_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input30_A memory_dmem_request_put[56] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5426__A2 _5425_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4229__A3 input33/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5977__A3 _4891_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4634__B1 _4224_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3988__A2 _3347_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output117_A _3076_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3003__A _3003_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3938__A _4042_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3657__B _3657_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5898__C1 _4403_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4769__A _4769_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3673__A _3673_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3912__A2 _3847_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4340_ _6138_/Q VGND VGND VPWR VPWR _4340_/Y sky130_fd_sc_hd__inv_2
X_4271_ _4811_/A VGND VGND VPWR VPWR _5971_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5114__A1 _5101_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3125__A0 _6051_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3222_ _3648_/B VGND VGND VPWR VPWR _4065_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__5665__A2 _4864_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6010_ _3060_/S _5291_/X _6206_/Q VGND VGND VPWR VPWR _6011_/C sky130_fd_sc_hd__a21bo_1
X_3153_ _3397_/A _3609_/B VGND VGND VPWR VPWR _3157_/C sky130_fd_sc_hd__nand2_4
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3676__A1 _3139_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4625__B1 _4613_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_67_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3084_ _3084_/A VGND VGND VPWR VPWR _3084_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3979__A2 _4004_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6032__CLK _6202_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5050__B1 _4747_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6182__CLK _6196_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3986_ _3839_/X _3986_/B _4088_/C _4088_/D VGND VGND VPWR VPWR _3986_/X sky130_fd_sc_hd__and4b_1
XFILLER_50_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5725_ _5725_/A _5725_/B _5725_/C VGND VGND VPWR VPWR _5725_/Y sky130_fd_sc_hd__nand3_2
XFILLER_22_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5656_ _4924_/X _5653_/Y _5654_/X _5655_/Y _4420_/A VGND VGND VPWR VPWR _5656_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__5889__C1 _5006_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4607_ _4459_/A _4547_/Y _4890_/C _4369_/Y VGND VGND VPWR VPWR _4607_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4156__A2 _4155_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5353__A1 _6090_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3583__A _3583_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4679__A _4924_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5587_ _5587_/A VGND VGND VPWR VPWR _6153_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4538_ _4937_/D _4536_/X _4297_/X _4882_/A VGND VGND VPWR VPWR _4538_/X sky130_fd_sc_hd__a31o_2
XANTENNA__3903__A2 _3834_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4561__C1 _4432_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5105__B2 _4971_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5105__A1 _4692_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4469_ _4457_/X _4306_/Y _4468_/Y VGND VGND VPWR VPWR _4469_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3116__A0 _6048_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5656__A2 _5653_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6139_ _6146_/CLK _6139_/D VGND VGND VPWR VPWR _6139_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5303__A _5303_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3419__B2 _3178_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3419__A1 _3831_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5959__A3 _5755_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4919__A1 _5745_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5041__B1 _6118_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5592__A1 _6024_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5973__A _5973_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4147__A2 _3967_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3493__A _3606_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4589__A _4589_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3355__B1 _3508_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input78_A memory_imem_request_put[4] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5344__A1 _6086_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5895__A2 _4960_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4698__A3 _4890_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3658__A1 _3621_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6055__CLK _6074_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_67_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4607__B1 _4890_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4851__A1_N _4799_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5804__C1 _5673_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5867__B _5899_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4622__A3 _4290_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5280__B1 _5279_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3668__A _3668_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5359__S _5361_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5032__B1 _4999_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3840_ _3828_/X _3837_/X _3839_/X VGND VGND VPWR VPWR _3840_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3387__B _3387_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5583__A1 _6020_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3771_ _3759_/X _3770_/Y _3727_/X _6026_/Q _3728_/X VGND VGND VPWR VPWR _6026_/D
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4791__C1 _4318_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5510_ _5510_/A VGND VGND VPWR VPWR _6127_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4138__A2 _4137_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5441_ _4977_/X _5412_/X _5440_/X _5398_/X _6109_/Q VGND VGND VPWR VPWR _5442_/A
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5335__A1 _6082_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3897__A1 _3882_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5886__A2 _5885_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5372_ _5508_/A VGND VGND VPWR VPWR _6011_/B sky130_fd_sc_hd__buf_4
XFILLER_99_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4323_ _4354_/B VGND VGND VPWR VPWR _4527_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__5099__B1 _5098_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4846__B1 _5133_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3649__A1 _4048_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4254_ _6136_/Q VGND VGND VPWR VPWR _4254_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5123__A _5761_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3205_ _3847_/C VGND VGND VPWR VPWR _3205_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__4310__A2 _4308_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4185_ _4405_/D VGND VGND VPWR VPWR _4859_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3136_ _3609_/A VGND VGND VPWR VPWR _3687_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_82_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3067_ _3067_/A VGND VGND VPWR VPWR _3067_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4613__A3 _4612_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5271__B1 _6062_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5810__A2 _4511_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5023__B1 _4948_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3969_ _3967_/X _3444_/X _3968_/X VGND VGND VPWR VPWR _3969_/Y sky130_fd_sc_hd__o21ai_1
X_5708_ _5145_/X _5706_/Y _5707_/Y _4924_/X VGND VGND VPWR VPWR _5708_/Y sky130_fd_sc_hd__o2bb2ai_4
XANTENNA__6104__D _6104_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4129__A2 _3305_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5326__A1 _6078_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5639_ _5639_/A VGND VGND VPWR VPWR _6177_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5877__A2 _5008_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3888__A1 _3636_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4202__A _4976_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3352__A3 _3338_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6078__CLK _6176_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4837__B1 _4834_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4872__A _4929_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5968__A _5968_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5801__A2 _4762_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5262__B1 _5045_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5687__B _5687_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3812__A1 _3238_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3488__A _4044_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5014__B1 _5013_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4773__C1 _5188_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5317__A1 _6074_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5868__A2 _4474_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3879__A1 _3517_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_4_0_CLK clkbuf_4_5_0_CLK/A VGND VGND VPWR VPWR _6045_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_68_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5878__A _5878_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5253__B1 _4393_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4056__B2 _4055_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4056__A1 _3603_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5990_ _6198_/Q _5570_/X _5288_/X VGND VGND VPWR VPWR _5990_/Y sky130_fd_sc_hd__o21ai_1
X_4941_ _4422_/X _4423_/X _4939_/Y _4940_/X VGND VGND VPWR VPWR _4941_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_91_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3803__A1 _3468_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4872_ _4929_/C VGND VGND VPWR VPWR _5240_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3398__A _3657_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3823_ _3816_/X _3820_/Y _3821_/X _6030_/Q _3822_/X VGND VGND VPWR VPWR _6030_/D
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5556__A1 _5405_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3754_ _3754_/A _3754_/B VGND VGND VPWR VPWR _3962_/A sky130_fd_sc_hd__nor2_8
XFILLER_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3685_ _3959_/D VGND VGND VPWR VPWR _3685_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5118__A _5118_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5859__A2 _4778_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5424_ input14/X _5395_/X _5405_/A VGND VGND VPWR VPWR _5424_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4516__C1 _4978_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4531__A2 _5687_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4957__A _4957_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5355_ _6048_/Q _6091_/Q _5361_/S VGND VGND VPWR VPWR _5356_/A sky130_fd_sc_hd__mux2_1
X_4306_ _4890_/B _5971_/A _4290_/Y _4305_/Y VGND VGND VPWR VPWR _4306_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_87_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5286_ _6064_/Q _5286_/B VGND VGND VPWR VPWR _5286_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__5380__A2_N _5377_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3072__S _3072_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4237_ _4229_/X _6125_/Q _4633_/S VGND VGND VPWR VPWR _4237_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5492__B1 _5491_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4168_ _4168_/A _4168_/B VGND VGND VPWR VPWR _4205_/A sky130_fd_sc_hd__nor2_1
XANTENNA__5244__B1 _5228_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4692__A _4692_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5003__D _5152_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4099_ _3668_/X _3551_/A _3418_/X _3673_/A VGND VGND VPWR VPWR _4099_/X sky130_fd_sc_hd__a211o_1
XFILLER_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4047__A1 _3477_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3119_ _6061_/Q _6092_/Q _3127_/S VGND VGND VPWR VPWR _3120_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5795__A1 _4422_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5795__B2 _5794_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5011__A3 _5010_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4770__A2 _4883_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5028__A _5028_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3730__B1 _3657_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4286__A1 _4293_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5483__B1 _5445_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3494__C1 _3588_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4038__B2 _4014_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5786__A1 _5944_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3767__A_N _3308_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3011__A _3011_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3564__A3 _3799_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3384__C _3983_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3470_ _3611_/A VGND VGND VPWR VPWR _3470_/X sky130_fd_sc_hd__buf_2
XANTENNA__5473__A1_N _4994_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4777__A _4777_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5171__C1 _5029_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2996__S _2998_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5140_ _5140_/A _5140_/B _5140_/C _5140_/D VGND VGND VPWR VPWR _5140_/X sky130_fd_sc_hd__or4_1
XANTENNA__3721__B1 _3749_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5071_ _5944_/D _4739_/X _4927_/X _5070_/Y _4403_/X VGND VGND VPWR VPWR _5071_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__5069__A3 _5068_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4022_ _3666_/X _3194_/X _3767_/B _3764_/X _3990_/X VGND VGND VPWR VPWR _4022_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__5488__A1_N _6122_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4029__A1 _4027_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5226__B1 _5013_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5777__A1 _4953_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5973_ _5973_/A _5973_/B _5973_/C VGND VGND VPWR VPWR _5973_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__5401__A _5401_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5777__B2 _5903_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4924_ _4924_/A VGND VGND VPWR VPWR _4924_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_52_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3788__B1 _3778_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4855_ _4855_/A _4996_/A _5761_/C _4855_/D VGND VGND VPWR VPWR _4855_/Y sky130_fd_sc_hd__nand4_4
X_4786_ _5061_/A VGND VGND VPWR VPWR _4786_/X sky130_fd_sc_hd__clkbuf_4
X_3806_ _3806_/A _3806_/B _3816_/D _3805_/X VGND VGND VPWR VPWR _3806_/X sky130_fd_sc_hd__or4b_1
XFILLER_118_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4752__A2 _4652_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3737_ _3519_/X _3847_/C _3756_/A _3871_/A _3911_/A VGND VGND VPWR VPWR _3737_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_20_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3960__B1 _3959_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3668_ _3668_/A VGND VGND VPWR VPWR _3668_/X sky130_fd_sc_hd__buf_2
XANTENNA__4687__A _4937_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3591__A _3591_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5407_ _5640_/D _2986_/B _5162_/A _4800_/A VGND VGND VPWR VPWR _5482_/A sky130_fd_sc_hd__a22o_1
X_3599_ _3579_/X _3598_/Y _3453_/X _6020_/Q _3541_/X VGND VGND VPWR VPWR _6020_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_102_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3712__B1 _3491_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5338_ _5338_/A VGND VGND VPWR VPWR _6083_/D sky130_fd_sc_hd__clkbuf_1
X_5269_ _5286_/B input3/X VGND VGND VPWR VPWR _5269_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5465__B1 _5540_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6116__CLK _6123_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5217__B1 _5074_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5768__A1 _6113_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3243__A2 _3215_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4991__A2 _5968_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4743__A2 _4740_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5940__A1 _5643_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3951__B1 _3950_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input60_A memory_dmem_request_put[86] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4597__A _4926_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4900__C1 _4580_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output147_A _3009_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5456__B1 _5256_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5208__B1 _4785_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5759__A1 _5756_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4482__D _4986_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5759__B2 _5739_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3785__A3 _4116_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4982__A2 _4980_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4640_ _4640_/A VGND VGND VPWR VPWR _5710_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4719__C1 _4978_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5931__A1 _5237_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4571_ _5715_/B _4859_/B _4859_/C _4800_/A VGND VGND VPWR VPWR _4571_/X sky130_fd_sc_hd__and4b_2
XANTENNA__6202__D _6202_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3522_ _3522_/A VGND VGND VPWR VPWR _3522_/X sky130_fd_sc_hd__buf_2
XFILLER_116_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5144__C1 _4555_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3453_ _4103_/C VGND VGND VPWR VPWR _3453_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4300__A _4354_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5695__B1 _4296_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6139__CLK _6146_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6172_ _6176_/CLK _6172_/D VGND VGND VPWR VPWR _6172_/Q sky130_fd_sc_hd__dfxtp_1
X_5123_ _5761_/A _5123_/B _5123_/C _5228_/A VGND VGND VPWR VPWR _5124_/B sky130_fd_sc_hd__and4_1
X_3384_ _3956_/B _3956_/C _3983_/C VGND VGND VPWR VPWR _3919_/A sky130_fd_sc_hd__or3_4
XFILLER_85_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5054_ _4865_/D _4865_/A _4937_/D _4937_/A VGND VGND VPWR VPWR _5720_/B sky130_fd_sc_hd__o211ai_4
X_4005_ _3299_/B _4124_/A _3223_/X _4004_/X _3476_/B VGND VGND VPWR VPWR _4005_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_65_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5131__A _5131_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5214__A3 _4750_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5956_ input15/X _5431_/B _5163_/X _4984_/X VGND VGND VPWR VPWR _5956_/X sky130_fd_sc_hd__a211o_1
X_5887_ _4890_/B _5761_/C _5170_/X _4923_/A _4534_/X VGND VGND VPWR VPWR _5887_/Y
+ sky130_fd_sc_hd__a32oi_2
X_4907_ input23/X _4718_/X _4906_/X _4717_/X _4978_/A VGND VGND VPWR VPWR _4907_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3586__A _3586_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4838_ _4480_/C _4437_/A _4865_/C _4937_/D VGND VGND VPWR VPWR _4838_/X sky130_fd_sc_hd__a31o_4
XFILLER_21_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4769_ _4769_/A _4769_/B _4769_/C VGND VGND VPWR VPWR _5005_/A sky130_fd_sc_hd__nand3_4
XANTENNA__6112__D _6112_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5922__A1 input13/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3933__B1 _3429_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5686__B1 _4656_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4210__A _5818_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4894__D1 _4551_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4864__B _4864_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3449__C1 _3815_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4110__B1 _3847_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4256__A4 _4309_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5976__A _5976_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4949__C1 _5973_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5610__A0 _6164_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5913__A1 _4332_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5913__B2 _4931_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3924__B1 _3860_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6022__D _6022_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5126__C1 _5175_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5141__A2 _5138_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4101__B1 _3862_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5794__A2_N _5062_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4404__A1 _4482_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5601__A0 _6160_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5810_ _6116_/Q _4511_/X _5676_/A _5809_/X VGND VGND VPWR VPWR _5811_/B sky130_fd_sc_hd__o211a_1
X_5741_ _4649_/A _4929_/C _4883_/A VGND VGND VPWR VPWR _5741_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3758__A3 _3756_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5672_ _4633_/S _4501_/X _5676_/A VGND VGND VPWR VPWR _5673_/A sky130_fd_sc_hd__a21oi_4
X_4623_ _4623_/A VGND VGND VPWR VPWR _4819_/A sky130_fd_sc_hd__buf_2
XANTENNA__5904__A1 _4794_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4554_ _4680_/A _5079_/C _4551_/Y _4552_/X _4744_/A VGND VGND VPWR VPWR _4554_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3915__B1 _3914_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3505_ _3479_/X _3483_/Y _3490_/X _3492_/X _3504_/Y VGND VGND VPWR VPWR _3505_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5668__B1 _4827_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4485_ _4485_/A VGND VGND VPWR VPWR _4485_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_89_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4668__C _4852_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3930__A3 _3925_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3436_ _3802_/B _3436_/B VGND VGND VPWR VPWR _3756_/A sky130_fd_sc_hd__nor2_4
X_3367_ _3582_/B VGND VGND VPWR VPWR _3631_/A sky130_fd_sc_hd__buf_2
XFILLER_85_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _6155_/CLK _6155_/D VGND VGND VPWR VPWR _6155_/Q sky130_fd_sc_hd__dfxtp_1
X_5106_ _5008_/X _5009_/A _4873_/A _4692_/A VGND VGND VPWR VPWR _5106_/X sky130_fd_sc_hd__a22o_2
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3694__A2 _3223_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ _6203_/CLK _6086_/D VGND VGND VPWR VPWR _6086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5037_ _4964_/X _5019_/Y _5024_/Y _4685_/X _5036_/Y VGND VGND VPWR VPWR _5037_/Y
+ sky130_fd_sc_hd__o311ai_4
X_3298_ _3353_/A VGND VGND VPWR VPWR _3491_/A sky130_fd_sc_hd__buf_2
XANTENNA__5840__B1 _5982_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5386__A_N _5383_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5199__A2 _5175_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6107__D _6107_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3841__C_N _3593_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5939_ _4679_/X _5935_/X _5937_/Y _5938_/X VGND VGND VPWR VPWR _5939_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4205__A _4205_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4159__B1 _3910_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3906__B1 _3205_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5108__C1 _4305_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4859__B _4859_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5659__B1 _4422_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4331__B1 _4329_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4875__A _4875_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput99 _3061_/X VGND VGND VPWR VPWR memory_dmem_response_get[1] sky130_fd_sc_hd__buf_2
Xoutput88 _3059_/X VGND VGND VPWR VPWR memory_dmem_response_get[0] sky130_fd_sc_hd__buf_2
XFILLER_88_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input23_A memory_dmem_request_put[49] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5831__B1 _5828_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4634__B2 _4633_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3842__C1 _3841_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6017__D _6017_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3938__B _3938_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3657__C _3657_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3070__A0 _6194_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5898__B1 _5878_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4769__B _4769_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3673__B _3673_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4570__B1 _6140_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output91_A _3087_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4270_ _4601_/A _4602_/A _4759_/A VGND VGND VPWR VPWR _4811_/A sky130_fd_sc_hd__o21ai_4
XFILLER_98_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5114__A2 _5104_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3221_ _3344_/A _3437_/C VGND VGND VPWR VPWR _3648_/B sky130_fd_sc_hd__and2_4
XFILLER_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5665__A3 _4864_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3125__A1 _6095_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3152_ _3275_/B VGND VGND VPWR VPWR _3609_/B sky130_fd_sc_hd__buf_2
XFILLER_79_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3676__A2 _3671_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4625__A1 _4606_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4625__B2 _4622_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3083_ _6184_/Q _6076_/Q _3083_/S VGND VGND VPWR VPWR _3084_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4389__B1 _4388_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5050__A1 _4777_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3985_ _3962_/X _3583_/X _3623_/B _3984_/X _3242_/X VGND VGND VPWR VPWR _3986_/B
+ sky130_fd_sc_hd__a2111o_1
XFILLER_50_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5724_ _5715_/X _4390_/X _5716_/X _5723_/Y VGND VGND VPWR VPWR _5725_/B sky130_fd_sc_hd__o22ai_1
X_5655_ _4459_/A _4461_/X _4937_/Y _5145_/A VGND VGND VPWR VPWR _5655_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__5889__B1 _5888_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4606_ _4600_/X _4605_/X _4395_/A VGND VGND VPWR VPWR _4606_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__3864__A _4083_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3583__B _3773_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4010__C1 _4009_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5586_ _6153_/Q _6021_/Q _5594_/S VGND VGND VPWR VPWR _5587_/A sky130_fd_sc_hd__mux2_1
X_4537_ _4585_/A VGND VGND VPWR VPWR _4882_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4561__B1 _4341_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3903__A3 _3902_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3075__S _3083_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5105__A2 _4328_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4468_ _4459_/X _4461_/X _4918_/A _4464_/X _4948_/A VGND VGND VPWR VPWR _4468_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5656__A3 _5654_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4695__A _4707_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3419_ _3831_/A _3418_/X _4004_/B _3178_/X _3308_/A VGND VGND VPWR VPWR _3420_/C
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3116__A1 _6091_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6207_ _6207_/CLK _6207_/D VGND VGND VPWR VPWR _6207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4399_ _4266_/A _4272_/X _4233_/A _6135_/Q VGND VGND VPWR VPWR _4442_/A sky130_fd_sc_hd__a22oi_4
X_6138_ _6146_/CLK _6138_/D VGND VGND VPWR VPWR _6138_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4077__C1 _3926_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3419__A2 _3418_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3104__A _3104_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6069_ _6074_/CLK _6069_/D VGND VGND VPWR VPWR _6069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4919__A2 _5078_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5041__A1 _4984_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3052__A0 _6043_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5973__B _5973_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4001__C1 _3562_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3355__A1 _3324_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5895__A3 _5028_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4698__A4 _5971_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4304__B1 _4543_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3658__A2 _3773_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4607__A1 _4459_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3014__A _3014_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5804__B1 _5803_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5280__A1 _5269_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5867__C _5867_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5032__A1 _4551_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3043__A0 _6039_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3770_ _3760_/X _3457_/X _3762_/X _3763_/X _3769_/X VGND VGND VPWR VPWR _3770_/Y
+ sky130_fd_sc_hd__o311ai_2
XANTENNA__4791__B1 _4738_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5440_ input17/X _5437_/X _5439_/X input9/X VGND VGND VPWR VPWR _5440_/X sky130_fd_sc_hd__a22o_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5371_ _5371_/A _6097_/Q VGND VGND VPWR VPWR _5371_/Y sky130_fd_sc_hd__nand2_1
X_4322_ _4354_/A VGND VGND VPWR VPWR _4527_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__3897__A2 _3703_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5099__A1 _5102_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4253_ _4282_/A VGND VGND VPWR VPWR _4268_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__4846__A1 _4483_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3204_ _3956_/A _3632_/A VGND VGND VPWR VPWR _3847_/C sky130_fd_sc_hd__nor2_2
XANTENNA__3649__A2 _3648_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4310__A3 _4309_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4184_ _4301_/D VGND VGND VPWR VPWR _4405_/D sky130_fd_sc_hd__buf_2
XANTENNA__5123__B _5123_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3135_ _3754_/B VGND VGND VPWR VPWR _3609_/A sky130_fd_sc_hd__inv_2
XANTENNA__4059__C1 _3867_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3066_ _6192_/Q _6068_/Q _3072_/S VGND VGND VPWR VPWR _3067_/A sky130_fd_sc_hd__mux2_2
XANTENNA__3859__A _3859_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5271__A1 _5269_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5023__A1 _4931_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3968_ _3968_/A _4042_/D _3968_/C VGND VGND VPWR VPWR _3968_/X sky130_fd_sc_hd__or3_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5707_ _4378_/A _5079_/B _4956_/A _4680_/A VGND VGND VPWR VPWR _5707_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__4782__B1 _4781_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3594__A _3594_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3899_ _3546_/X _3892_/Y _3894_/X _3898_/Y _3838_/X VGND VGND VPWR VPWR _3899_/X
+ sky130_fd_sc_hd__o311a_1
X_5638_ _6177_/Q _6045_/Q _5638_/S VGND VGND VPWR VPWR _5639_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4534__B1 _4483_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5877__A3 _5009_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4911__A1_N _2986_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5569_ _5569_/A VGND VGND VPWR VPWR _6147_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3888__A2 _3522_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6120__D _6120_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4837__A1 _4964_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5314__A _5314_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5968__B _5968_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5798__C1 _4821_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5262__A1 _4716_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5687__C _5687_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3812__A2 _3426_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5014__A1 _4633_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5984__A _6197_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4773__B1 _4353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5722__C1 _4765_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6022__CLK _6155_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3879__A2 _3869_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3009__A _3009_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6030__D _6030_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6172__CLK _6176_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5878__B _5878_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5253__A1 _5242_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3679__A _3679_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5789__C1 _5788_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4056__A2 _3300_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4940_ _4680_/X _4935_/X _5971_/D _5878_/C _4618_/X VGND VGND VPWR VPWR _4940_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_91_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3803__A2 _3746_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4871_ _4565_/A _5711_/B _4956_/D _5078_/A VGND VGND VPWR VPWR _4871_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_60_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3822_ _3822_/A VGND VGND VPWR VPWR _3822_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__6205__D _6205_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5556__A2 _5555_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3753_ _3622_/X _3734_/Y _3577_/X VGND VGND VPWR VPWR _3759_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__4303__A _4700_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3684_ _3681_/X _3683_/X _3580_/A VGND VGND VPWR VPWR _3684_/X sky130_fd_sc_hd__a21o_1
XFILLER_9_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5118__B _5118_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5859__A3 _4581_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5713__C1 _5712_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4516__B1 _4718_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5423_ _5423_/A VGND VGND VPWR VPWR _6105_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5354_ _5354_/A VGND VGND VPWR VPWR _6090_/D sky130_fd_sc_hd__clkbuf_1
X_4305_ _4347_/A _4296_/X _4378_/A VGND VGND VPWR VPWR _4305_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__5134__A _5235_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5285_ _5285_/A _5285_/B VGND VGND VPWR VPWR _5285_/X sky130_fd_sc_hd__and2_1
XFILLER_114_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4236_ _5013_/S VGND VGND VPWR VPWR _4633_/S sky130_fd_sc_hd__buf_4
XFILLER_4_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4167_ _4405_/A VGND VGND VPWR VPWR _4520_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4973__A _4973_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5492__B2 _6123_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5492__A1 _4803_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_83_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3118_ _5294_/A VGND VGND VPWR VPWR _3127_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__5244__A1 _4563_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4098_ _4105_/A _3859_/A _3704_/X _3546_/A _4097_/Y VGND VGND VPWR VPWR _4102_/B
+ sky130_fd_sc_hd__o311a_1
XANTENNA__3996__A2_N _3994_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3589__A _3611_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4047__A2 _4036_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5795__A2 _4423_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3049_ _3049_/A VGND VGND VPWR VPWR _3049_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6115__D _6115_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4755__B1 _5034_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6045__CLK _6045_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4213__A _4307_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5180__B1 _4998_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6195__CLK _6196_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3730__A1 _3437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5044__A _5044_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4883__A _4883_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4286__A2 _4246_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5483__B2 _5131_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4691__C1 _4690_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3494__B1 _3468_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3499__A _3499_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5786__A2 _4960_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6025__D _6025_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5943__C1 _5942_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3444__A1_N _3802_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3962__A _3962_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5171__B1 _5018_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3305__C_N _3475_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3721__A1 _4124_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5070_ _5096_/A _4369_/D _4843_/B _5152_/B VGND VGND VPWR VPWR _5070_/Y sky130_fd_sc_hd__o211ai_4
XANTENNA__4793__A _5903_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4021_ _4019_/X _3139_/X _3161_/X _4020_/X VGND VGND VPWR VPWR _4021_/X sky130_fd_sc_hd__a211o_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4682__C1 _5734_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4029__A2 _4028_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5226__A1 _6124_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5777__A2 _5761_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5972_ _5061_/X _5062_/X _5720_/A _5971_/Y VGND VGND VPWR VPWR _5973_/A sky130_fd_sc_hd__o211ai_1
XANTENNA__5401__B _5422_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4923_ _4923_/A VGND VGND VPWR VPWR _5123_/B sky130_fd_sc_hd__buf_2
XANTENNA__3202__A _3966_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3788__B2 _3785_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3788__A1 _3777_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6068__CLK _6202_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4854_ _4854_/A VGND VGND VPWR VPWR _5761_/C sky130_fd_sc_hd__buf_2
XFILLER_60_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4737__B1 _4736_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4785_ _4742_/A _4472_/X _4864_/A _4865_/C _4835_/A VGND VGND VPWR VPWR _4785_/X
+ sky130_fd_sc_hd__a41o_4
X_3805_ _3934_/C _3798_/Y _3800_/Y _3804_/X VGND VGND VPWR VPWR _3805_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5934__C1 _5734_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3736_ _3735_/X _3645_/A _3246_/X _3281_/A VGND VGND VPWR VPWR _3736_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_20_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4752__A3 _4751_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3960__A1 _3359_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3667_ _3870_/A _3667_/B _3966_/B VGND VGND VPWR VPWR _3668_/A sky130_fd_sc_hd__or3_4
XFILLER_69_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3598_ _3580_/X _3597_/X _3539_/X VGND VGND VPWR VPWR _3598_/Y sky130_fd_sc_hd__o21ai_1
X_5406_ input10/X _5395_/X _5405_/X VGND VGND VPWR VPWR _5406_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_102_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3712__A1 _3710_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3083__S _3083_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5337_ _6055_/Q _6083_/Q _5339_/S VGND VGND VPWR VPWR _5338_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5268_ _5570_/C VGND VGND VPWR VPWR _5286_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_102_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4219_ _4219_/A _4219_/B _4219_/C _4219_/D VGND VGND VPWR VPWR _4220_/D sky130_fd_sc_hd__nor4_1
XANTENNA__5465__A1 _5444_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5199_ _5174_/Y _5175_/X _5186_/Y _5198_/Y VGND VGND VPWR VPWR _5199_/Y sky130_fd_sc_hd__o31ai_4
XANTENNA__5217__A1 _5050_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4208__A _4282_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5768__A2 _5643_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4991__A3 _4990_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_3_0_CLK clkbuf_4_3_0_CLK/A VGND VGND VPWR VPWR _6203_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_8_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3951__A1 _3139_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5940__A2 _4501_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4878__A _4878_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5153__B1 _5240_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4900__B1 _4873_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input53_A memory_dmem_request_put[79] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5456__A1 _6112_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5456__B2 _5260_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5502__A _5502_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5208__A1 _4882_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5759__A2 _5757_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3022__A _3022_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5648__S _5648_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4719__B1 _4718_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4570_ _4800_/A _5203_/A _6140_/Q VGND VGND VPWR VPWR _4570_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_30_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3521_ _3519_/X _3520_/X _3161_/A VGND VGND VPWR VPWR _3521_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5931__A2 _5930_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3942__A1 _3940_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4788__A _4926_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3692__A _3692_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5144__B1 _4364_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3452_ _3359_/A _3408_/X _3421_/X _3450_/X _3744_/A VGND VGND VPWR VPWR _3452_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3383_ _3383_/A VGND VGND VPWR VPWR _3983_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__5695__A1 _4404_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5695__B2 _4668_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6171_ _6203_/CLK _6171_/D VGND VGND VPWR VPWR _6171_/Q sky130_fd_sc_hd__dfxtp_1
X_5122_ _5116_/Y _5119_/Y _5121_/Y _4744_/X VGND VGND VPWR VPWR _5124_/A sky130_fd_sc_hd__o2bb2ai_2
XFILLER_97_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5053_ _4437_/A _4937_/A _5152_/C _4369_/C VGND VGND VPWR VPWR _5720_/A sky130_fd_sc_hd__o211ai_4
XANTENNA__4655__C1 _4835_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5412__A _5432_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4004_ _4004_/A _4004_/B _4004_/C VGND VGND VPWR VPWR _4004_/X sky130_fd_sc_hd__and3_1
XFILLER_53_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5131__B _5444_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5214__A4 _4642_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4958__B1 _4957_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5955_ _5955_/A _5955_/B _5955_/C _5955_/D VGND VGND VPWR VPWR _5955_/Y sky130_fd_sc_hd__nand4_2
XANTENNA__3867__A _3867_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5886_ _4665_/X _5885_/X _5237_/X VGND VGND VPWR VPWR _5886_/Y sky130_fd_sc_hd__o21ai_1
X_4906_ _5438_/C _4227_/A input15/X VGND VGND VPWR VPWR _4906_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3586__B _3663_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4837_ _4964_/A _4826_/Y _4834_/Y _4836_/X VGND VGND VPWR VPWR _4837_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5907__C1 _5906_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3607__A_N _3781_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4768_ _4732_/Y _4746_/Y _4252_/X _4766_/Y _4767_/X VGND VGND VPWR VPWR _4797_/A
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__5922__A2 _5420_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3719_ _3998_/A _3719_/B VGND VGND VPWR VPWR _3720_/A sky130_fd_sc_hd__nor2_2
XANTENNA__3933__A1 _4083_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4699_ _4699_/A VGND VGND VPWR VPWR _4699_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5135__B1 _5743_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5686__A1 _5706_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4894__C1 _5034_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3697__B1 _6023_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3107__A _5294_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4864__C _4864_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3449__B1 _3448_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4110__A1 _3260_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4949__B1 _4947_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5976__B _5976_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5071__C1 _4403_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5610__A1 _6032_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5913__A2 _5080_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5374__B1 _6097_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3924__A1 _3581_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5126__B1 _5124_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3688__B1 _3687_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4101__A1 _4099_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4404__A2 _4308_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5601__A1 _6028_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3687__A _3687_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5740_ _5683_/Y _5739_/Y _4746_/A VGND VGND VPWR VPWR _5740_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_50_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5671_ _5664_/X _5670_/X _4498_/X VGND VGND VPWR VPWR _5674_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__5365__A0 _6052_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4622_ _4617_/Y _4618_/X _4290_/Y _4619_/X _5755_/B VGND VGND VPWR VPWR _4622_/Y
+ sky130_fd_sc_hd__a32oi_4
XANTENNA__5904__A2 _5903_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6106__CLK _6146_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3915__A1 _3799_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4553_ _4555_/B VGND VGND VPWR VPWR _4744_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5117__B1 _5721_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4484_ _4482_/A _4308_/X _4309_/X _6136_/Q VGND VGND VPWR VPWR _4485_/A sky130_fd_sc_hd__o31a_2
X_3504_ _3363_/X _3496_/Y _3497_/X _3502_/X _3724_/B VGND VGND VPWR VPWR _3504_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__4311__A _4405_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5668__A1 _5078_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3435_ _3315_/A _3513_/A _3345_/A VGND VGND VPWR VPWR _3732_/D sky130_fd_sc_hd__o21a_1
XFILLER_89_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4634__A1_N _4239_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3366_ _3366_/A _3440_/B VGND VGND VPWR VPWR _3582_/B sky130_fd_sc_hd__nand2_2
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _6155_/CLK _6154_/D VGND VGND VPWR VPWR _6154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5105_ _4692_/X _4328_/X _5755_/B _4971_/X _5068_/X VGND VGND VPWR VPWR _5105_/X
+ sky130_fd_sc_hd__o221a_1
X_3297_ _3864_/B VGND VGND VPWR VPWR _3537_/B sky130_fd_sc_hd__buf_2
XFILLER_57_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3694__A3 _3183_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ _6203_/CLK _6085_/D VGND VGND VPWR VPWR _6085_/Q sky130_fd_sc_hd__dfxtp_1
X_5036_ _4998_/X _5027_/X _5030_/X _5031_/X _5035_/Y VGND VGND VPWR VPWR _5036_/Y
+ sky130_fd_sc_hd__o311ai_4
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5840__A1 _4498_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3851__B1 _3868_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5053__C1 _4369_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5199__A3 _5186_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5938_ _4657_/X _5913_/X _5756_/X _5757_/X VGND VGND VPWR VPWR _5938_/X sky130_fd_sc_hd__o211a_1
XFILLER_41_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5869_ _4487_/Y _4891_/X _4931_/X _5102_/A VGND VGND VPWR VPWR _5869_/Y sky130_fd_sc_hd__a31oi_4
XANTENNA__4159__A1 _4124_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4205__B _4205_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6123__D _6123_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4159__B2 _3553_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3906__B2 _4152_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3906__A1 _3666_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5108__B1 _4666_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4859__C _4859_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4221__A _4309_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5659__A1 _5018_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4331__B2 _4330_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput89 _3082_/X VGND VGND VPWR VPWR memory_dmem_response_get[10] sky130_fd_sc_hd__buf_2
XFILLER_48_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5831__A1 _5228_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4095__B1 _4094_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input16_A memory_dmem_request_put[42] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5831__B2 _5830_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3842__B1 _4105_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4891__A _4891_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3938__C _3938_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3300__A _3881_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6129__CLK _6145_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3070__A1 _6070_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6033__D _6033_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5898__A1 _4353_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4769__C _4769_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4570__A1 _4800_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output84_A _2987_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3220_ _3461_/B VGND VGND VPWR VPWR _3437_/C sky130_fd_sc_hd__clkbuf_2
X_3151_ _3315_/A VGND VGND VPWR VPWR _3397_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3530__C1 _3529_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3676__A3 _3672_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4625__A2 _4607_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4086__B1 _4085_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3082_ _3082_/A VGND VGND VPWR VPWR _3082_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3833__B1 _3488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4389__A1 _4361_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5586__A0 _6153_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5050__A2 _4778_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3210__A _3864_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3984_ _3414_/X _3983_/X _3701_/A _3692_/A VGND VGND VPWR VPWR _3984_/X sky130_fd_sc_hd__o211a_1
X_5723_ _5719_/X _5722_/Y _4950_/X VGND VGND VPWR VPWR _5723_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5932__A1_N _5925_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5654_ _4369_/A _5867_/C _4621_/A _4999_/A VGND VGND VPWR VPWR _5654_/X sky130_fd_sc_hd__o211a_1
XFILLER_30_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5889__A1 _4823_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4605_ _4777_/A _4778_/A _4864_/A _4960_/A _4604_/X VGND VGND VPWR VPWR _4605_/X
+ sky130_fd_sc_hd__o311a_2
XANTENNA__3864__B _3864_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3583__C _3583_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4561__A1 _4340_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4010__B1 _3763_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5585_ _5618_/A VGND VGND VPWR VPWR _5594_/S sky130_fd_sc_hd__buf_2
XFILLER_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4536_ _4536_/A VGND VGND VPWR VPWR _4536_/X sky130_fd_sc_hd__buf_2
X_4467_ _4875_/A VGND VGND VPWR VPWR _4948_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4976__A _4976_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4398_ _5240_/B VGND VGND VPWR VPWR _4398_/X sky130_fd_sc_hd__clkbuf_8
X_3418_ _3588_/B VGND VGND VPWR VPWR _3418_/X sky130_fd_sc_hd__buf_2
X_6206_ _6207_/CLK _6206_/D VGND VGND VPWR VPWR _6206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3349_ _4073_/B VGND VGND VPWR VPWR _3350_/A sky130_fd_sc_hd__clkbuf_4
X_6137_ _6146_/CLK _6137_/D VGND VGND VPWR VPWR _6137_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_input8_A memory_dmem_request_put[34] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4077__B1 _4089_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6068_ _6202_/CLK _6068_/D VGND VGND VPWR VPWR _6068_/Q sky130_fd_sc_hd__dfxtp_1
X_5019_ _4931_/X _5017_/X _4870_/X _4652_/X _5018_/Y VGND VGND VPWR VPWR _5019_/Y
+ sky130_fd_sc_hd__a311oi_4
XANTENNA__3824__B1 _3479_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6118__D _6118_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5600__A _5600_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5577__A0 _6149_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4216__A _4246_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3120__A _3120_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5041__A2 _5757_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3052__A1 _6175_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5973__C _5973_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4001__B1 _4000_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3355__A2 _3352_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4304__A1 _4297_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3658__A3 _3583_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3475__A_N _3911_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_67_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4607__A2 _4547_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4068__B1 _3902_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5804__A1 _5175_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output122_A _3018_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6028__D _6028_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5280__A2 _5272_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5510__A _5510_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_83_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5032__A2 _5073_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4126__A _4126_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3579__C1 _3744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3043__A1 _6171_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4791__A1 _4243_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5740__B1 _4746_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5370_ _4189_/A _5369_/X _5381_/B VGND VGND VPWR VPWR _5371_/A sky130_fd_sc_hd__a21o_1
XFILLER_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4321_ _4942_/A VGND VGND VPWR VPWR _5687_/A sky130_fd_sc_hd__buf_2
XANTENNA__3897__A3 _3418_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5099__A2 _5097_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4252_ _4950_/A VGND VGND VPWR VPWR _4252_/X sky130_fd_sc_hd__buf_4
XFILLER_101_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4846__A2 _4485_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3203_ _3344_/A VGND VGND VPWR VPWR _3956_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3205__A _3847_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4183_ _4265_/A _4265_/C VGND VGND VPWR VPWR _4301_/D sky130_fd_sc_hd__nor2_2
XANTENNA__5123__C _5123_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4059__B1 _3362_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3134_ _3918_/A _3918_/C _4002_/A _3822_/A VGND VGND VPWR VPWR _3134_/X sky130_fd_sc_hd__or4_1
XFILLER_103_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3065_ _3065_/A VGND VGND VPWR VPWR _3065_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5420__A _5420_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5271__A2 _5270_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5023__A2 _4740_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4036__A _4036_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3967_ _3967_/A VGND VGND VPWR VPWR _3967_/X sky130_fd_sc_hd__buf_2
XFILLER_10_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4782__A1 _4457_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5706_ _5706_/A _5706_/B _5706_/C VGND VGND VPWR VPWR _5706_/Y sky130_fd_sc_hd__nand3_2
XFILLER_109_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3990__C1 _3600_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3898_ _3998_/C _3731_/D _3896_/Y _3699_/A _3897_/X VGND VGND VPWR VPWR _3898_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_5637_ _5637_/A VGND VGND VPWR VPWR _6176_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3086__S _3094_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4534__A1 _4929_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4534__B2 _4485_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5568_ _5568_/A _5568_/B VGND VGND VPWR VPWR _5569_/A sky130_fd_sc_hd__and2_1
XFILLER_117_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4519_ _5203_/A VGND VGND VPWR VPWR _5968_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__3888__A3 _3882_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5499_ _5499_/A VGND VGND VPWR VPWR _5499_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4837__A2 _4826_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3115__A _3115_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5247__C1 _5118_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5798__B1 _4744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5968__C _5968_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5209__A1_N _5207_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5330__A _5352_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5262__A2 _4513_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5014__A2 _4501_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4222__B1 _6147_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5984__B _5998_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4773__A1 _4945_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input83_A memory_imem_request_put[9] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5970__B1 _5968_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3981__C1 _3242_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5722__B1 _5973_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3879__A3 _3872_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3025__A _3025_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5878__C _5878_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5789__B1 _5673_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5240__A _5240_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5253__A2 _5245_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3803__A3 _3593_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4870_ _5018_/A VGND VGND VPWR VPWR _4870_/X sky130_fd_sc_hd__buf_4
XFILLER_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3821_ _4103_/C VGND VGND VPWR VPWR _3821_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3695__A _3695_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5961__B1 _4316_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3752_ _3744_/X _3751_/X _3727_/X _6025_/Q _3728_/X VGND VGND VPWR VPWR _6025_/D
+ sky130_fd_sc_hd__a32o_1
X_3683_ _3682_/X _3350_/X _3649_/Y VGND VGND VPWR VPWR _3683_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3972__C1 _3302_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5118__C _5118_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5713__B1 _5237_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4516__B2 input18/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4516__A1 input10/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5422_ _5422_/A _5422_/B VGND VGND VPWR VPWR _5423_/A sky130_fd_sc_hd__and2_1
X_5353_ _6047_/Q _6090_/Q _5361_/S VGND VGND VPWR VPWR _5354_/A sky130_fd_sc_hd__mux2_1
X_4304_ _4297_/X _4536_/A _5008_/A _5009_/A _4543_/A VGND VGND VPWR VPWR _4378_/A
+ sky130_fd_sc_hd__a41oi_4
XANTENNA__5415__A _5415_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5284_ _5284_/A VGND VGND VPWR VPWR _6063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4235_ _4363_/A VGND VGND VPWR VPWR _5013_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4166_ _4301_/A VGND VGND VPWR VPWR _4405_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4973__B _4973_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5492__A2 _5433_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3117_ _3117_/A VGND VGND VPWR VPWR _3117_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5244__A2 _4673_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4097_ _3512_/A _4152_/B _3573_/X _3873_/X _3470_/X VGND VGND VPWR VPWR _4097_/Y
+ sky130_fd_sc_hd__o221ai_1
XANTENNA__5150__A _5150_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3589__B _3589_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4047__A3 _4039_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3048_ _6041_/Q _6173_/Q _3054_/S VGND VGND VPWR VPWR _3049_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4999_ _4999_/A VGND VGND VPWR VPWR _5971_/C sky130_fd_sc_hd__buf_4
XANTENNA__4755__A1 _5761_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5952__B1 _4395_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5704__B1 _4652_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6131__D _6131_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5180__A1 _4871_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5325__A _5325_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3730__A2 _3446_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4286__A3 _4308_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4140__C1 _3828_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4691__B1 _5829_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3494__A1 _3592_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5786__A3 _4693_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5943__B1 _4364_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6041__D _6041_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5171__A1 _5170_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5171__B2 _4661_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5235__A _5235_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3721__A2 _3720_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4020_ _3195_/B _3829_/X _3720_/X _3489_/X _3934_/C VGND VGND VPWR VPWR _4020_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_65_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4682__B1 _4657_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5226__A2 _4807_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5971_ _5971_/A _5971_/B _5971_/C _5971_/D VGND VGND VPWR VPWR _5971_/Y sky130_fd_sc_hd__nand4_2
XFILLER_92_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4922_ _5976_/C _5971_/A _5148_/B _4708_/A VGND VGND VPWR VPWR _4922_/X sky130_fd_sc_hd__a22o_1
XFILLER_33_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3788__A2 _3638_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2996__A0 _6018_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4853_ _4317_/A _4234_/A _4255_/Y _4585_/A VGND VGND VPWR VPWR _4855_/A sky130_fd_sc_hd__o211a_4
XFILLER_60_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4737__A1 _4735_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4737__B2 _5152_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3804_ _4044_/A _4044_/B _3801_/X _3803_/X _3282_/A VGND VGND VPWR VPWR _3804_/X
+ sky130_fd_sc_hd__a311o_1
X_4784_ _4243_/X _4362_/A _4910_/A _4815_/D _4364_/A VGND VGND VPWR VPWR _5761_/A
+ sky130_fd_sc_hd__o311a_4
XANTENNA__5934__B1 _5704_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4314__A _4405_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3735_ _3780_/A _4092_/B _3904_/C _3663_/A VGND VGND VPWR VPWR _3735_/X sky130_fd_sc_hd__or4b_2
XFILLER_109_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3960__A2 _3952_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3666_ _3666_/A VGND VGND VPWR VPWR _3666_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5698__C1 _4685_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5405_ _5405_/A VGND VGND VPWR VPWR _5405_/X sky130_fd_sc_hd__buf_2
XANTENNA__5145__A _5145_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3173__B1 _3359_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3597_ _3584_/Y _3590_/X _3596_/Y VGND VGND VPWR VPWR _3597_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3712__A2 _3992_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4370__C1 _4369_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5336_ _5336_/A VGND VGND VPWR VPWR _6082_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5267_ input4/X VGND VGND VPWR VPWR _5570_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4984__A _4984_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4218_ _4218_/A _4218_/B _4218_/C _4218_/D VGND VGND VPWR VPWR _4220_/C sky130_fd_sc_hd__nor4_1
XANTENNA__5465__A2 _5445_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5198_ _5196_/Y _5197_/Y _5015_/A VGND VGND VPWR VPWR _5198_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_18_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5217__A2 _5944_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4149_ _4149_/A _4149_/B _4152_/A _4149_/D VGND VGND VPWR VPWR _4149_/X sky130_fd_sc_hd__or4_1
XFILLER_71_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4208__B _4244_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6126__D _6126_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5925__B1 _5924_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6162__CLK _6197_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4224__A _4224_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3936__C1 _3350_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4878__B _4878_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5689__C1 _5756_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3951__A2 _3946_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5153__B2 _5152_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5153__A1 _4855_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4900__A1 _4297_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4361__C1 _4360_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input46_A memory_dmem_request_put[72] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4113__C1 _3607_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5456__A2 _5222_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3303__A _4073_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5208__A2 _4461_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6036__D _6036_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5916__B1 _5976_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4719__B2 input21/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4719__A1 input13/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3520_ _3732_/D VGND VGND VPWR VPWR _3520_/X sky130_fd_sc_hd__buf_4
XANTENNA__4788__B _4788_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3942__A2 _3492_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5144__A1 _4243_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3451_ _3538_/A VGND VGND VPWR VPWR _3744_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5695__A2 _4405_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3382_ _3841_/A _4149_/D _3779_/C _3382_/D VGND VGND VPWR VPWR _3382_/X sky130_fd_sc_hd__or4_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6170_ _6203_/CLK _6170_/D VGND VGND VPWR VPWR _6170_/Q sky130_fd_sc_hd__dfxtp_1
X_5121_ _4882_/X _5118_/Y _5120_/X VGND VGND VPWR VPWR _5121_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_97_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4104__C1 _4103_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5052_ _5049_/X _4748_/X _5020_/X _5051_/Y _4665_/X VGND VGND VPWR VPWR _5052_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_84_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4655__B1 _5061_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6035__CLK _6197_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4309__A _4309_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4003_ _3867_/X _3831_/X _3512_/X _4152_/B _3934_/B VGND VGND VPWR VPWR _4003_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_37_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4958__A1 _4954_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5080__B1 _4259_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5954_ _4671_/X _5944_/C _5148_/A _4657_/X VGND VGND VPWR VPWR _5955_/C sky130_fd_sc_hd__a31o_1
XFILLER_53_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6185__CLK _6204_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5885_ _4870_/X _5859_/X _5883_/X _5884_/X VGND VGND VPWR VPWR _5885_/X sky130_fd_sc_hd__o31a_2
X_4905_ _4767_/X _4868_/X _4503_/A _4904_/Y VGND VGND VPWR VPWR _4905_/X sky130_fd_sc_hd__o211a_1
XFILLER_21_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3586__C _3876_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4044__A _4044_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4836_ _4856_/A VGND VGND VPWR VPWR _4836_/X sky130_fd_sc_hd__buf_4
XANTENNA__5907__B1 _5905_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4767_ _4767_/A VGND VGND VPWR VPWR _4767_/X sky130_fd_sc_hd__buf_4
XANTENNA__4591__C1 _4369_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4698_ _4673_/Y _4563_/A _4890_/A _5971_/D _4819_/A VGND VGND VPWR VPWR _4698_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__3933__A2 _3932_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3718_ _3410_/A _3215_/X _3482_/X _3510_/X _3717_/X VGND VGND VPWR VPWR _3718_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5135__A1 _5006_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3649_ _4048_/A _3648_/Y _3749_/B VGND VGND VPWR VPWR _3649_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__3094__S _3094_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5686__A2 _5706_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4894__B1 _4887_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3697__B2 _3541_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3697__A1 _3691_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5319_ _5365_/S VGND VGND VPWR VPWR _5328_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_0_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3449__A1 _3161_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4110__A2 _3708_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4864__D _4864_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5843__C1 _5031_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4219__A _4219_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4949__A1 _4943_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5976__C _5976_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5071__B1 _5070_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5374__A1 _5373_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3924__A2 _3882_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5126__A1 _4252_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3688__A1 _3603_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6058__CLK _6207_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5834__C1 _4440_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4101__A2 _4100_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3033__A _3033_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3968__A _3968_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3231__A_N _3226_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3687__B _3687_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4404__A3 _4309_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5670_ _4652_/X _5666_/Y _5669_/Y _5031_/X VGND VGND VPWR VPWR _5670_/X sky130_fd_sc_hd__o211a_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4621_ _4621_/A VGND VGND VPWR VPWR _5755_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__5365__A1 _6096_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4799__A _5646_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4552_ _4815_/C VGND VGND VPWR VPWR _4552_/X sky130_fd_sc_hd__buf_2
XANTENNA__4573__C1 _4378_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3915__A2 _3583_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5117__A1 _4551_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4483_ _4483_/A VGND VGND VPWR VPWR _4483_/X sky130_fd_sc_hd__clkbuf_4
X_3503_ _3537_/B VGND VGND VPWR VPWR _3724_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__4311__B _4333_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5668__A2 _5687_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3434_ _3904_/C VGND VGND VPWR VPWR _4092_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3208__A _3509_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3365_ _3461_/A _3272_/A VGND VGND VPWR VPWR _3686_/A sky130_fd_sc_hd__or2b_2
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _6155_/CLK _6153_/D VGND VGND VPWR VPWR _6153_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5423__A _5423_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5104_ _4998_/X _5102_/Y _5103_/X _4584_/X VGND VGND VPWR VPWR _5104_/X sky130_fd_sc_hd__a31o_1
X_3296_ _3799_/A VGND VGND VPWR VPWR _3299_/A sky130_fd_sc_hd__buf_2
XFILLER_58_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4628__B1 _4523_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_4_2_0_CLK clkbuf_4_3_0_CLK/A VGND VGND VPWR VPWR _6176_/CLK sky130_fd_sc_hd__clkbuf_2
X_6084_ _6202_/CLK _6084_/D VGND VGND VPWR VPWR _6084_/Q sky130_fd_sc_hd__dfxtp_1
X_5035_ _5033_/Y _5034_/X _4744_/X VGND VGND VPWR VPWR _5035_/Y sky130_fd_sc_hd__o21ai_2
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4039__A _4039_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5840__A2 _5831_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3851__A1 _4135_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5053__B1 _5152_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5937_ _5652_/Y _5936_/X _4765_/X VGND VGND VPWR VPWR _5937_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_41_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3806__D_N _3805_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5868_ _5867_/X _4474_/X _4765_/A VGND VGND VPWR VPWR _5868_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4205__C _4205_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5799_ _5732_/A _4765_/A _5973_/C _5798_/X VGND VGND VPWR VPWR _5799_/Y sky130_fd_sc_hd__a31oi_2
X_4819_ _4819_/A VGND VGND VPWR VPWR _4964_/A sky130_fd_sc_hd__buf_2
XANTENNA__4159__A2 _3844_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3906__A2 _3567_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5108__A1 _5106_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4859__D _4859_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5659__A2 _4864_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3118__A _5294_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3119__A0 _6061_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6200__CLK _6201_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4867__B1 _4863_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5816__C1 _5725_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5831__A2 _5825_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4095__A1 _3687_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3842__A1 _3814_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4412__A _4614_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5898__A2 _5021_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5508__A _5508_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3358__B1 _6017_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4570__A2 _5203_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4858__B1 _6139_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3150_ _3443_/B VGND VGND VPWR VPWR _3315_/A sky130_fd_sc_hd__buf_2
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3530__B1 _3241_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3081_ _6183_/Q _6075_/Q _3083_/S VGND VGND VPWR VPWR _3082_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4086__A1 _3975_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3272__B_N _3330_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3698__A _3749_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3833__B2 _3439_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3833__A1 _3831_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5035__B1 _4744_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4389__A2 _4370_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5586__A1 _6021_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3983_ _3983_/A _3983_/B _3983_/C VGND VGND VPWR VPWR _3983_/X sky130_fd_sc_hd__and3_2
X_5722_ _4675_/X _5720_/Y _5973_/C _4765_/A VGND VGND VPWR VPWR _5722_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__3597__B1 _3596_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5914__A2_N _5912_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5653_ _4855_/D _4673_/A _5107_/A VGND VGND VPWR VPWR _5653_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4604_ _4604_/A VGND VGND VPWR VPWR _4604_/X sky130_fd_sc_hd__buf_6
XANTENNA__5889__A2 _5887_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4322__A _4354_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5418__A _5422_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4010__A1 _3895_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5584_ _5584_/A VGND VGND VPWR VPWR _6152_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4535_ _4543_/A VGND VGND VPWR VPWR _4937_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__4116__C_N _3911_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4561__A2 _5818_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4466_ _4835_/A VGND VGND VPWR VPWR _4875_/A sky130_fd_sc_hd__buf_2
XANTENNA__4849__B1 _4837_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4397_ _5188_/B VGND VGND VPWR VPWR _5240_/B sky130_fd_sc_hd__clkbuf_2
X_3417_ _3781_/A VGND VGND VPWR VPWR _3588_/B sky130_fd_sc_hd__buf_2
X_6205_ _6205_/CLK _6205_/D VGND VGND VPWR VPWR _6205_/Q sky130_fd_sc_hd__dfxtp_1
X_3348_ _3687_/A VGND VGND VPWR VPWR _4073_/B sky130_fd_sc_hd__buf_2
XANTENNA__3521__B1 _3161_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6136_ _6146_/CLK _6136_/D VGND VGND VPWR VPWR _6136_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ _3279_/A VGND VGND VPWR VPWR _3359_/C sky130_fd_sc_hd__buf_4
XANTENNA__4077__A1 _3195_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4077__B2 _3835_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6067_ _6074_/CLK _6067_/D VGND VGND VPWR VPWR _6067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5018_ _5018_/A _5018_/B _5018_/C _5018_/D VGND VGND VPWR VPWR _5018_/Y sky130_fd_sc_hd__nor4_4
XFILLER_54_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3824__A1 _3628_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5026__B1 _4472_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5577__A1 _6016_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6134__D _6134_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5041__A3 _5757_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4001__A1 _3376_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4232__A input1/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4304__A2 _4536_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5998__A _5998_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4068__A1 _3893_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5265__B1 _5264_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5804__A2 _5797_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4407__A _4926_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output115_A _3071_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3311__A _3461_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5017__B1 _5899_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_83_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3579__B1 _3578_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4126__B _4126_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6044__D _6044_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4776__C1 _4811_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4791__A2 _4482_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5740__A1 _5683_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4320_ _4566_/A VGND VGND VPWR VPWR _4942_/A sky130_fd_sc_hd__buf_2
XANTENNA__3751__B1 _3750_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5099__A3 _5102_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4251_ _4584_/A VGND VGND VPWR VPWR _4950_/A sky130_fd_sc_hd__buf_2
XFILLER_4_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4846__A3 _5028_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3202_ _3966_/B VGND VGND VPWR VPWR _4135_/B sky130_fd_sc_hd__buf_2
XFILLER_67_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4182_ _4231_/A _4231_/B _4231_/C _4231_/D VGND VGND VPWR VPWR _4265_/C sky130_fd_sc_hd__nand4_4
XANTENNA__5123__D _5228_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_67_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4059__A1 _3832_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5701__A _5772_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3133_ _3918_/B VGND VGND VPWR VPWR _3822_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3064_ _6191_/Q _6067_/Q _3072_/S VGND VGND VPWR VPWR _3065_/A sky130_fd_sc_hd__mux2_2
XANTENNA__4317__A _4317_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3221__A _3344_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4036__B _4036_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3966_ _4042_/A _3966_/B _3966_/C VGND VGND VPWR VPWR _4105_/C sky130_fd_sc_hd__or3_4
XANTENNA__5023__A3 _5782_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4782__A2 _4771_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5705_ _5683_/Y _5704_/X _4950_/X VGND VGND VPWR VPWR _5705_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3990__B1 _3657_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5148__A _5148_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3897_ _3882_/C _3703_/A _3418_/X _3470_/X _3975_/B VGND VGND VPWR VPWR _3897_/X
+ sky130_fd_sc_hd__a311o_1
X_5636_ _6176_/Q _6044_/Q _5638_/S VGND VGND VPWR VPWR _5637_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4534__A2 _4754_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4987__A _6146_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5567_ _4199_/X _5433_/A _4803_/X _5499_/X _6147_/Q VGND VGND VPWR VPWR _5568_/A
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3891__A _3891_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3742__B1 _3741_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4518_ _4518_/A VGND VGND VPWR VPWR _5203_/A sky130_fd_sc_hd__buf_2
X_5498_ _5529_/A VGND VGND VPWR VPWR _5498_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4449_ _4422_/X _4423_/X _4431_/X _5712_/C _4448_/X VGND VGND VPWR VPWR _4449_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__6119__CLK _6147_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5247__B1 _4843_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6129__D _6129_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ _6147_/CLK _6119_/D VGND VGND VPWR VPWR _6119_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5798__A1 _4786_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5611__A _5611_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4227__A _4227_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5262__A3 input36/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3131__A _3538_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4222__A1 _5757_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4773__A2 _4852_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5970__A1 _4629_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3981__B1 _3980_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5970__B2 _5969_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3442__A_N _3272_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5183__C1 _5170_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5722__A1 _4675_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input76_A memory_imem_request_put[2] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3306__A _3687_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5238__B1 _5237_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6039__D _6039_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5789__A1 _5175_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5240__B _5240_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5878__D _5971_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3820_ _3760_/X _3457_/X _3762_/X _3763_/X _3819_/X VGND VGND VPWR VPWR _3820_/Y
+ sky130_fd_sc_hd__o311ai_2
XFILLER_60_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3695__B _3695_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3751_ _3748_/X _3749_/X _3635_/X _3750_/Y VGND VGND VPWR VPWR _3751_/X sky130_fd_sc_hd__a31o_1
XFILLER_32_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5961__A1 _5076_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3972__B1 _3762_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3682_ _3668_/X _3666_/A _3631_/X _3749_/C VGND VGND VPWR VPWR _3682_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5118__D _5118_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5713__A1 _5708_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4516__A2 _4717_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5421_ input13/X _5412_/X _5431_/B _5398_/X _6105_/Q VGND VGND VPWR VPWR _5422_/A
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4921__C1 _5734_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5352_ _5352_/A VGND VGND VPWR VPWR _5361_/S sky130_fd_sc_hd__buf_2
XFILLER_114_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4303_ _4700_/A VGND VGND VPWR VPWR _4543_/A sky130_fd_sc_hd__buf_2
XFILLER_102_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3216__A _3275_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5283_ _5285_/B _6014_/B _5283_/C VGND VGND VPWR VPWR _5284_/A sky130_fd_sc_hd__and3_1
XANTENNA__5477__B1 _5093_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4234_ _4234_/A VGND VGND VPWR VPWR _4363_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4165_ input1/X VGND VGND VPWR VPWR _4301_/A sky130_fd_sc_hd__buf_2
XANTENNA__5492__A3 _5490_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_83_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5229__B1 _4685_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3116_ _6048_/Q _6091_/Q _3116_/S VGND VGND VPWR VPWR _3117_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5431__A _5431_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5244__A3 _5878_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5150__B _5150_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4096_ _3340_/X _4090_/X _4091_/Y _3707_/X _4095_/Y VGND VGND VPWR VPWR _4096_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_82_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3047_ _3047_/A VGND VGND VPWR VPWR _3047_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4988__C1 _4987_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5577__S _5583_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4998_ _5006_/A VGND VGND VPWR VPWR _4998_/X sky130_fd_sc_hd__buf_4
XFILLER_51_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4755__A2 _4437_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5952__A1 _5721_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3949_ _4124_/B _3720_/A _3701_/A _3369_/X VGND VGND VPWR VPWR _3949_/Y sky130_fd_sc_hd__a211oi_1
XANTENNA__3097__S _3105_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3963__B1 _3468_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5704__A1 _4474_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5165__C1 _5164_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5619_ _6168_/Q _6036_/Q _5627_/S VGND VGND VPWR VPWR _5620_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5180__A2 _5706_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3715__B1 _3714_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5606__A _5606_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4510__A _5648_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3126__A _3126_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4286__A4 _4246_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4140__B1 _3142_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6091__CLK _6204_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4691__A1 _4686_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3494__A2 _3462_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5341__A _5352_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4979__C1 _4978_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5943__A1 _5093_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3954__B1 _4004_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4903__C1 _4902_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4420__A _4420_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3706__B1 _3661_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5171__A2 _5971_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3036__A _3036_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5459__B1 _5451_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4131__B1 _3663_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4682__A1 _4679_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4682__B2 _4681_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5255__A1_N _6059_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3890__C1 _3889_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5970_ _4629_/A _4975_/X _5968_/X _5969_/Y VGND VGND VPWR VPWR _5970_/X sky130_fd_sc_hd__o22a_1
X_4921_ _4916_/X _4812_/X _4917_/X _4920_/X _5734_/A VGND VGND VPWR VPWR _4934_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_45_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4852_ _4852_/A _5048_/A _4852_/C _4878_/C VGND VGND VPWR VPWR _4852_/Y sky130_fd_sc_hd__nand4_4
XFILLER_60_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2996__A1 _6150_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3803_ _3468_/A _3746_/A _3593_/D _3962_/A _3802_/X VGND VGND VPWR VPWR _3803_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__4737__A2 _4610_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4783_ _4864_/C VGND VGND VPWR VPWR _4783_/X sky130_fd_sc_hd__buf_4
XANTENNA__4314__B _4341_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5934__A1 _4785_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3945__B1 _3319_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3734_ _3238_/X _3733_/Y _3680_/X VGND VGND VPWR VPWR _3734_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5147__C1 _5032_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3665_ _3646_/X _3656_/X _3664_/Y _3562_/X _3744_/A VGND VGND VPWR VPWR _3665_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4330__A _4602_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5698__B1 _5664_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3960__A3 _3953_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5404_ _4232_/B _4859_/B _4232_/D _5403_/X VGND VGND VPWR VPWR _5405_/A sky130_fd_sc_hd__a31o_1
XANTENNA__3173__A1 _3161_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3596_ _3593_/X _3595_/X _3724_/B VGND VGND VPWR VPWR _3596_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3712__A3 _3711_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4370__B1 _4364_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5335_ _6054_/Q _6082_/Q _5339_/S VGND VGND VPWR VPWR _5336_/A sky130_fd_sc_hd__mux2_1
X_5266_ _6061_/Q _5166_/A _4224_/X _5265_/X VGND VGND VPWR VPWR _6061_/D sky130_fd_sc_hd__a22o_1
X_4217_ _4217_/A _4217_/B _4217_/C _4217_/D VGND VGND VPWR VPWR _4220_/B sky130_fd_sc_hd__nor4_1
XANTENNA__5465__A3 _5772_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4122__B1 _4121_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5870__B1 _5868_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5197_ _4420_/X _4464_/X _4793_/X _5176_/X _4685_/A VGND VGND VPWR VPWR _5197_/Y
+ sky130_fd_sc_hd__a41oi_1
X_4148_ _3695_/A _4143_/X _4144_/X _4146_/Y _4147_/X VGND VGND VPWR VPWR _4148_/X
+ sky130_fd_sc_hd__a32o_1
X_4079_ _4124_/A _4077_/Y _3223_/X _3517_/X _4078_/X VGND VGND VPWR VPWR _4079_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_16_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4208__C _4264_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5925__A1 _5915_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3936__B1 _3543_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6142__D _6142_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5138__C1 _5137_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4878__C _4878_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5689__B1 _4882_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3951__A3 _3947_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4240__A _5648_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5336__A _5336_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5153__A2 _5034_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4900__A2 _4536_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4361__B1 _4353_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4113__B1 _3589_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input39_A memory_dmem_request_put[65] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5861__B1 _4765_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3872__C1 _3871_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5208__A3 _4931_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4415__A _4415_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5916__A1 _5140_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4719__A2 _4717_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6052__D _6052_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5129__C1 _4987_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4788__C _5744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5144__A2 _4362_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3450_ _4102_/A _3426_/X _3431_/Y _3340_/X _3449_/Y VGND VGND VPWR VPWR _3450_/X
+ sky130_fd_sc_hd__o311a_1
X_3381_ _4034_/B VGND VGND VPWR VPWR _4149_/D sky130_fd_sc_hd__buf_2
X_5120_ _5711_/B _5078_/D _5667_/B _5152_/D VGND VGND VPWR VPWR _5120_/X sky130_fd_sc_hd__a211o_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5051_ _5123_/B _4735_/Y _5050_/Y _4736_/Y VGND VGND VPWR VPWR _5051_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_85_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4278__A2_N _4268_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4104__B1 _4088_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5852__B1 _4572_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4655__A1 _4333_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4002_ _4002_/A _4002_/B _4001_/X VGND VGND VPWR VPWR _4002_/X sky130_fd_sc_hd__or3b_1
XANTENNA__3863__C1 _4039_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3213__B _3440_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5080__A1 _4864_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4958__A2 _4956_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5953_ _5951_/X _4957_/X _5952_/X VGND VGND VPWR VPWR _5955_/B sky130_fd_sc_hd__a21o_1
X_5884_ _5878_/A _4956_/D _5829_/A _5878_/C _4618_/X VGND VGND VPWR VPWR _5884_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4325__A _4747_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4904_ _4881_/Y _4889_/X _4685_/X _4903_/Y VGND VGND VPWR VPWR _4904_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4044__B _4044_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4835_ _4835_/A VGND VGND VPWR VPWR _4856_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5907__A1 _6104_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5368__C1 _4188_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5132__A1_N _5129_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4766_ _4749_/X _4752_/X _4763_/Y _4765_/X VGND VGND VPWR VPWR _4766_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__4591__B1 _4572_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3717_ _4048_/A VGND VGND VPWR VPWR _3717_/X sky130_fd_sc_hd__clkbuf_2
X_4697_ _4697_/A VGND VGND VPWR VPWR _5971_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5135__A2 _4878_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3648_ _3648_/A _3648_/B VGND VGND VPWR VPWR _3648_/Y sky130_fd_sc_hd__nand2_2
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5686__A3 _5706_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3579_ _3547_/X _3560_/X _3562_/X _3578_/Y _3744_/A VGND VGND VPWR VPWR _3579_/X
+ sky130_fd_sc_hd__a311o_2
XANTENNA__5590__S _5594_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4894__A1 _4843_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5318_ _5318_/A VGND VGND VPWR VPWR _6074_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3697__A2 _3290_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3735__D_N _3663_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5700__A1_N _6182_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5249_ _4547_/Y _5246_/Y _5247_/X _5248_/X VGND VGND VPWR VPWR _5249_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__3404__A _3437_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5843__B1 _5842_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3449__A2 _3439_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4219__B _4219_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6137__D _6137_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4949__A2 _4944_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5071__A1 _5944_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4971__A1_N _4297_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4235__A _4363_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5374__A2 _5371_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3924__A3 _3674_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5126__A2 _5124_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4334__B1 _6137_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3688__A2 _3686_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5834__B1 _4827_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4098__C1 _4097_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output145_A _3005_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6047__D _6047_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3968__B _4042_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4620_ _4640_/A VGND VGND VPWR VPWR _4621_/A sky130_fd_sc_hd__buf_2
XANTENNA__4022__C1 _3990_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4551_ _4551_/A _4692_/A VGND VGND VPWR VPWR _4551_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__4573__B1 _4572_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3915__A3 _3594_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5117__A2 _4996_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3502_ _4083_/C _3457_/X _3501_/Y _3428_/X VGND VGND VPWR VPWR _3502_/X sky130_fd_sc_hd__o31a_1
X_4482_ _4482_/A _4482_/B _4985_/A _4986_/A VGND VGND VPWR VPWR _4483_/A sky130_fd_sc_hd__nor4_4
XANTENNA__4311__C _4313_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5668__A3 _5003_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3433_ _3904_/B VGND VGND VPWR VPWR _3660_/B sky130_fd_sc_hd__buf_2
XANTENNA__5522__C1 _5521_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _6197_/CLK _6152_/D VGND VGND VPWR VPWR _6152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5103_ _5048_/X _5018_/D _5944_/B _4757_/X VGND VGND VPWR VPWR _5103_/X sky130_fd_sc_hd__a31o_1
X_3364_ _4034_/A VGND VGND VPWR VPWR _4042_/A sky130_fd_sc_hd__buf_2
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3224__A _3226_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3295_ _3983_/A VGND VGND VPWR VPWR _3799_/A sky130_fd_sc_hd__buf_2
XFILLER_85_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6083_ _6202_/CLK _6083_/D VGND VGND VPWR VPWR _6083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5825__B1 _5824_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5034_ _5971_/C _5034_/B _5034_/C VGND VGND VPWR VPWR _5034_/X sky130_fd_sc_hd__and3_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4039__B _4039_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4628__B2 _4627_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6152__CLK _6197_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3851__A2 _3659_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5053__A1 _4437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5936_ _5097_/X _4917_/A _4708_/A _4610_/X _4823_/X VGND VGND VPWR VPWR _5936_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_53_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3064__A0 _6191_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5867_ _5899_/A _5899_/C _5867_/C VGND VGND VPWR VPWR _5867_/X sky130_fd_sc_hd__and3_1
XANTENNA__4205__D _4205_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6002__B1 _5293_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4818_ _5140_/A _5976_/A _4456_/X _4817_/Y VGND VGND VPWR VPWR _4818_/X sky130_fd_sc_hd__o31a_1
X_5798_ _4786_/X _5062_/A _4744_/A _4821_/Y VGND VGND VPWR VPWR _5798_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4013__C1 _4012_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4749_ _4551_/Y _5976_/B _5123_/C _5755_/D _4748_/X VGND VGND VPWR VPWR _4749_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_31_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5086__A1_N _6054_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5108__A2 _5680_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5659__A3 _4865_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3119__A1 _6092_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4867__A1 _4858_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4867__B2 _4866_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4723__A2_N _4721_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5816__B1 _5815_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3134__A _3918_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4095__A2 _4093_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3842__A2 _3573_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5039__A1_N _4799_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3358__A1 _3287_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4412__B _4543_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5898__A3 _5192_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6025__CLK _6045_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3358__B2 _3357_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3309__A _3956_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4858__A1 _4859_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6175__CLK _6201_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3530__A1 _3521_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3080_ _3080_/A VGND VGND VPWR VPWR _3080_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3044__A _3044_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5807__B1 _5769_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4086__A2 _4083_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3833__A2 _3975_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5035__A1 _5033_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3046__A0 _6040_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3982_ _4088_/C _3976_/X _3982_/C _4088_/D VGND VGND VPWR VPWR _3982_/X sky130_fd_sc_hd__and4bb_1
X_5721_ _5721_/A _5721_/B _5721_/C VGND VGND VPWR VPWR _5973_/C sky130_fd_sc_hd__nand3_2
XANTENNA__3597__A1 _3584_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5652_ _5026_/X _5680_/C _4823_/X VGND VGND VPWR VPWR _5652_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_31_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4603_ _4329_/X _4330_/X _4728_/A _4462_/A VGND VGND VPWR VPWR _4604_/A sky130_fd_sc_hd__o211ai_4
X_5583_ _6152_/Q _6020_/Q _5583_/S VGND VGND VPWR VPWR _5584_/A sky130_fd_sc_hd__mux2_1
X_4534_ _4929_/C _4754_/A _4483_/X _4485_/X VGND VGND VPWR VPWR _4534_/X sky130_fd_sc_hd__o22a_2
XANTENNA__3219__A _3387_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4010__A2 _3760_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4849__B2 _4848_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4849__A1 _4685_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4465_ _4340_/Y _4209_/A _4341_/Y VGND VGND VPWR VPWR _4835_/A sky130_fd_sc_hd__o21a_2
X_4396_ _4734_/A VGND VGND VPWR VPWR _5188_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_89_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3416_ _3680_/A VGND VGND VPWR VPWR _4036_/A sky130_fd_sc_hd__buf_4
X_6204_ _6204_/CLK _6204_/D VGND VGND VPWR VPWR _6204_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3347_ _3499_/A VGND VGND VPWR VPWR _3347_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3521__A1 _3519_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6135_ _6146_/CLK _6135_/D VGND VGND VPWR VPWR _6135_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _6203_/CLK _6066_/D VGND VGND VPWR VPWR _6066_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ _4565_/A _4668_/B _4852_/C _5899_/C VGND VGND VPWR VPWR _5017_/X sky130_fd_sc_hd__a31o_2
X_3278_ _3278_/A _4073_/C VGND VGND VPWR VPWR _3279_/A sky130_fd_sc_hd__nor2_1
XANTENNA__4077__A2 _3831_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3824__A2 _3674_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5026__A1 _4437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3037__A0 _6036_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4785__B1 _4835_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5919_ _5028_/X _5880_/X _5779_/X _4374_/X VGND VGND VPWR VPWR _5919_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5609__A _5609_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6048__CLK _6205_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4513__A _4513_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6010__B1_N _6206_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4232__B _4232_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4001__A2 _3996_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6198__CLK _6201_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6150__D _6150_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4304__A3 _5008_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5998__B _5998_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4068__A2 _3653_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3799__A _3799_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input21_A memory_dmem_request_put[47] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5265__A1 _4801_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5017__A1 _4565_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3311__B _3311_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_83_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3028__A0 _6032_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3579__A1 _3547_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output108_A _3122_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4776__B1 _4640_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4791__A3 _4247_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4423__A _4699_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5519__A _5519_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_1_0_CLK clkbuf_4_1_0_CLK/A VGND VGND VPWR VPWR _6197_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_32_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6060__D _6060_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5740__A2 _5739_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3200__B1 _6016_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3751__A1 _3748_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4250_ _4243_/X _4654_/A _4910_/A _5756_/A VGND VGND VPWR VPWR _4584_/A sky130_fd_sc_hd__o31a_4
XFILLER_101_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3201_ _3330_/A _3442_/B VGND VGND VPWR VPWR _3966_/B sky130_fd_sc_hd__and2b_4
X_4181_ _4219_/C _4219_/D VGND VGND VPWR VPWR _4231_/D sky130_fd_sc_hd__nor2_1
XFILLER_95_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3132_ input3/X VGND VGND VPWR VPWR _3918_/B sky130_fd_sc_hd__clkinv_2
XFILLER_67_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4059__A2 _3583_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3267__B1 _3266_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5701__B _5772_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3063_ _3096_/A VGND VGND VPWR VPWR _3072_/S sky130_fd_sc_hd__buf_2
XANTENNA__3221__B _3437_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3019__A0 _6028_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4036__C _4036_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3965_ _3871_/B _3457_/A _4073_/D VGND VGND VPWR VPWR _3965_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_50_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3896_ _3895_/X _3457_/A _3403_/X _3410_/A _3537_/A VGND VGND VPWR VPWR _3896_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_5704_ _4474_/X _5661_/B _4652_/A VGND VGND VPWR VPWR _5704_/X sky130_fd_sc_hd__a21o_2
XANTENNA__4333__A _4333_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5429__A _5429_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3990__A1 _3397_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3990__B2 _3582_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5148__B _5148_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4782__A3 _4773_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5635_ _5635_/A VGND VGND VPWR VPWR _6175_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5192__B1 _5899_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5566_ _5566_/A VGND VGND VPWR VPWR _6146_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3742__A1 _3534_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4517_ _4716_/A _4513_/X input34/X _5805_/B _4516_/X VGND VGND VPWR VPWR _4522_/A
+ sky130_fd_sc_hd__o311ai_4
X_5497_ _5201_/X _5405_/X _5224_/Y _5288_/X _5496_/X VGND VGND VPWR VPWR _6124_/D
+ sky130_fd_sc_hd__o311ai_1
X_4448_ _4437_/Y _4440_/Y _5903_/B _5079_/C _5020_/A VGND VGND VPWR VPWR _4448_/X
+ sky130_fd_sc_hd__a221o_2
X_4379_ _4379_/A VGND VGND VPWR VPWR _4462_/A sky130_fd_sc_hd__buf_2
XFILLER_58_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5247__A1 _4347_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ _6147_/CLK _6118_/D VGND VGND VPWR VPWR _6118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5798__A2 _5062_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6049_ _6205_/CLK _6049_/D VGND VGND VPWR VPWR _6049_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4508__A _5805_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3412__A _3582_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6145__D _6145_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4222__A2 _4985_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4243__A _4243_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3981__A1 _3628_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5970__A2 _4975_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5183__B1 _5903_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5722__A2 _5720_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3733__A1 _3731_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input69_A memory_dmem_request_put[95] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4694__C1 _4290_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3497__B1 _3571_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5238__A1 _5232_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5789__A2 _5784_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5240__C _5240_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4997__B1 _4736_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3322__A _3589_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5013__S _5013_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6055__D _6055_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5928__A2_N _4604_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4749__B1 _4748_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3695__C _3695_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3421__B1 _3420_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3750_ _3537_/X _3716_/X _3816_/A VGND VGND VPWR VPWR _3750_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5961__A2 _4971_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3972__A1 _3142_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3992__A _3992_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3681_ _3830_/D _3429_/X _3679_/X _3645_/Y _3680_/X VGND VGND VPWR VPWR _3681_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__3972__B2 _3300_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5174__B1 _5172_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5713__A2 _5709_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5420_ _5420_/A VGND VGND VPWR VPWR _5431_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__4921__B1 _4920_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5351_ _5351_/A VGND VGND VPWR VPWR _6089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4302_ _4354_/B VGND VGND VPWR VPWR _5009_/A sky130_fd_sc_hd__buf_2
X_5282_ _5985_/A _3822_/A _5272_/Y _5279_/Y VGND VGND VPWR VPWR _5283_/C sky130_fd_sc_hd__o211ai_1
XFILLER_102_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4233_ _4233_/A VGND VGND VPWR VPWR _4234_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_4_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5477__A1 _6118_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5477__B2 _4802_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5712__A _5712_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5229__A1 _4894_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4164_ _4157_/X _4163_/Y _3290_/X _6045_/Q _3891_/X VGND VGND VPWR VPWR _6045_/D
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4328__A _5667_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_83_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4095_ _3687_/Y _4093_/X _4094_/X VGND VGND VPWR VPWR _4095_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3115_ _3115_/A VGND VGND VPWR VPWR _3115_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5431__B _5431_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3232__A _3667_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5150__C _5150_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4988__B1 _6117_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3046_ _6040_/Q _6172_/Q _3054_/S VGND VGND VPWR VPWR _3047_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5244__A4 _4692_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4997_ _5976_/C _5102_/C _4736_/Y VGND VGND VPWR VPWR _4997_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_11_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4755__A3 _4754_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5952__A2 _4965_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3948_ _3403_/X _3519_/X _3673_/B VGND VGND VPWR VPWR _3948_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3963__A1 _3867_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4998__A _5006_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3879_ _3517_/X _3869_/Y _3872_/X _3685_/X _3878_/Y VGND VGND VPWR VPWR _3879_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__5704__A2 _5661_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5618_ _5618_/A VGND VGND VPWR VPWR _5627_/S sky130_fd_sc_hd__buf_2
XANTENNA__5165__B1 _5013_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5549_ _5523_/X _4218_/D _5529_/X _5499_/X _6141_/Q VGND VGND VPWR VPWR _5550_/A
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3715__A1 _3699_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5180__A3 _5179_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4676__C1 _4675_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3716__A2_N _3911_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5622__A _5622_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4140__A1 _3760_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4140__B2 _4139_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4691__A2 _5755_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_86_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4238__A _4238_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3142__A _3695_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4979__B1 _4718_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3954__A1 _3932_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5943__A2 _4362_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5156__B1 _5155_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4701__A _5016_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4903__B1 _5237_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3706__A1 _3701_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3317__A _3779_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5459__B2 _6113_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5459__A1 _4977_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5532__A _5532_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4131__A1 _4061_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4682__A2 _4619_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3890__B1 _3880_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4920_ _5148_/B _5148_/D _4672_/X _4919_/Y VGND VGND VPWR VPWR _4920_/X sky130_fd_sc_hd__a31o_1
XFILLER_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5919__C1 _4374_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4851_ _4799_/X _6050_/Q _4809_/X _4850_/Y VGND VGND VPWR VPWR _6050_/D sky130_fd_sc_hd__a2bb2oi_1
XFILLER_33_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3802_ _3802_/A _3802_/B _3895_/A _3802_/D VGND VGND VPWR VPWR _3802_/X sky130_fd_sc_hd__or4_4
XFILLER_60_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4782_ _4457_/X _4771_/X _4773_/Y _4781_/X VGND VGND VPWR VPWR _4782_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5934__A2 _5933_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4314__C _4518_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6109__CLK _6123_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3733_ _3731_/X _3732_/X _3528_/A VGND VGND VPWR VPWR _3733_/Y sky130_fd_sc_hd__a21boi_4
XANTENNA__3945__A1 _3666_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4611__A _4729_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5147__B1 _5102_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3664_ _3536_/X _3636_/X _3594_/X _3662_/Y _3663_/X VGND VGND VPWR VPWR _3664_/Y
+ sky130_fd_sc_hd__o311ai_1
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5698__A1 _5694_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5403_ _5757_/A VGND VGND VPWR VPWR _5403_/X sky130_fd_sc_hd__buf_2
XANTENNA__3227__A _3437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4370__A1 _4362_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3173__A2 _3170_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3595_ _3271_/A _3594_/X _3249_/X _3748_/B VGND VGND VPWR VPWR _3595_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5334_ _5334_/A VGND VGND VPWR VPWR _6081_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5265_ _4801_/X _5260_/X _5262_/X _5264_/X VGND VGND VPWR VPWR _5265_/X sky130_fd_sc_hd__a31o_1
X_5196_ _5187_/X _5189_/X _4494_/X _5195_/Y VGND VGND VPWR VPWR _5196_/Y sky130_fd_sc_hd__o211ai_4
X_4216_ _4246_/B VGND VGND VPWR VPWR _4985_/A sky130_fd_sc_hd__buf_2
XANTENNA__5442__A _5442_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4122__A1 _3357_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4122__B2 _3453_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5870__A1 _5794_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5870__B2 _5869_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4147_ _3533_/X _3967_/X _3218_/X _3621_/C VGND VGND VPWR VPWR _4147_/X sky130_fd_sc_hd__a211o_1
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5083__C1 _5082_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3432__A_N _3440_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_83_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4078_ _3679_/X _4089_/B _3919_/X _3428_/X _3488_/X VGND VGND VPWR VPWR _4078_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5588__S _5594_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4208__D _4245_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3029_ _3029_/A VGND VGND VPWR VPWR _3029_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5925__A2 _5921_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3936__A1 _3418_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5138__B1 _5732_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4521__A _4800_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5617__A _5617_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4878__D _4878_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5689__B2 _4652_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5689__A1 _5757_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5153__A3 _5240_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3137__A _3687_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4361__B2 _5140_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4361__A1 _5976_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2976__A _6100_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4113__A1 _3527_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5352__A _5352_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4088__A_N _3839_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5861__A1 _5706_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3872__B1 _3161_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5074__C1 _5078_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3600__A _3600_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5916__A2 _4840_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5377__B1 _5371_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4431__A _5706_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5129__B1 _6120_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4788__D _5016_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4888__C1 _5240_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5144__A3 _4247_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3047__A _3047_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5201__B_N _4200_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3380_ _3603_/D _3781_/B _4034_/B _3904_/C VGND VGND VPWR VPWR _3380_/X sky130_fd_sc_hd__or4_4
XFILLER_69_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3560__C1 _3559_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5050_ _4777_/A _4778_/A _4747_/A _4937_/A VGND VGND VPWR VPWR _5050_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_69_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4104__A1 _6042_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5852__A1 _5079_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4001_ _3376_/X _3996_/X _4000_/X _3562_/A VGND VGND VPWR VPWR _4001_/X sky130_fd_sc_hd__a211o_2
XANTENNA__4655__A2 _5818_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3863__B1 _3861_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5952_ _5721_/A _4965_/Y _5782_/A _4395_/A VGND VGND VPWR VPWR _5952_/X sky130_fd_sc_hd__a31o_1
XFILLER_37_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4812__C1 _5761_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5080__A2 _5008_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4903_ _4890_/X _4892_/X _5237_/A _4902_/Y VGND VGND VPWR VPWR _4903_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__3510__A _3586_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5883_ _5211_/X _5878_/B _4783_/X _4680_/A _5878_/A VGND VGND VPWR VPWR _5883_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4834_ _5102_/A _4831_/X _4833_/X _4794_/X VGND VGND VPWR VPWR _4834_/Y sky130_fd_sc_hd__o211ai_4
XANTENNA__4044__C _4044_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5907__A2 _4975_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5368__B1 input2/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4040__B1 _4042_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4765_ _4765_/A VGND VGND VPWR VPWR _4765_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__6081__CLK _6203_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4591__A1 _5971_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4341__A _4405_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3716_ _3832_/A _3911_/B _3418_/X _3674_/C VGND VGND VPWR VPWR _3716_/X sky130_fd_sc_hd__o2bb2a_2
XANTENNA__5437__A _5437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4696_ _4696_/A VGND VGND VPWR VPWR _4697_/A sky130_fd_sc_hd__buf_2
XFILLER_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5135__A3 _4852_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3647_ _3647_/A VGND VGND VPWR VPWR _4048_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3578_ _4126_/B _3569_/X _3571_/X _3576_/Y _3577_/X VGND VGND VPWR VPWR _3578_/Y
+ sky130_fd_sc_hd__a221oi_2
XFILLER_115_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4894__A2 _4565_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5317_ _6182_/Q _6074_/Q _5317_/S VGND VGND VPWR VPWR _5318_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3697__A3 _3696_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5248_ _5118_/A _5003_/B _5003_/C _5152_/D VGND VGND VPWR VPWR _5248_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5843__A1 _5176_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5179_ _5179_/A VGND VGND VPWR VPWR _5179_/X sky130_fd_sc_hd__buf_4
XFILLER_68_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3854__B1 _3853_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4219__C _4219_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5056__C1 _5055_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5071__A2 _4739_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3420__A _4036_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6153__D _6153_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5359__A0 _6049_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4031__B1 _4030_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4251__A _4584_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5347__A _5347_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4334__A1 _4293_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input51_A memory_dmem_request_put[77] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_86_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5834__A1 _5899_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4098__B1 _3546_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5295__C1 _5294_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3845__B1 _3301_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output138_A _3051_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4426__A _4759_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3330__A _3330_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3968__C _3968_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4270__B1 _4759_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4103__A_N _3286_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6063__D _6063_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4573__A1 _5148_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4022__B1 _3764_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5257__A input5/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4550_ _4769_/C VGND VGND VPWR VPWR _4692_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5770__B1 _5769_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5117__A3 _4887_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3501_ _3499_/X _3911_/C _3475_/D VGND VGND VPWR VPWR _3501_/Y sky130_fd_sc_hd__a21oi_4
X_4481_ _4642_/A VGND VGND VPWR VPWR _4665_/A sky130_fd_sc_hd__buf_2
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5668__A4 _4887_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3432_ _3440_/A _3432_/B VGND VGND VPWR VPWR _3904_/B sky130_fd_sc_hd__and2b_1
XANTENNA__5522__B1 _5447_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3363_ _3847_/B _3557_/A _3382_/D _3362_/Y _4004_/A VGND VGND VPWR VPWR _3363_/X
+ sky130_fd_sc_hd__o221a_4
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6151_ _6197_/CLK _6151_/D VGND VGND VPWR VPWR _6151_/Q sky130_fd_sc_hd__dfxtp_1
X_5102_ _5102_/A _5102_/B _5102_/C _5102_/D VGND VGND VPWR VPWR _5102_/Y sky130_fd_sc_hd__nand4_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5825__A1 _4829_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3294_ _3802_/A VGND VGND VPWR VPWR _3983_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _6202_/CLK _6082_/D VGND VGND VPWR VPWR _6082_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5825__B2 _4875_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_85_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5033_ _4786_/X _5062_/A _5721_/B _5032_/Y VGND VGND VPWR VPWR _5033_/Y sky130_fd_sc_hd__a2bb2oi_4
XANTENNA__3836__B1 _3347_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5720__A _5720_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3851__A3 _3215_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5038__C1 _5037_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5053__A2 _4937_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4336__A _4432_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3240__A _3687_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5935_ _5829_/B _4930_/X _5080_/X _5102_/B _5167_/X VGND VGND VPWR VPWR _5935_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_41_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3064__A1 _6067_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5866_ _5240_/A _5903_/A _4875_/A _4792_/A _4924_/A VGND VGND VPWR VPWR _5866_/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_61_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4817_ _4657_/A _4812_/X _4813_/X _4816_/X VGND VGND VPWR VPWR _4817_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__6002__B2 _6202_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5167__A _5167_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5797_ _5754_/Y _5792_/Y _5796_/Y VGND VGND VPWR VPWR _5797_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__4013__B1 _4036_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4748_ _5899_/B _4621_/A _5711_/A _5022_/A VGND VGND VPWR VPWR _4748_/X sky130_fd_sc_hd__a31o_2
XFILLER_5_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4679_ _4924_/A VGND VGND VPWR VPWR _4679_/X sky130_fd_sc_hd__buf_2
XANTENNA__5513__B1 _6129_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4867__A2 _4859_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3415__A _3754_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5816__A1 _4952_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6148__D _6148_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3827__B1 _3826_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3134__B _3918_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3842__A3 _3807_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3150__A _3443_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4246__A _4246_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5752__B1 _5706_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3358__A2 _3290_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5805__A _5805_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4858__A2 _5203_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3325__A _3621_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3530__A2 _3522_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5807__A1 _5676_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6058__D _6058_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5540__A _5540_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3818__B1 _3695_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4491__B1 _5240_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5035__A2 _5034_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3981_ _3628_/A _3998_/C _3977_/X _3980_/X _3242_/X VGND VGND VPWR VPWR _3982_/C
+ sky130_fd_sc_hd__a311o_2
XFILLER_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3046__A1 _6172_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5720_ _5720_/A _5720_/B VGND VGND VPWR VPWR _5720_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3597__A2 _3590_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5991__B1 _5990_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5651_ _5811_/A _5651_/B VGND VGND VPWR VPWR _5651_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4602_ _4602_/A VGND VGND VPWR VPWR _4778_/A sky130_fd_sc_hd__buf_2
X_5582_ _5582_/A VGND VGND VPWR VPWR _6151_/D sky130_fd_sc_hd__clkbuf_1
X_4533_ _4533_/A VGND VGND VPWR VPWR _4929_/C sky130_fd_sc_hd__buf_2
XANTENNA__4010__A3 _3722_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5715__A _5715_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4464_ _5903_/B VGND VGND VPWR VPWR _4464_/X sky130_fd_sc_hd__buf_4
XANTENNA__4849__A2 _4818_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6203_ _6203_/CLK _6203_/D VGND VGND VPWR VPWR _6203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3235__A _3904_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4395_ _4395_/A VGND VGND VPWR VPWR _4732_/B sky130_fd_sc_hd__buf_4
X_3415_ _3754_/B VGND VGND VPWR VPWR _3680_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3346_ _3711_/B VGND VGND VPWR VPWR _3410_/B sky130_fd_sc_hd__buf_4
XANTENNA__3521__A2 _3520_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6134_ _6146_/CLK _6134_/D VGND VGND VPWR VPWR _6134_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _6203_/CLK _6065_/D VGND VGND VPWR VPWR _6065_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _5016_/A VGND VGND VPWR VPWR _5899_/C sky130_fd_sc_hd__buf_2
XFILLER_85_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3277_ _3500_/A VGND VGND VPWR VPWR _4073_/C sky130_fd_sc_hd__clkbuf_2
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3809__B1 _3492_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3690__D1 _3689_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5026__A2 _5009_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3037__A1 _6168_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4785__A1 _4742_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5918_ _5021_/X _5167_/X _5068_/X _5880_/X VGND VGND VPWR VPWR _5918_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3993__C1 _3992_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5849_ _6190_/Q _4629_/X _4630_/X _5848_/X VGND VGND VPWR VPWR _6190_/D sky130_fd_sc_hd__o31a_1
XFILLER_22_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4232__C _4301_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3745__C1 _3594_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3129__B _6063_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3145__A _3437_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4304__A4 _5009_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5998__C _5998_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2984__A _5381_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4068__A3 _3668_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3799__B _3847_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_67_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5360__A _5360_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5265__A2 _5260_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5670__C1 _5031_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input14_A memory_dmem_request_put[40] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5017__A2 _4668_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3028__A1 _6164_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4776__A1 _4926_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3579__A2 _3560_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3984__C1 _3692_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5519__B _5531_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6142__CLK _6145_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3200__B2 _5388_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3751__A2 _3749_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5489__C1 _5488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4180_ _4219_/A _4219_/B VGND VGND VPWR VPWR _4231_/C sky130_fd_sc_hd__nor2_1
XANTENNA__3055__A _3055_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3200_ _3134_/X _3197_/X _6016_/Q _5388_/B VGND VGND VPWR VPWR _6016_/D sky130_fd_sc_hd__a2bb2o_1
X_3131_ _3538_/A VGND VGND VPWR VPWR _4002_/A sky130_fd_sc_hd__buf_2
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5270__A _5286_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5110__D1 _4574_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3267__A1 _3246_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5701__C _5701_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3062_ _5294_/A VGND VGND VPWR VPWR _3096_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3019__A1 _6160_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4036__D _4036_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4614__A _4614_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5964__B1 _5753_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3964_ _3195_/B _3194_/X _3767_/B _3687_/Y _3512_/X VGND VGND VPWR VPWR _3964_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_16_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3895_ _3895_/A VGND VGND VPWR VPWR _3895_/X sky130_fd_sc_hd__buf_4
X_5703_ _5676_/X _5702_/X _5811_/A VGND VGND VPWR VPWR _5703_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5429__B _5468_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3990__A2 _3781_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5148__C _5148_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5716__B1 _4950_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5634_ _6175_/Q _6043_/Q _5638_/S VGND VGND VPWR VPWR _5635_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5192__A1 _4404_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5565_ _5988_/A _5565_/B VGND VGND VPWR VPWR _5566_/A sky130_fd_sc_hd__or2_1
XANTENNA__5445__A _5445_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3742__A2 _3938_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4516_ input10/X _4717_/A _4718_/A input18/X _4978_/A VGND VGND VPWR VPWR _4516_/X
+ sky130_fd_sc_hd__a221o_1
X_5496_ _6124_/Q _4239_/X _5495_/X _5092_/X VGND VGND VPWR VPWR _5496_/X sky130_fd_sc_hd__a2bb2o_1
X_4447_ _4869_/A VGND VGND VPWR VPWR _5020_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4378_ _4378_/A _4673_/B _4673_/A VGND VGND VPWR VPWR _4378_/Y sky130_fd_sc_hd__nand3_4
XANTENNA_input6_A memory_dmem_request_put[32] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6117_ _6145_/CLK _6117_/D VGND VGND VPWR VPWR _6117_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5247__A2 _4369_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3329_ _4092_/A VGND VGND VPWR VPWR _4083_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4455__B1 _5756_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6048_ _6205_/CLK _6048_/D VGND VGND VPWR VPWR _6048_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3412__B _3446_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4524__A _5667_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6165__CLK _6176_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4222__A3 _4986_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5707__B1 _4956_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3981__A2 _3998_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6161__D _6161_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5183__A1 _5745_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3718__C1 _3717_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3733__A2 _3732_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4694__B1 _5179_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3497__A1 _3299_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3603__A _3603_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5238__A2 _5236_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5240__D _5240_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4997__A1 _5976_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output120_A _2993_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4434__A _4890_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4749__A1 _4551_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5946__B1 _5945_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3421__A1 _3327_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5961__A3 _4395_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6071__D _6071_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3972__A2 _3971_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3992__B _3992_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3680_ _3680_/A VGND VGND VPWR VPWR _3680_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5174__B2 _5173_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5174__A1 _5168_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4921__A1 _4916_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5350_ _6046_/Q _6089_/Q _5350_/S VGND VGND VPWR VPWR _5351_/A sky130_fd_sc_hd__mux2_1
X_4301_ _4301_/A _4405_/B _4301_/C _4301_/D VGND VGND VPWR VPWR _4354_/B sky130_fd_sc_hd__nand4_4
X_5281_ input4/X VGND VGND VPWR VPWR _5985_/A sky130_fd_sc_hd__inv_2
XFILLER_114_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4232_ input1/X _4232_/B _4301_/C _4232_/D VGND VGND VPWR VPWR _4233_/A sky130_fd_sc_hd__nand4_4
XANTENNA__5477__A2 _4239_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5712__B _5746_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6038__CLK _6202_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3513__A _3513_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4163_ _3300_/X _3807_/A _3828_/X _4162_/X VGND VGND VPWR VPWR _4163_/Y sky130_fd_sc_hd__o211ai_1
X_4094_ _3762_/A _3254_/X _3549_/X _3868_/A _3414_/X VGND VGND VPWR VPWR _4094_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__5229__A2 _5228_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3114_ _6047_/Q _6090_/Q _3116_/S VGND VGND VPWR VPWR _3115_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3045_ _5985_/B VGND VGND VPWR VPWR _3054_/S sky130_fd_sc_hd__buf_2
XANTENNA__4988__A1 _4984_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6188__CLK _6205_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4996_ _4996_/A VGND VGND VPWR VPWR _5102_/C sky130_fd_sc_hd__buf_2
XANTENNA__4344__A _4780_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5937__B1 _4765_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3947_ _4083_/C _3975_/D _3548_/X _3799_/X VGND VGND VPWR VPWR _3947_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4070__D1 _3230_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5952__A3 _5782_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3963__A2 _3249_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3878_ _3548_/X _3874_/X _3877_/Y _3241_/X VGND VGND VPWR VPWR _3878_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__5175__A _5175_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5617_ _5617_/A VGND VGND VPWR VPWR _6167_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5165__A1 _6121_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5548_ _5548_/A VGND VGND VPWR VPWR _6140_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3715__A2 _3477_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5903__A _5903_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5479_ _4803_/X _5090_/X _5445_/A _5451_/X _6119_/Q VGND VGND VPWR VPWR _5480_/A
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4676__B1 _4672_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5873__C1 _5872_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3423__A _3447_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4519__A _5203_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4140__A2 _3919_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_0_0_CLK clkbuf_4_1_0_CLK/A VGND VGND VPWR VPWR _6201_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_104_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4979__A1 _5431_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6156__D _6156_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4979__B2 input24/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2981__B _6098_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5928__B1 _5098_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4254__A _6136_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4600__B1 _5022_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5943__A3 _5529_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3954__A2 _3847_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input81_A memory_imem_request_put[7] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5156__A1 _5151_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4701__B _5191_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4903__A1 _4890_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3706__A2 _3705_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5813__A _5955_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5459__A2 _5433_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4429__A _4860_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5864__C1 _4824_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4131__A2 _3904_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3333__A _3437_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6066__D _6066_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3890__A1 _3357_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5919__B1 _5779_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4850_ _4850_/A _4974_/C VGND VGND VPWR VPWR _4850_/Y sky130_fd_sc_hd__nand2_1
X_3801_ _3614_/A _3447_/C _3571_/B VGND VGND VPWR VPWR _3801_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4781_ _5829_/C _4967_/A _4928_/A _4779_/Y _5006_/A VGND VGND VPWR VPWR _4781_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_33_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3732_ _4034_/B _3904_/B _3904_/C _3732_/D VGND VGND VPWR VPWR _3732_/X sky130_fd_sc_hd__or4_4
XANTENNA__3945__A2 _3573_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5147__A1 _5061_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3663_ _3663_/A _3711_/A _3663_/C _3938_/C VGND VGND VPWR VPWR _3663_/X sky130_fd_sc_hd__or4_4
XANTENNA__5698__A2 _5697_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3508__A _3508_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5402_ _5402_/A VGND VGND VPWR VPWR _6101_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3227__B _3606_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3594_ _3594_/A VGND VGND VPWR VPWR _3594_/X sky130_fd_sc_hd__clkbuf_4
X_5333_ _6053_/Q _6081_/Q _5339_/S VGND VGND VPWR VPWR _5334_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4370__A2 _5263_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4658__B1 _4777_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5264_ _5643_/A _5643_/B _6128_/Q VGND VGND VPWR VPWR _5264_/X sky130_fd_sc_hd__and3_1
XFILLER_87_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5195_ _4812_/X _5190_/X _4541_/X _5194_/Y VGND VGND VPWR VPWR _5195_/Y sky130_fd_sc_hd__o211ai_4
X_4215_ _4264_/C VGND VGND VPWR VPWR _4246_/B sky130_fd_sc_hd__buf_2
XANTENNA__5442__B _5468_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4122__A2 _6043_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5870__A2 _5866_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4146_ _4146_/A _4146_/B VGND VGND VPWR VPWR _4146_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5083__B1 _4746_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4077_ _3195_/B _3831_/X _4089_/B _3835_/X _3926_/X VGND VGND VPWR VPWR _4077_/Y
+ sky130_fd_sc_hd__o221ai_1
X_3028_ _6032_/Q _6164_/Q _3032_/S VGND VGND VPWR VPWR _3029_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4830__B1 _5182_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4074__A _4074_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5925__A3 _5845_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4979_ _5431_/A _4717_/X _4718_/X input24/X _4978_/X VGND VGND VPWR VPWR _4979_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_11_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3936__A2 _4074_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4802__A _5203_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5138__A1 _4403_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6203__CLK _6203_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3418__A _3588_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5689__A2 _5013_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4897__B1 _4945_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4361__A2 _5018_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5633__A _5633_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4113__A2 _3703_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5846__C1 _5093_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3153__A _3397_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5861__A2 _5706_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3872__A1 _4083_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5074__B1 _4946_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4821__B1 _4820_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5916__A3 _4890_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5377__A1 _6097_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5129__A1 _4984_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3328__A _3781_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4888__B1 _5761_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5543__A _5543_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3560__B1 _3628_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_7_0_CLK clkbuf_3_7_0_CLK/A VGND VGND VPWR VPWR clkbuf_3_7_0_CLK/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4104__A2 _3891_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5852__A2 _4534_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4000_ _3992_/A _3998_/X _3999_/X _3962_/A VGND VGND VPWR VPWR _4000_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3063__A _3096_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3998__A _3998_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3863__A1 _3161_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5065__B1 _5063_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3613__C_N _3612_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5951_ _4459_/X _4918_/A _5098_/X _5721_/A _4619_/X VGND VGND VPWR VPWR _5951_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_65_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4812__B1 _5078_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4902_ _4403_/X _4894_/X _4898_/Y _4901_/X VGND VGND VPWR VPWR _4902_/Y sky130_fd_sc_hd__o31ai_1
XANTENNA__5080__A3 _5009_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3510__B _3719_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5882_ _5879_/Y _5881_/Y _4765_/X VGND VGND VPWR VPWR _5882_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3002__S _3010_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4833_ _5899_/B _4843_/C _5118_/A _4675_/A VGND VGND VPWR VPWR _4833_/X sky130_fd_sc_hd__a31o_1
XFILLER_60_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5368__A1 _6143_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4040__A1 _4073_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4764_ _4875_/A VGND VGND VPWR VPWR _4765_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__4591__A2 _4437_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4040__B2 _3543_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4341__B _4341_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3715_ _3699_/X _3477_/X _3706_/X _3714_/X VGND VGND VPWR VPWR _3715_/X sky130_fd_sc_hd__a31o_1
XFILLER_107_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4695_ _4707_/D VGND VGND VPWR VPWR _4890_/A sky130_fd_sc_hd__buf_2
X_3646_ _3548_/X _4135_/A _3938_/C _3645_/Y _3546_/X VGND VGND VPWR VPWR _3646_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_20_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3577_ _3838_/A VGND VGND VPWR VPWR _3577_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5453__A _5453_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5316_ _5316_/A VGND VGND VPWR VPWR _6073_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5247_ _4347_/A _4369_/D _4843_/B _5118_/D VGND VGND VPWR VPWR _5247_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5828__C1 _5827_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5843__A2 _4971_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5178_ _4772_/A _4788_/B _5191_/A _5188_/B VGND VGND VPWR VPWR _5706_/C sky130_fd_sc_hd__o211ai_4
XANTENNA__3854__A1 _3701_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5599__S _5605_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5056__B1 _4771_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4129_ _3835_/X _3305_/A _3762_/A _3876_/X _3350_/A VGND VGND VPWR VPWR _4129_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__4219__D _4219_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3701__A _3701_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5071__A3 _4927_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3420__B _3838_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5359__A1 _6093_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5221__A2_N _5040_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4031__A1 _3685_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5628__A _5628_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3148__A _3446_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5236__A2_N _5233_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3790__B1 _4146_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4334__A2 _4244_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2987__A _2987_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3542__B1 _6019_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input44_A memory_dmem_request_put[70] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5834__A2 _5745_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4098__A1 _4105_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5295__B1 _5293_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3845__A1 _3844_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4707__A _4865_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3611__A _3611_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5302__S _5306_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5047__B1 _4241_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4270__A1 _4601_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4442__A _4442_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5538__A _5538_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4022__A1 _3666_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4573__A2 _4332_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3500_ _3500_/A VGND VGND VPWR VPWR _3911_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__5770__A1 _5676_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4480_ _5711_/A _4725_/A _4480_/C _4960_/A VGND VGND VPWR VPWR _4480_/X sky130_fd_sc_hd__and4_1
X_3431_ _3428_/X _3410_/A _3429_/X _3653_/B VGND VGND VPWR VPWR _3431_/Y sky130_fd_sc_hd__a211oi_1
XANTENNA__5522__A1 _6132_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4730__C1 _4923_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3362_ _3632_/A _3858_/A _3983_/B VGND VGND VPWR VPWR _3362_/Y sky130_fd_sc_hd__o21ai_4
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6150_ _6197_/CLK _6150_/D VGND VGND VPWR VPWR _6150_/Q sky130_fd_sc_hd__dfxtp_1
X_5101_ _5004_/A _5099_/X _5100_/X VGND VGND VPWR VPWR _5101_/Y sky130_fd_sc_hd__a21oi_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3293_ _3526_/A VGND VGND VPWR VPWR _3293_/X sky130_fd_sc_hd__buf_6
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ _6203_/CLK _6081_/D VGND VGND VPWR VPWR _6081_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5825__A2 _4316_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5032_ _4551_/A _5073_/A _4999_/A _4472_/X VGND VGND VPWR VPWR _5032_/Y sky130_fd_sc_hd__o211ai_4
XANTENNA__3836__A1 _4135_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5720__B _5720_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3836__B2 _3975_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5038__B1 _5220_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5934_ _4785_/X _5933_/X _5704_/X _5734_/X VGND VGND VPWR VPWR _5934_/Y sky130_fd_sc_hd__o211ai_1
X_5865_ _5863_/Y _5864_/X _5734_/A VGND VGND VPWR VPWR _5865_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_80_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4352__A _4832_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4816_ _4814_/X _4815_/X _4819_/A VGND VGND VPWR VPWR _4816_/X sky130_fd_sc_hd__o21a_1
X_5796_ _4858_/Y _4859_/X _5704_/X _5795_/Y VGND VGND VPWR VPWR _5796_/Y sky130_fd_sc_hd__a2bb2oi_2
XANTENNA__5210__B1 _4498_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4013__A1 _3536_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4747_ _4747_/A VGND VGND VPWR VPWR _5123_/C sky130_fd_sc_hd__buf_2
XFILLER_107_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4678_ _4421_/A _4699_/A _4643_/A VGND VGND VPWR VPWR _4924_/A sky130_fd_sc_hd__o21ai_4
X_3629_ _3687_/B _3687_/A VGND VGND VPWR VPWR _3663_/C sky130_fd_sc_hd__nand2_2
XANTENNA__5513__B2 _5503_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5513__A1 _5495_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5816__A2 _5814_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3827__A1 _5388_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3134__C _4002_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4527__A _4527_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4246__B _4246_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6164__D _6164_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5790__A2_N _5646_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5358__A _5358_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5752__B2 _5145_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5752__A1 _5743_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3358__A3 _3356_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5805__B _5805_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3606__A _3606_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5093__A _5093_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3818__A1 _3807_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5807__A2 _5806_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4437__A _4437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5540__B _5540_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6071__CLK _6074_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4491__A1 _4487_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3341__A _3468_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6074__D _6074_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4779__C1 _4369_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3980_ _3338_/Y _3978_/Y _3546_/A _3979_/X VGND VGND VPWR VPWR _3980_/X sky130_fd_sc_hd__o211a_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5128__A2_N _5040_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5991__A1 _6198_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5440__B1 _5439_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5268__A _5570_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4172__A _4205_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5650_ _6109_/Q _4511_/X _5676_/A _5649_/X VGND VGND VPWR VPWR _5651_/B sky130_fd_sc_hd__o211a_1
X_4601_ _4601_/A VGND VGND VPWR VPWR _4777_/A sky130_fd_sc_hd__buf_2
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5581_ _6151_/Q _6019_/Q _5583_/S VGND VGND VPWR VPWR _5582_/A sky130_fd_sc_hd__mux2_1
X_4532_ _4431_/X _4524_/X _4374_/X _4531_/X VGND VGND VPWR VPWR _4532_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__4951__C1 _4950_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4463_ _4649_/A _5744_/A _4815_/D VGND VGND VPWR VPWR _4918_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__5715__B _5715_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3414_ _4004_/B _3527_/C _3708_/A VGND VGND VPWR VPWR _3414_/X sky130_fd_sc_hd__and3_4
X_6202_ _6202_/CLK _6202_/D VGND VGND VPWR VPWR _6202_/Q sky130_fd_sc_hd__dfxtp_1
X_4394_ _4642_/A VGND VGND VPWR VPWR _4395_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_97_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3345_ _3345_/A VGND VGND VPWR VPWR _3711_/B sky130_fd_sc_hd__clkbuf_2
X_6133_ _6146_/CLK _6133_/D VGND VGND VPWR VPWR _6133_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__5259__B1 _5388_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3276_ _3657_/A VGND VGND VPWR VPWR _3674_/B sky130_fd_sc_hd__buf_4
XANTENNA__5731__A _5731_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3809__A1 _3766_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _6201_/CLK _6064_/D VGND VGND VPWR VPWR _6064_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5015_/A VGND VGND VPWR VPWR _5220_/C sky130_fd_sc_hd__buf_4
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4347__A _4347_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_85_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3251__A _3275_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3690__C1 _3685_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5026__A3 _5008_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5917_ _5123_/C _5123_/B _5179_/X _5916_/X VGND VGND VPWR VPWR _5917_/Y sky130_fd_sc_hd__a31oi_4
XFILLER_41_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4785__A2 _4472_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3993__B1 _3562_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5848_ _5843_/X _5844_/X _5845_/X _5847_/X _5769_/X VGND VGND VPWR VPWR _5848_/X
+ sky130_fd_sc_hd__a311o_1
X_5779_ _5078_/D _5745_/B _4843_/B VGND VGND VPWR VPWR _5779_/X sky130_fd_sc_hd__a21o_2
XANTENNA__5195__C1 _5194_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4810__A _5188_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3745__B1 _3271_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4232__D _4232_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3129__C _6062_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6094__CLK _6204_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6159__D _6159_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5998__D _6201_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5265__A3 _5262_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4257__A _4700_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5670__B1 _5669_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3799__C _4149_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3161__A _3161_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3681__C1 _3680_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5017__A3 _4852_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4776__A2 _4926_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3579__A3 _3562_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5088__A _5093_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3984__B1 _3701_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5186__C1 _5185_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3736__B1 _3281_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3336__A _3582_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3751__A3 _3635_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5489__B1 _6011_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4161__B1 _4160_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6069__D _6069_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5551__A _5551_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3130_ _3301_/A VGND VGND VPWR VPWR _3538_/A sky130_fd_sc_hd__buf_2
XFILLER_121_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5270__B input3/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5110__C1 _4829_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3267__A2 _3249_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4167__A _4405_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3071__A _3071_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3061_ _3061_/A VGND VGND VPWR VPWR _3061_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3672__C1 _3327_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5413__B1 _5398_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5964__A1 _5176_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3963_ _3867_/X _3249_/X _3773_/C _3468_/X VGND VGND VPWR VPWR _3963_/X sky130_fd_sc_hd__a31o_1
XFILLER_50_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3894_ _3178_/X _3183_/X _3218_/X _3893_/X VGND VGND VPWR VPWR _3894_/X sky130_fd_sc_hd__o211a_1
X_5702_ _6111_/Q _4721_/X _5701_/X VGND VGND VPWR VPWR _5702_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3010__S _3010_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5148__D _5148_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5177__C1 _5070_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5716__A1 _5076_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5633_ _5633_/A VGND VGND VPWR VPWR _6174_/D sky130_fd_sc_hd__clkbuf_1
X_5564_ _5256_/A _5968_/B _4990_/X _4987_/X _5482_/A VGND VGND VPWR VPWR _5565_/B
+ sky130_fd_sc_hd__o32a_1
XANTENNA__3942__B1_N _3806_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4630__A _4630_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5192__A2 _4405_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4515_ _4515_/A VGND VGND VPWR VPWR _4978_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3246__A _3468_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3742__A3 _3608_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5495_ _5715_/A VGND VGND VPWR VPWR _5495_/X sky130_fd_sc_hd__clkbuf_2
X_4446_ _4585_/A VGND VGND VPWR VPWR _4869_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4377_ _4854_/A VGND VGND VPWR VPWR _4673_/A sky130_fd_sc_hd__clkbuf_4
X_3328_ _3781_/A VGND VGND VPWR VPWR _4092_/A sky130_fd_sc_hd__buf_2
XANTENNA__5461__A _5461_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ _6123_/CLK _6116_/D VGND VGND VPWR VPWR _6116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ _3802_/A _3437_/A VGND VGND VPWR VPWR _3260_/A sky130_fd_sc_hd__and2_1
XFILLER_73_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5652__B1 _4823_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4455__A1 _4654_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6047_ _6205_/CLK _6047_/D VGND VGND VPWR VPWR _6047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5404__B1 _5403_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5707__A1 _4378_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5707__B2 _4680_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5168__C1 _5020_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4540__A _4835_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3981__A3 _3977_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3718__B1 _3482_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5183__A2 _4777_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3156__A _3603_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4391__B1 _4390_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2995__A _2995_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5891__B1 _5213_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4694__A1 _4692_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3497__A2 _3362_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5371__A _5371_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3603__B _3603_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4997__A2 _5102_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output113_A _3067_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4715__A _5646_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4749__A2 _5976_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5946__A1 _5693_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3957__B1 _3700_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3421__A2 _3934_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4002__C_N _4001_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3992__C _3992_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3709__B1 _4105_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5174__A2 _5169_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4921__A2 _4812_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4300_ _4354_/A VGND VGND VPWR VPWR _5008_/A sky130_fd_sc_hd__buf_2
XFILLER_5_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5280_ _5269_/Y _5272_/Y _5279_/Y VGND VGND VPWR VPWR _5285_/B sky130_fd_sc_hd__a21o_1
XFILLER_114_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4134__B1 _3286_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4231_ _4231_/A _4231_/B _4231_/C _4231_/D VGND VGND VPWR VPWR _4232_/D sky130_fd_sc_hd__and4_2
XANTENNA__5882__B1 _4765_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5281__A input4/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5712__C _5712_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4162_ _4158_/Y _4159_/X _4161_/Y _3517_/X _3580_/A VGND VGND VPWR VPWR _4162_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_95_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4093_ _3567_/X _3932_/Y _3992_/A _4092_/X VGND VGND VPWR VPWR _4093_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5229__A3 _4563_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5634__A0 _6175_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3113_ _3113_/A VGND VGND VPWR VPWR _3113_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3044_ _3044_/A VGND VGND VPWR VPWR _3044_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4988__A2 _5757_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5937__A1 _5652_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4995_ _4988_/X _4991_/X _4241_/X _4994_/X VGND VGND VPWR VPWR _4995_/X sky130_fd_sc_hd__a2bb2o_2
XANTENNA__4070__C1 _3648_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3948__B1 _3673_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3946_ _3428_/X _3895_/X _3720_/X _3945_/X VGND VGND VPWR VPWR _3946_/X sky130_fd_sc_hd__o31a_1
XFILLER_51_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3963__A3 _3773_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3877_ _3343_/X _3875_/X _3844_/X _3876_/X _3350_/X VGND VGND VPWR VPWR _3877_/Y
+ sky130_fd_sc_hd__o221ai_1
X_5616_ _6167_/Q _6035_/Q _5616_/S VGND VGND VPWR VPWR _5617_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5165__A2 _4511_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5547_ _5988_/A _5547_/B VGND VGND VPWR VPWR _5548_/A sky130_fd_sc_hd__or2_1
XANTENNA__3715__A3 _3706_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3181__B_N _3442_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5478_ _5444_/X _5046_/A _5445_/X _5540_/A _5477_/X VGND VGND VPWR VPWR _6118_/D
+ sky130_fd_sc_hd__a311o_1
X_4429_ _4860_/C _4462_/A _4769_/B VGND VGND VPWR VPWR _4955_/A sky130_fd_sc_hd__nand3_4
XANTENNA__5903__B _5903_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4125__B1 _3359_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5191__A _5191_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4676__A1 _5755_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4676__B2 _4673_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5873__B1 _5905_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3423__B _3870_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5625__A0 _6171_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6132__CLK _6205_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4979__A2 _4717_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4535__A _4543_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2981__C _6097_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5928__B2 _4967_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3939__B1 _3938_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6172__D _6172_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4600__A1 _4347_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5366__A _5366_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5156__A2 _5154_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4903__A2 _4892_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input74_A memory_imem_request_put[10] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4798__A2_N _6049_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5813__B _5813_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5459__A3 _5767_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5864__B1 _4890_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3614__A _3614_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4429__B _4462_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3875__C1 _3631_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5616__A0 _6167_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5077__D1 _4943_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3890__A2 _6033_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3627__C1 _3594_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4445__A _4815_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5919__A1 _5028_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4780_ _4780_/A VGND VGND VPWR VPWR _5006_/A sky130_fd_sc_hd__buf_2
X_3800_ _3799_/X _3522_/X _3464_/X VGND VGND VPWR VPWR _3800_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_33_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6082__D _6082_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3731_ _3956_/A _3873_/B _3966_/C _3731_/D VGND VGND VPWR VPWR _3731_/X sky130_fd_sc_hd__or4_1
XANTENNA__4052__C1 _3621_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3945__A3 _4089_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5276__A _5276_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5147__A2 _5062_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3662_ _3658_/X _3661_/Y _3376_/X VGND VGND VPWR VPWR _3662_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4180__A _4219_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3593_ _4073_/B _3659_/D _3614_/A _3593_/D VGND VGND VPWR VPWR _3593_/X sky130_fd_sc_hd__and4b_2
X_5401_ _5401_/A _5422_/B VGND VGND VPWR VPWR _5402_/A sky130_fd_sc_hd__and2_1
X_5332_ _5332_/A VGND VGND VPWR VPWR _6080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4107__B1 _3509_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5855__B1 _5853_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4658__B2 _4778_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3524__A _3583_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5263_ _5263_/A VGND VGND VPWR VPWR _5643_/A sky130_fd_sc_hd__buf_2
X_5194_ _4305_/Y _5192_/X _5193_/X VGND VGND VPWR VPWR _5194_/Y sky130_fd_sc_hd__o21bai_2
X_4214_ _4243_/A VGND VGND VPWR VPWR _5757_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__6155__CLK _6155_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4145_ _3460_/X _3762_/A _3910_/B _3875_/X _3868_/A VGND VGND VPWR VPWR _4146_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_95_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5083__A1 _5075_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4076_ _4073_/X _4075_/X _3479_/X _3838_/X VGND VGND VPWR VPWR _4076_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4830__A1 _4929_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4355__A _4729_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3027_ _3027_/A VGND VGND VPWR VPWR _3027_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3094__A0 _6053_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4074__B _4074_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4978_ _4978_/A VGND VGND VPWR VPWR _4978_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4594__B1 _4744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3929_ _3732_/X _3926_/X _3781_/X _3928_/Y _3376_/X VGND VGND VPWR VPWR _3929_/Y
+ sky130_fd_sc_hd__a311oi_4
XANTENNA__3936__A3 _3519_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5138__A2 _5102_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4346__B1 _4339_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4897__B2 _5096_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4897__A1 _4483_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3434__A _3904_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4113__A3 _4074_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5846__B1 _5163_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3153__B _3609_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5861__A3 _5032_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6167__D _6167_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3872__A2 _3460_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5074__A1 _4865_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4821__A1 _4369_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4265__A _4265_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5377__A2 _5368_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5096__A _5096_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6028__CLK _6155_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3609__A _3609_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5129__A2 _5757_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4888__B2 _5687_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4888__A1 _4488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6178__CLK _6207_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3344__A _3344_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3560__A1 _3548_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5543__B _5568_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5837__B1 _4345_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3201__A_N _3330_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6077__D _6077_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3998__B _4092_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3863__A2 _3857_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5065__A1 _5061_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5065__B2 _5064_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5950_ _6194_/Q _4799_/X _5941_/Y _5949_/X VGND VGND VPWR VPWR _6194_/D sky130_fd_sc_hd__o22a_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4175__A _4217_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4812__A1 _4843_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4901_ _4899_/X _4900_/X _4856_/A _4563_/A VGND VGND VPWR VPWR _4901_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3510__C _3983_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5881_ _5025_/Y _5880_/X _4930_/X _4305_/Y _5004_/A VGND VGND VPWR VPWR _5881_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4832_ _4832_/A VGND VGND VPWR VPWR _5118_/A sky130_fd_sc_hd__buf_4
XANTENNA__4025__C1 _3911_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5368__A2 _4211_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4763_ _4755_/X _5829_/B _4757_/X _4762_/Y VGND VGND VPWR VPWR _4763_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__4576__B1 _5029_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4040__A2 _4149_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4694_ _4692_/X _4693_/X _5179_/A _4290_/Y VGND VGND VPWR VPWR _4694_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3519__A _4092_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3714_ _3613_/B _3707_/X _3538_/A _3713_/Y VGND VGND VPWR VPWR _3714_/X sky130_fd_sc_hd__a211o_1
XFILLER_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3238__B _3557_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4341__C _4405_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5734__A _5734_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3645_ _3645_/A _3645_/B VGND VGND VPWR VPWR _3645_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3576_ _3934_/C _3576_/B VGND VGND VPWR VPWR _3576_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4628__A2_N _4190_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5315_ _6181_/Q _6073_/Q _5317_/S VGND VGND VPWR VPWR _5316_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5453__B _5468_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5246_ _5687_/A _4604_/X _5079_/B _5829_/C VGND VGND VPWR VPWR _5246_/Y sky130_fd_sc_hd__a31oi_1
XANTENNA__5828__B1 _5732_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3254__A _3847_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5843__A3 _4793_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5177_ _5061_/X _5062_/X _4668_/X _5176_/X _5070_/Y VGND VGND VPWR VPWR _5177_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_56_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3854__A2 _3241_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5056__A1 _4461_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4128_ _4128_/A _4128_/B VGND VGND VPWR VPWR _4128_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5056__B2 _5020_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4059_ _3832_/A _3583_/C _3362_/Y _3867_/A VGND VGND VPWR VPWR _4059_/X sky130_fd_sc_hd__o211a_1
XFILLER_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3420__C _3420_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6005__B1 _6004_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4016__C1 _4124_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4567__B1 _4580_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3429__A _3574_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4031__A2 _3962_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4319__B1 _4318_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4123__A1_N _3773_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3790__A1 _3607_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4334__A3 _4308_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3542__A1 _3507_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3542__B2 _3541_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3164__A _3876_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4098__A2 _3859_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5295__A1 _5291_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input37_A memory_dmem_request_put[63] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5834__A3 _5710_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3845__A2 _3687_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4707__B _4862_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3058__A0 _6189_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5047__B2 _5046_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3103__S _3105_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4270__A2 _4602_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5819__A _5819_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4007__C1 _3860_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4558__B1 _4252_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3339__A _3864_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4022__A2 _3194_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5770__A2 _5768_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5554__A _5554_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3430_ _3746_/B VGND VGND VPWR VPWR _3653_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_7_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5522__A2 _5504_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4730__B1 _5687_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3361_ _3254_/X _4135_/C _3208_/X VGND VGND VPWR VPWR _3361_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_112_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5100_ _5004_/D _4675_/X _5080_/X _4642_/X VGND VGND VPWR VPWR _5100_/X sky130_fd_sc_hd__a31o_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6080_ _6176_/CLK _6080_/D VGND VGND VPWR VPWR _6080_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3074__A _3096_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3292_ _3366_/A _3432_/B VGND VGND VPWR VPWR _3526_/A sky130_fd_sc_hd__or2_2
X_5031_ _5140_/C VGND VGND VPWR VPWR _5031_/X sky130_fd_sc_hd__clkbuf_4
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5825__A3 _5823_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3802__A _3802_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3836__A2 _3834_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5038__A1 _4952_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3013__S _3021_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5933_ _4360_/X _4740_/X _4771_/X _4957_/X VGND VGND VPWR VPWR _5933_/X sky130_fd_sc_hd__o211a_1
XFILLER_53_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5729__A _5811_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5864_ _4693_/X _5123_/C _4953_/X _4890_/C _4824_/X VGND VGND VPWR VPWR _5864_/X
+ sky130_fd_sc_hd__a311o_1
X_4815_ _4862_/A _4929_/A _4815_/C _4815_/D VGND VGND VPWR VPWR _4815_/X sky130_fd_sc_hd__and4_1
XANTENNA__3249__A _3603_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5795_ _4422_/X _4423_/X _5060_/X _5794_/Y VGND VGND VPWR VPWR _5795_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__5210__A1 _5011_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4013__A2 _3701_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4746_ _4746_/A _4746_/B VGND VGND VPWR VPWR _4746_/Y sky130_fd_sc_hd__nand2_1
XFILLER_107_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4677_ _5004_/A _4669_/Y _4676_/X VGND VGND VPWR VPWR _4677_/Y sky130_fd_sc_hd__a21oi_1
X_3628_ _3628_/A _3748_/B _3628_/C VGND VGND VPWR VPWR _3628_/X sky130_fd_sc_hd__or3_1
XANTENNA__5483__A1_N _5482_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5513__A2 _4720_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3559_ _3438_/X _3558_/X _3308_/X VGND VGND VPWR VPWR _3559_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5229_ _4894_/X _5228_/X _4563_/X _4685_/A VGND VGND VPWR VPWR _5229_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3827__A2 _6031_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3134__D _3822_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4527__B _4536_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4505__A2_N _4190_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4246__C _4246_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3460__B1 _3468_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4543__A _4543_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5639__A _5639_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5737__C1 _5018_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_CLK clkbuf_3_7_0_CLK/A VGND VGND VPWR VPWR clkbuf_3_6_0_CLK/X sky130_fd_sc_hd__clkbuf_2
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3159__A _3647_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6180__D _6180_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5752__A2 _5743_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5805__C _5805_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4712__B1 _4503_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4000__A1_N _3992_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5313__S _5317_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4718__A _4718_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output143_A _2999_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3818__A2 _3767_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4491__A2 _4488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4437__B _5048_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4228__C1 _4804_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4779__B1 _4369_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5440__A1 input17/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5440__B2 input9/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5991__A2 _5570_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5728__C1 _5727_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4600_ _4347_/A _5867_/C _4946_/A _5022_/A VGND VGND VPWR VPWR _4600_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3069__A _3069_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6090__D _6090_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4172__B _4205_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5580_ _5580_/A VGND VGND VPWR VPWR _6150_/D sky130_fd_sc_hd__clkbuf_1
X_4531_ _5878_/B _5687_/C _5107_/A VGND VGND VPWR VPWR _4531_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4951__B1 _4949_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4462_ _4462_/A VGND VGND VPWR VPWR _4649_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5715__C _5968_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5284__A _5284_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3413_ _3642_/A VGND VGND VPWR VPWR _3708_/A sky130_fd_sc_hd__clkbuf_2
X_6201_ _6201_/CLK _6201_/D VGND VGND VPWR VPWR _6201_/Q sky130_fd_sc_hd__dfxtp_1
X_4393_ _4685_/A VGND VGND VPWR VPWR _4393_/X sky130_fd_sc_hd__buf_4
XANTENNA__3008__S _3010_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3344_ _3344_/A _3432_/B VGND VGND VPWR VPWR _3345_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5259__A1 _5256_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6132_ _6205_/CLK _6132_/D VGND VGND VPWR VPWR _6132_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3275_ _3513_/A _3275_/B VGND VGND VPWR VPWR _3657_/A sky130_fd_sc_hd__and2_1
XANTENNA__5731__B _5731_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _6201_/CLK _6063_/D VGND VGND VPWR VPWR _6063_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3532__A _4065_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5014_ _4633_/S _4501_/X _5013_/X VGND VGND VPWR VPWR _5015_/A sky130_fd_sc_hd__a21oi_4
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3809__A2 _3808_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3690__B1 _3612_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5916_ _5140_/B _4840_/X _4890_/A _5976_/B VGND VGND VPWR VPWR _5916_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4363__A _4363_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4785__A3 _4864_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3993__A1 _3748_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5847_ _6102_/Q _4807_/A _5905_/A _5846_/X VGND VGND VPWR VPWR _5847_/X sky130_fd_sc_hd__o211a_1
X_5778_ _5776_/Y _4457_/X _5006_/X _5777_/X VGND VGND VPWR VPWR _5778_/X sky130_fd_sc_hd__a211o_2
XANTENNA__5195__B1 _4541_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4729_ _4895_/A _4729_/B _4926_/A VGND VGND VPWR VPWR _4923_/A sky130_fd_sc_hd__nand3_4
XANTENNA__3745__A1 _4089_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3707__A _3707_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5670__A1 _4652_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6175__D _6175_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3681__B1 _3645_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5958__C1 _5957_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4273__A _6135_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3984__A1 _3414_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5186__B1 _4950_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4933__B1 _4932_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3736__A1 _3735_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3617__A _3754_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3336__B _3437_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5489__A1 _5201_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4161__A1 _3868_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5110__B1 _4882_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4449__C1 _4448_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3060_ _6190_/Q _6066_/Q _3060_/S VGND VGND VPWR VPWR _3061_/A sky130_fd_sc_hd__mux2_2
XFILLER_95_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3267__A3 _3612_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6085__D _6085_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3672__B1 _3653_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5949__C1 _5948_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4183__A _4265_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5279__A _5285_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5413__B2 _6103_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5413__A1 input11/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5964__A2 _5179_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3962_ _3962_/A VGND VGND VPWR VPWR _3962_/X sky130_fd_sc_hd__buf_2
X_5701_ _5772_/A _5772_/B _5701_/C VGND VGND VPWR VPWR _5701_/X sky130_fd_sc_hd__and3_1
X_3893_ _4149_/A _3932_/B _3893_/C VGND VGND VPWR VPWR _3893_/X sky130_fd_sc_hd__or3_1
XFILLER_31_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5177__B1 _4668_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5716__A2 _4459_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5632_ _6174_/Q _6042_/Q _5638_/S VGND VGND VPWR VPWR _5633_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5563_ _5563_/A VGND VGND VPWR VPWR _6145_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5192__A3 _4865_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3527__A _3773_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4514_ _4976_/A VGND VGND VPWR VPWR _5805_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__3246__B _3780_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5494_ _5494_/A VGND VGND VPWR VPWR _6123_/D sky130_fd_sc_hd__clkbuf_1
X_4445_ _4815_/D VGND VGND VPWR VPWR _5079_/C sky130_fd_sc_hd__clkbuf_2
X_4376_ _4860_/A _4860_/B VGND VGND VPWR VPWR _4854_/A sky130_fd_sc_hd__nand2_4
XANTENNA__4358__A _4358_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_85_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3327_ _3571_/A VGND VGND VPWR VPWR _3327_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_58_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6115_ _6123_/CLK _6115_/D VGND VGND VPWR VPWR _6115_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3262__A _3657_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5101__B1 _5100_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _3344_/A VGND VGND VPWR VPWR _3802_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5652__A1 _5026_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4455__A2 _4363_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6046_ _6205_/CLK _6046_/D VGND VGND VPWR VPWR _6046_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3189_ _3344_/A VGND VGND VPWR VPWR _3781_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5404__A1 _4232_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4612__C1 _4619_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5707__A2 _5079_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5168__B1 _4927_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_3_7_0_CLK_A clkbuf_3_7_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3718__B2 _3510_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3718__A1 _3410_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4915__B1 _4905_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5742__A2_N _4378_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5183__A3 _4778_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3437__A _3437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4391__A1 _5715_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6061__CLK _6204_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5891__A1 _5211_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4694__A2 _4693_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3497__A3 _3305_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3351__C1 _3350_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5371__B _6097_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4268__A _4268_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3172__A _4044_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3603__C _3612_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4603__C1 _4462_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4749__A3 _5123_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5946__A2 _5943_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output106_A _3117_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3957__A1 _3612_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3421__A3 _3414_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5159__B1 _5132_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3709__A1 _4074_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4906__B1 input15/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3347__A _3499_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4921__A3 _4917_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5562__A _5562_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4134__A1 _4127_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4230_ _4230_/A _4230_/B _4230_/C VGND VGND VPWR VPWR _4232_/B sky130_fd_sc_hd__and3_2
XFILLER_4_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5331__A0 _6188_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5882__A1 _5879_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4161_ _3868_/X _3653_/X _3910_/X _4160_/Y VGND VGND VPWR VPWR _4161_/Y sky130_fd_sc_hd__o31ai_1
XANTENNA__5712__D _5712_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4178__A _4218_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3082__A _3082_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4092_ _4092_/A _4092_/B _4092_/C _4092_/D VGND VGND VPWR VPWR _4092_/X sky130_fd_sc_hd__or4_1
XFILLER_67_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3112_ _6046_/Q _6089_/Q _3116_/S VGND VGND VPWR VPWR _3113_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5634__A1 _6043_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3043_ _6039_/Q _6171_/Q _3043_/S VGND VGND VPWR VPWR _3044_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4988__A3 _5757_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5937__A2 _5936_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3021__S _3021_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4994_ input6/X _4994_/B _4200_/B VGND VGND VPWR VPWR _4994_/X sky130_fd_sc_hd__or3b_2
XFILLER_23_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4070__B1 _3962_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3945_ _3666_/A _3573_/X _4089_/B _3319_/X VGND VGND VPWR VPWR _3945_/X sky130_fd_sc_hd__o31a_1
XANTENNA__3948__A1 _3403_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6084__CLK _6202_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3876_ _3876_/A _3876_/B VGND VGND VPWR VPWR _3876_/X sky130_fd_sc_hd__or2_4
X_5615_ _5615_/A VGND VGND VPWR VPWR _6166_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3257__A _3462_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5546_ _5093_/X _5715_/B _4802_/X _6140_/Q _5482_/X VGND VGND VPWR VPWR _5547_/B
+ sky130_fd_sc_hd__o32a_1
X_5477_ _6118_/Q _4239_/X _5093_/X _4802_/X VGND VGND VPWR VPWR _5477_/X sky130_fd_sc_hd__o22a_1
X_4428_ _4705_/A VGND VGND VPWR VPWR _4769_/B sky130_fd_sc_hd__buf_2
XANTENNA__5903__C _5903_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5858__D1 _5857_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4125__A1 _3178_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4125__B2 _3904_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5322__A0 _6184_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4676__A2 _4671_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5873__A1 _6103_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4359_ _4878_/C VGND VGND VPWR VPWR _4668_/B sky130_fd_sc_hd__buf_2
XFILLER_59_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5625__A1 _6039_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6029_ _6155_/CLK _6029_/D VGND VGND VPWR VPWR _6029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3720__A _3720_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_67_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5389__B1 _4859_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3939__A1 _4105_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4551__A _4551_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4600__A2 _5867_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5647__A _5822_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5010__C1 _5711_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3167__A _3437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5561__B1 _5499_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input67_A memory_dmem_request_put[93] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5813__C _5813_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5313__A0 _6196_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5382__A _6099_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5864__A1 _4693_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3324__C1 _4146_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4429__C _4769_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3875__B1 _3462_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5077__C1 _4824_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4726__A _4726_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5616__A1 _6035_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3630__A _3663_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3627__B1 _3271_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5919__A2 _5880_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4052__B1 _3934_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4461__A _4461_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3730_ _3437_/A _3446_/B _3657_/B VGND VGND VPWR VPWR _3731_/D sky130_fd_sc_hd__o21ai_4
XFILLER_13_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3661_ _3659_/X _3660_/X _3429_/X VGND VGND VPWR VPWR _3661_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__4180__B _4219_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3592_ _3592_/A VGND VGND VPWR VPWR _3593_/D sky130_fd_sc_hd__buf_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5552__B1 _6142_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5400_ input5/X VGND VGND VPWR VPWR _5422_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5331_ _6188_/Q _6080_/Q _5339_/S VGND VGND VPWR VPWR _5332_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4107__A1 _3537_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4107__B2 _4040_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5292__A _6204_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5304__A0 _6192_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5855__A1 _5852_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5262_ _4716_/X _4513_/X input36/X _5045_/A _5261_/X VGND VGND VPWR VPWR _5262_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_114_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5855__B2 _5854_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5193_ _5118_/B _5711_/A _4697_/A _4869_/A VGND VGND VPWR VPWR _5193_/X sky130_fd_sc_hd__a31o_1
X_4213_ _4307_/A VGND VGND VPWR VPWR _4243_/A sky130_fd_sc_hd__clkbuf_2
X_4144_ _3910_/C _3299_/A _3369_/X _3603_/A _3537_/A VGND VGND VPWR VPWR _4144_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4636__A _4860_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5083__A2 _5077_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4075_ _3834_/X _3428_/X _3938_/C _4074_/X VGND VGND VPWR VPWR _4075_/X sky130_fd_sc_hd__a211o_1
XFILLER_36_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3026_ _6031_/Q _6163_/Q _3032_/S VGND VGND VPWR VPWR _3027_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3094__A1 _6081_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4830__A2 _4883_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4074__C _4074_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4594__A1 _4668_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4043__B1 _3648_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4977_ _5772_/B VGND VGND VPWR VPWR _4977_/X sky130_fd_sc_hd__clkbuf_2
X_3928_ _4124_/A _3895_/X _3847_/X _3701_/A VGND VGND VPWR VPWR _3928_/Y sky130_fd_sc_hd__a211oi_2
XANTENNA__5138__A3 _4574_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3859_ _3859_/A VGND VGND VPWR VPWR _4124_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_50_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5159__A1_N _4799_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4346__B2 _4345_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4346__A1 _4306_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4897__A2 _4485_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5529_ _5529_/A VGND VGND VPWR VPWR _5529_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5846__A1 input10/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3857__B1 _3447_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5861__A4 _5068_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4546__A _4854_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5074__A2 _4865_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4806__C1 _4805_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4265__B _4283_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4983__A1_N _4974_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4821__A2 _4480_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6183__D _6183_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5231__C1 _4675_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4281__A _4738_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3609__B _3609_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3793__C1 _3674_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5129__A3 _5757_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4888__A2 _4887_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5837__A1 _5834_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3560__A2 _3554_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6001__A _6207_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3344__B _3432_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3848__B1 _3847_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3998__C _3998_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3360__A _3711_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4456__A _5667_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5065__A2 _5062_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4175__B _4217_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4812__A2 _4843_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4900_ _4297_/X _4536_/X _4873_/A _4580_/A VGND VGND VPWR VPWR _4900_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3510__D _4092_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5880_ _5880_/A VGND VGND VPWR VPWR _5880_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6093__D _6093_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4831_ _5745_/C _4843_/B _4829_/Y _5880_/A VGND VGND VPWR VPWR _4831_/X sky130_fd_sc_hd__o211a_1
XFILLER_33_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4025__B1 _3205_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5368__A3 _5367_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5287__A input5/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4762_ _5152_/B _4956_/D _4923_/A _4761_/X VGND VGND VPWR VPWR _4762_/Y sky130_fd_sc_hd__a31oi_4
XANTENNA__4576__A1 _4480_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4191__A input8/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5773__B1 _5772_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4693_ _5188_/C VGND VGND VPWR VPWR _4693_/X sky130_fd_sc_hd__buf_2
XANTENNA__4040__A3 _3998_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3713_ _3621_/X _3709_/X _3712_/X VGND VGND VPWR VPWR _3713_/Y sky130_fd_sc_hd__a21oi_1
X_3644_ _3633_/A _3711_/B _3499_/A _3543_/B VGND VGND VPWR VPWR _3645_/B sky130_fd_sc_hd__o22a_2
XANTENNA__3238__C _3549_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4341__D _4405_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6122__CLK _6147_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3575_ _3910_/B _3519_/X _3573_/X _3520_/X _3574_/X VGND VGND VPWR VPWR _3576_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5314_ _5314_/A VGND VGND VPWR VPWR _6072_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5828__A1 _4360_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5245_ _4541_/X _4464_/X _5243_/X _5244_/X VGND VGND VPWR VPWR _5245_/X sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_4_6_0_CLK_A clkbuf_4_7_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3839__B1 _3838_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5176_ _5944_/D VGND VGND VPWR VPWR _5176_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_56_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3854__A3 _3848_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5056__A2 _4576_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3270__A _4074_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4127_ _3636_/X _4123_/X _4124_/X _3685_/X _4126_/Y VGND VGND VPWR VPWR _4127_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_83_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4058_ _3338_/Y _3564_/X _3546_/X VGND VGND VPWR VPWR _4058_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_45_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3009_ _3009_/A VGND VGND VPWR VPWR _3009_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__6005__A1 _6203_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4016__B1 _3194_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4571__A_N _5715_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4567__A1 _4929_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5764__B1 _5228_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4031__A3 _3414_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4319__A1 _4482_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3790__A2 _3733_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5516__B1 _5504_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4334__A4 _4245_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3542__A2 _3540_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6178__D _6178_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4098__A3 _3704_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5295__A2 _5292_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3845__A3 _3534_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4276__A _4769_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3180__A _3226_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4707__C _4707_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4255__B1 _4254_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3058__A1 _6065_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4007__B1 _3660_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5204__C1 _5260_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4558__A1 _4542_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6145__CLK _6145_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4022__A3 _3767_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3944__A2_N _3943_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5507__B1 _6127_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output98_A _3102_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4730__A1 _5078_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3360_ _3711_/B VGND VGND VPWR VPWR _4135_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_112_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6088__D _6088_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3291_ _3387_/B VGND VGND VPWR VPWR _3432_/B sky130_fd_sc_hd__clkbuf_2
X_5030_ _4761_/X _5028_/X _4927_/A _4726_/A _5029_/X VGND VGND VPWR VPWR _5030_/X
+ sky130_fd_sc_hd__o221a_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3802__B _3802_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3836__A3 _3835_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4186__A _4186_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5038__A2 _5012_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5932_ _5925_/Y _5931_/Y _4190_/X _6193_/Q VGND VGND VPWR VPWR _6193_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_80_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5994__B1 _5986_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5863_ _4726_/A _5070_/Y _4742_/X _4387_/X VGND VGND VPWR VPWR _5863_/Y sky130_fd_sc_hd__a31oi_1
XANTENNA__5729__B _5729_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4814_ _4864_/C _4643_/A _4864_/A _4780_/A VGND VGND VPWR VPWR _4814_/X sky130_fd_sc_hd__a31o_1
X_5794_ _4786_/X _5062_/A _5721_/B _5793_/Y VGND VGND VPWR VPWR _5794_/Y sky130_fd_sc_hd__a2bb2oi_4
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4745_ _5712_/C _4737_/Y _4743_/Y _4744_/X VGND VGND VPWR VPWR _4746_/B sky130_fd_sc_hd__o211ai_1
XANTENNA__5210__A2 _5209_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4013__A3 _3501_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5745__A _5745_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4676_ _5755_/B _4671_/X _4672_/X _4673_/Y _4675_/X VGND VGND VPWR VPWR _4676_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3265__A _3574_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3627_ _3626_/X _3342_/X _3271_/A _3594_/X VGND VGND VPWR VPWR _3628_/C sky130_fd_sc_hd__o211a_1
XANTENNA__5513__A3 _5498_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5438__B_N _4227_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3558_ _3968_/A _4149_/B _3660_/B VGND VGND VPWR VPWR _3558_/X sky130_fd_sc_hd__or3_2
XFILLER_1_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3489_ _3648_/A _4074_/B _4135_/C VGND VGND VPWR VPWR _3489_/X sky130_fd_sc_hd__or3_2
XANTENNA__5480__A _5480_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5228_ _5228_/A VGND VGND VPWR VPWR _5228_/X sky130_fd_sc_hd__buf_4
XFILLER_103_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5159_ _4799_/X _6056_/Q _5132_/X _5158_/Y VGND VGND VPWR VPWR _6056_/D sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__6018__CLK _6155_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4527__C _4527_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4237__A0 _4229_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6168__CLK _6203_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3460__A1 _3663_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5737__B1 _4864_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3175__A _3440_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4712__A1 _4685_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5390__A _5432_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3818__A3 _3817_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output136_A _3047_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4491__A3 _4843_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3114__S _3116_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4228__B1 _4718_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4734__A _4734_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4779__A1 _4777_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5440__A2 _5437_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3987__C1 _3986_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5728__B1 _5676_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4172__C _4205_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5565__A _5988_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4530_ _4661_/A VGND VGND VPWR VPWR _5107_/A sky130_fd_sc_hd__buf_4
XANTENNA__4951__A1 _4938_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4461_ _4461_/A VGND VGND VPWR VPWR _4461_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_7_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_1_1_0_CLK_A clkbuf_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3412_ _3582_/C _3446_/B VGND VGND VPWR VPWR _3642_/A sky130_fd_sc_hd__nor2_2
X_6200_ _6201_/CLK _6200_/D VGND VGND VPWR VPWR _6200_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3085__A _3096_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5900__B1 _5235_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4392_ _4767_/A VGND VGND VPWR VPWR _4685_/A sky130_fd_sc_hd__clkbuf_2
X_6131_ _6145_/CLK _6131_/D VGND VGND VPWR VPWR _6131_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5392__A_N input7/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3343_ _3343_/A VGND VGND VPWR VPWR _3343_/X sky130_fd_sc_hd__buf_2
XANTENNA__4909__A _5757_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5259__A2 _2986_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3274_ _4152_/C VGND VGND VPWR VPWR _3815_/C sky130_fd_sc_hd__clkbuf_4
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6201_/CLK _6062_/D VGND VGND VPWR VPWR _6062_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5013_ _4990_/X _6146_/Q _5013_/S VGND VGND VPWR VPWR _5013_/X sky130_fd_sc_hd__mux2_8
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3024__S _3032_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3690__A1 _4124_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4644__A _4827_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5967__B1 _5958_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5915_ _5910_/X _5911_/X _5237_/X _5914_/Y VGND VGND VPWR VPWR _5915_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_53_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5719__B1 _5955_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3993__A2 _3988_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4785__A4 _4865_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5846_ input10/X _5395_/A _5163_/A _5093_/A VGND VGND VPWR VPWR _5846_/X sky130_fd_sc_hd__a211o_1
XFILLER_42_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5777_ _4953_/X _5761_/C _4574_/A _5903_/A _4572_/X VGND VGND VPWR VPWR _5777_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5195__A1 _4812_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2989_ _5294_/A VGND VGND VPWR VPWR _3060_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_21_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5475__A _5475_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4728_ _4728_/A VGND VGND VPWR VPWR _4926_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3745__A2 _3499_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4659_ _4728_/A VGND VGND VPWR VPWR _5188_/D sky130_fd_sc_hd__buf_4
XFILLER_1_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4819__A _4819_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3442__B _3442_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5655__C1 _5145_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_3_0_CLK_A clkbuf_3_3_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5670__A2 _5666_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3681__A1 _3830_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_83_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5958__B1 _5955_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6191__D _6191_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3984__A2 _3983_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5186__A1 _5177_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4933__A1 _4922_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4933__B2 _4563_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3736__A2 _3645_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3197__B1 _3173_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3602__B1_N _3330_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_4_14_0_CLK_A clkbuf_3_7_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5489__A2 _5202_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5894__C1 _5893_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4729__A _4895_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3633__A _3633_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4161__A2 _3653_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5324__S _5328_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5110__A1 _4761_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4449__B1 _4431_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3267__A4 _3998_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3121__A0 _6049_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3672__A1 _3223_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4464__A _5903_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5949__B1 _5822_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4183__B _4265_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3961_ _3508_/X _3951_/X _3960_/Y VGND VGND VPWR VPWR _3961_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5279__B _5279_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5413__A2 _5412_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5964__A3 _5025_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5700_ _6182_/Q _5646_/X _5679_/Y _5699_/Y VGND VGND VPWR VPWR _6182_/D sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__3387__A_N _3311_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3892_ _3829_/X _3720_/X _3512_/X _3464_/X _3882_/X VGND VGND VPWR VPWR _3892_/Y
+ sky130_fd_sc_hd__a311oi_1
XFILLER_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5177__B2 _5176_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5177__A1 _5061_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5716__A3 _5192_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5631_ _5631_/A VGND VGND VPWR VPWR _6173_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5562_ _5562_/A _5568_/B VGND VGND VPWR VPWR _5563_/A sky130_fd_sc_hd__and2_1
XANTENNA__3527__B _3588_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4513_ _4513_/A VGND VGND VPWR VPWR _4513_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_105_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3019__S _3021_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5493_ _5493_/A _5501_/B VGND VGND VPWR VPWR _5494_/A sky130_fd_sc_hd__and2_1
X_4444_ _4549_/A _4884_/A VGND VGND VPWR VPWR _5903_/B sky130_fd_sc_hd__nand2_4
XANTENNA__4639__A _4929_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4375_ _4811_/A VGND VGND VPWR VPWR _4673_/B sky130_fd_sc_hd__buf_4
XANTENNA__3896__D1 _3537_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3543__A _3847_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3326_ _3528_/A VGND VGND VPWR VPWR _3571_/A sky130_fd_sc_hd__clkbuf_2
X_6114_ _6123_/CLK _6114_/D VGND VGND VPWR VPWR _6114_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5101__A1 _5004_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_5_0_CLK clkbuf_3_5_0_CLK/A VGND VGND VPWR VPWR clkbuf_3_5_0_CLK/X sky130_fd_sc_hd__clkbuf_2
X_6045_ _6045_/CLK _6045_/D VGND VGND VPWR VPWR _6045_/Q sky130_fd_sc_hd__dfxtp_1
X_3257_ _3462_/B VGND VGND VPWR VPWR _3831_/A sky130_fd_sc_hd__buf_4
XFILLER_86_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5652__A2 _5680_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3112__A0 _6046_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3188_ _3233_/A VGND VGND VPWR VPWR _3344_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4374__A _5240_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5404__A2 _4859_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4612__B1 _4536_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5829_ _5829_/A _5829_/B _5829_/C VGND VGND VPWR VPWR _5829_/X sky130_fd_sc_hd__and3_1
XANTENNA__5168__A1 _5167_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5168__B2 _4838_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6206__CLK _6207_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3718__A2 _3215_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4915__B2 _4914_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4915__A1 _6051_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3437__B _3437_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4391__A2 _4211_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4549__A _4549_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5891__A2 _5745_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3351__B1 _3410_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3453__A _4103_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4268__B _4268_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3172__B _3282_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6186__D _6186_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3603__D _3603_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3103__A0 _6057_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4851__B1 _4809_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input12_A memory_dmem_request_put[38] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4603__B1 _4728_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4749__A4 _5755_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5800__C1 _4255_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3957__A2 _4035_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5159__B2 _5158_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3709__A2 _3157_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3628__A _3628_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4906__A1 _5438_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4119__C1 _4118_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4035__A_N _3350_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3590__B1 _4128_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4459__A _4459_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4134__A2 _4133_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5562__B _5568_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5331__A1 _6080_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5882__A2 _5881_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4160_ _3815_/C _3673_/B _3482_/X _3510_/X _3717_/X VGND VGND VPWR VPWR _4160_/Y
+ sky130_fd_sc_hd__o221ai_1
XANTENNA__5249__A2_N _5246_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6096__D _6096_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4178__B _4218_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3111_ _3111_/A VGND VGND VPWR VPWR _3111_/X sky130_fd_sc_hd__clkbuf_1
X_4091_ _3194_/X _3834_/X _3293_/X _3975_/D _3308_/X VGND VGND VPWR VPWR _4091_/Y
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__5095__B1 _5094_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3042_ _3042_/A VGND VGND VPWR VPWR _3042_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4842__B1 _4732_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4993_ input25/X _4978_/A _4992_/X VGND VGND VPWR VPWR _4994_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__4070__A1 _3967_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3948__A2 _3519_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3944_ _3866_/X _3943_/X _5388_/B _6035_/Q VGND VGND VPWR VPWR _6035_/D sky130_fd_sc_hd__a2bb2o_1
X_3875_ _3711_/A _3588_/C _3462_/B _3631_/A VGND VGND VPWR VPWR _3875_/X sky130_fd_sc_hd__o211a_2
XANTENNA__5817__A2_N _4715_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3538__A _3538_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5614_ _6166_/Q _6034_/Q _5616_/S VGND VGND VPWR VPWR _5615_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5545_ _5545_/A VGND VGND VPWR VPWR _5988_/A sky130_fd_sc_hd__buf_4
X_5476_ _5476_/A VGND VGND VPWR VPWR _6117_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4369__A _4369_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4427_ _4313_/A _4293_/Y _4261_/Y _4209_/A VGND VGND VPWR VPWR _4705_/A sky130_fd_sc_hd__o2bb2ai_2
XANTENNA__5858__C1 _5175_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4125__A2 _3767_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5322__A1 _6076_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3273__A _3437_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5903__D _5903_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5873__A2 _5805_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4358_ _4358_/A VGND VGND VPWR VPWR _4878_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_86_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4088__B _4088_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input4_A EN_memory_imem_response_get VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4289_ _4578_/A VGND VGND VPWR VPWR _4725_/A sky130_fd_sc_hd__buf_2
X_3309_ _3956_/A VGND VGND VPWR VPWR _3614_/A sky130_fd_sc_hd__clkbuf_2
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5086__B1 _5047_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6028_ _6155_/CLK _6028_/D VGND VGND VPWR VPWR _6028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4833__B1 _4675_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5389__A1 _4246_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4832__A _4832_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3939__A2 _3271_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4551__B _4692_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4600__A3 _4946_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5010__B1 _4353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5561__A1 _5968_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5561__B2 _6145_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4279__A _4379_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5313__A1 _6072_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5382__B _5382_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5864__A2 _5123_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3183__A _4004_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3324__B1 _3320_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3875__A1 _3711_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5077__B1 _4823_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3911__A _3911_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3627__A1 _3626_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_2_0_0_CLK_A clkbuf_2_1_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4824__B1 _4649_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4726__B _5148_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4742__A _4742_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4052__A1 _3919_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3660_ _3841_/A _3660_/B _4092_/D _4152_/C VGND VGND VPWR VPWR _3660_/X sky130_fd_sc_hd__or4_1
XANTENNA__5001__B1 _4742_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3591_ _3591_/A VGND VGND VPWR VPWR _3659_/D sky130_fd_sc_hd__buf_2
XANTENNA__5552__A1 _5256_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5552__B2 _5482_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5330_ _5352_/A VGND VGND VPWR VPWR _5339_/S sky130_fd_sc_hd__buf_2
XANTENNA__5573__A _5629_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4107__A2 _4106_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5261_ input12/X _4717_/X _4718_/X input20/X _4804_/X VGND VGND VPWR VPWR _5261_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5304__A1 _6068_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5855__A2 _5721_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4212_ _4282_/A VGND VGND VPWR VPWR _4307_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3093__A _3093_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4189__A _4189_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5192_ _4404_/X _4405_/X _4865_/A _5899_/A VGND VGND VPWR VPWR _5192_/X sky130_fd_sc_hd__o31a_4
XFILLER_110_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4917__A _4917_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4143_ _4143_/A _4143_/B _3645_/A VGND VGND VPWR VPWR _4143_/X sky130_fd_sc_hd__or3b_1
XFILLER_68_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4074_ _4074_/A _4074_/B _4074_/C VGND VGND VPWR VPWR _4074_/X sky130_fd_sc_hd__and3_1
XANTENNA__3821__A _4103_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6051__CLK _6205_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3025_ _3025_/A VGND VGND VPWR VPWR _3025_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3032__S _3032_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4652__A _4652_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4043__A1 _3967_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_2_0_CLK_A clkbuf_4_3_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4200__A_N input6/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4976_ _4976_/A VGND VGND VPWR VPWR _5772_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__4594__A2 _5000_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3927_ _4048_/B VGND VGND VPWR VPWR _4124_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3268__A _3268_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3858_ _3858_/A _3876_/B VGND VGND VPWR VPWR _3859_/A sky130_fd_sc_hd__nor2_2
XANTENNA__4346__A2 _4316_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3789_ _5388_/B _6027_/Q _3788_/X VGND VGND VPWR VPWR _6027_/D sky130_fd_sc_hd__a21o_1
X_5528_ _5528_/A _5528_/B VGND VGND VPWR VPWR _6134_/D sky130_fd_sc_hd__nand2_1
XANTENNA__3554__B1 _3910_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5459_ _4977_/X _5433_/A _5767_/C _5451_/X _6113_/Q VGND VGND VPWR VPWR _5460_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_59_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3857__A1 _3666_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5846__A2 _5395_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4827__A _4827_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_86_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3731__A _3956_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5059__B1 _4568_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4806__B1 _4803_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4265__C _4265_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6008__C1 _4715_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3490__C1 _3489_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4562__A _5903_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5231__B1 _5080_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3178__A _3780_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3793__B1 _3767_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6001__B _6203_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5298__A0 _6189_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5837__A2 _5836_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3848__A1 _3343_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6074__CLK _6074_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3641__A _4149_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3998__D _3998_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4456__B _5029_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5470__B1 _5439_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4830_ _4929_/B _4883_/A _5182_/A VGND VGND VPWR VPWR _5880_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__4472__A _4566_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5568__A _5568_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4025__A1 _3895_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4761_ _4946_/A VGND VGND VPWR VPWR _4761_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__4576__A2 _4668_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5773__A1 _6114_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4692_ _4692_/A VGND VGND VPWR VPWR _4692_/X sky130_fd_sc_hd__clkbuf_4
X_3712_ _3710_/X _3992_/A _3711_/X _3491_/A VGND VGND VPWR VPWR _3712_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3784__B1 _3695_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3643_ _3643_/A VGND VGND VPWR VPWR _3645_/A sky130_fd_sc_hd__buf_2
XANTENNA__3238__D _3847_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3816__A _3816_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3574_ _3574_/A VGND VGND VPWR VPWR _3574_/X sky130_fd_sc_hd__buf_2
X_5313_ _6196_/Q _6072_/Q _5317_/S VGND VGND VPWR VPWR _5314_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5289__B1 _5288_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5828__A2 _5826_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5244_ _4563_/A _4673_/Y _5878_/A _4692_/X _5228_/A VGND VGND VPWR VPWR _5244_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_88_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3839__A1 _3536_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4647__A _5022_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5175_ _5175_/A VGND VGND VPWR VPWR _5175_/X sky130_fd_sc_hd__buf_4
XANTENNA__3551__A _3551_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4126_ _4126_/A _4126_/B VGND VGND VPWR VPWR _4126_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4057_ _4047_/X _3787_/X _4056_/Y _6040_/Q _3822_/X VGND VGND VPWR VPWR _6040_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_24_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3008_ _6023_/Q _6155_/Q _3010_/S VGND VGND VPWR VPWR _3009_/A sky130_fd_sc_hd__mux2_2
XANTENNA__4382__A _4700_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6005__A2 _5293_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5213__B1 _4862_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4016__A1 _3343_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4016__B2 _3533_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4567__A2 _5744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4959_ _5020_/A VGND VGND VPWR VPWR _4959_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5764__A1 _5722_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3775__B1 _3774_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4319__A2 _4234_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5516__A1 _4806_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3542__A3 _3453_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6097__CLK _6207_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3461__A _3461_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4274__A2_N _4272_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3845__A4 _3293_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4707__D _4707_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4255__A1 _4268_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6194__D _6194_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5452__B1 _5451_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4292__A _4738_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5388__A _5388_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4007__A1 _4083_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4007__B2 _3876_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5204__B1 _5968_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4558__A2 _4557_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3766__B1 _3765_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5507__A1 _5495_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3636__A _4128_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5507__B2 _5499_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4730__A2 _4488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ _4103_/C VGND VGND VPWR VPWR _3290_/X sky130_fd_sc_hd__buf_2
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5570__B _6199_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3371__A _3437_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4467__A _4875_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5691__B1 _5684_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3802__C _3895_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4186__B _6178_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5931_ _5237_/X _5930_/X _5955_/A VGND VGND VPWR VPWR _5931_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_19_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5994__A1 _5998_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5862_ _5179_/X _5859_/X _5860_/X _5861_/Y VGND VGND VPWR VPWR _5862_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_33_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5793_ _4296_/X _5078_/D _4673_/A _5118_/A VGND VGND VPWR VPWR _5793_/Y sky130_fd_sc_hd__o211ai_2
X_4813_ _4290_/Y _4617_/Y _4924_/A VGND VGND VPWR VPWR _4813_/X sky130_fd_sc_hd__a21o_1
X_4744_ _4744_/A VGND VGND VPWR VPWR _4744_/X sky130_fd_sc_hd__buf_4
XANTENNA__4930__A _5098_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5745__B _5745_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4675_ _4675_/A VGND VGND VPWR VPWR _4675_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3546__A _3546_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5726__A1_N _6183_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3626_ _3841_/B VGND VGND VPWR VPWR _3626_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_115_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3557_ _3557_/A VGND VGND VPWR VPWR _4149_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_115_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5761__A _5761_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3488_ _4044_/A VGND VGND VPWR VPWR _3488_/X sky130_fd_sc_hd__buf_2
XFILLER_0_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5480__B _5501_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5227_ _5222_/X _4630_/A _5225_/X _5226_/Y VGND VGND VPWR VPWR _5227_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4377__A _4854_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5682__B1 _5140_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3281__A _3281_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5158_ _5141_/Y _5142_/X _5220_/C _5157_/Y VGND VGND VPWR VPWR _5158_/Y sky130_fd_sc_hd__o211ai_4
XANTENNA__3693__C1 _3380_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4527__D _4527_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4109_ _3580_/A _3911_/B _3533_/X _3962_/X _4108_/Y VGND VGND VPWR VPWR _4109_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__4237__A1 _6125_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5089_ _5256_/A _5757_/C _5757_/D _6119_/Q _4987_/X VGND VGND VPWR VPWR _5089_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_44_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5434__B1 _5968_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3460__A2 _3876_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3996__B1 _4044_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5737__A1 _4686_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4840__A _4882_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3456__A _3966_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5572__A2_N _5985_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4712__A2 _4711_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6189__D _6189_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3920__B1 _3917_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input42_A memory_dmem_request_put[68] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3191__A _3841_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4287__A _4301_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output129_A _3033_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4228__B2 input17/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4228__A1 input9/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5610__S _5616_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_4_10_0_CLK_A clkbuf_3_5_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6112__CLK _6123_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4779__A2 _4778_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3987__B1 _3982_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5728__A1 _6112_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4172__D _4205_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5565__B _5565_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4951__A2 _4941_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3366__A _3366_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4460_ _4860_/C _4462_/A _4769_/B _4734_/A VGND VGND VPWR VPWR _4461_/A sky130_fd_sc_hd__a31o_1
XANTENNA__5900__A1 _5006_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3411_ _3870_/B VGND VGND VPWR VPWR _3527_/C sky130_fd_sc_hd__clkbuf_2
X_4391_ _5715_/B _4211_/A _4390_/X VGND VGND VPWR VPWR _4767_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__6099__D _6099_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4164__B1 _6045_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3342_ _3515_/B VGND VGND VPWR VPWR _3342_/X sky130_fd_sc_hd__clkbuf_4
X_6130_ _6207_/CLK _6130_/D VGND VGND VPWR VPWR _6130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3273_ _3437_/B _3773_/B VGND VGND VPWR VPWR _4152_/C sky130_fd_sc_hd__nor2_2
XANTENNA__5113__C1 _5112_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6061_ _6204_/CLK _6061_/D VGND VGND VPWR VPWR _6061_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4197__A _4225_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5012_ _5002_/Y _5004_/Y _5007_/X _5011_/X VGND VGND VPWR VPWR _5012_/Y sky130_fd_sc_hd__a31oi_4
XANTENNA__5664__B1 _4584_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3690__A2 _3645_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5416__B1 _5405_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5967__B2 _5966_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5967__A1 _6195_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3978__B1 _3470_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5914_ _4657_/X _5912_/Y _5004_/A _5913_/X VGND VGND VPWR VPWR _5914_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_34_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5719__A1 _4666_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5845_ _4570_/Y _4571_/X _5982_/C VGND VGND VPWR VPWR _5845_/X sky130_fd_sc_hd__o21a_2
XFILLER_34_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3993__A3 _3989_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5756__A _5756_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5776_ _4353_/X _5775_/Y _5017_/X VGND VGND VPWR VPWR _5776_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5195__A2 _5190_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2988_ _6204_/Q VGND VGND VPWR VPWR _5294_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5475__B _5501_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4727_ _5188_/C VGND VGND VPWR VPWR _5078_/B sky130_fd_sc_hd__buf_2
XANTENNA__3276__A _3657_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4658_ _4297_/X _4536_/A _4777_/A _4778_/A VGND VGND VPWR VPWR _5167_/A sky130_fd_sc_hd__o2bb2a_2
XFILLER_107_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3609_ _3609_/A _3609_/B VGND VGND VPWR VPWR _3938_/B sky130_fd_sc_hd__and2_2
XANTENNA__4155__B1 _4154_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4589_ _4589_/A VGND VGND VPWR VPWR _5680_/B sky130_fd_sc_hd__buf_4
XANTENNA__5491__A _5499_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5655__B1 _4937_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6135__CLK _6146_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4835__A _4835_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3681__A2 _3429_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5407__B1 _5162_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5958__A1 _4629_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3969__B1 _3968_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4091__C1 _3308_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5186__A2 _5180_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3197__A1 _3139_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3186__A _3447_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4933__A2 _4925_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3736__A3 _3246_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3197__B2 _3196_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5489__A3 _5405_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5894__B1 _5845_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5605__S _5605_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4729__B _4729_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4161__A3 _3910_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4449__A1 _4422_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3633__B _3710_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3125__S _3127_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5110__A2 _4328_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4449__B2 _5712_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3121__A1 _6093_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3672__A2 _3230_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5949__A1 _5946_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3960_ _3359_/A _3952_/Y _3953_/X _3959_/X _4002_/A VGND VGND VPWR VPWR _3960_/Y
+ sky130_fd_sc_hd__a311oi_1
XFILLER_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5413__A3 _5395_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4082__C1 _3756_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5576__A _5576_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3891_ _3891_/A VGND VGND VPWR VPWR _3891_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4480__A _5711_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5177__A2 _5062_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5630_ _6173_/Q _6041_/Q _5638_/S VGND VGND VPWR VPWR _5631_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5716__A4 _4556_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5561_ _5968_/C _5529_/X _5560_/X _5499_/X _6145_/Q VGND VGND VPWR VPWR _5562_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3527__C _3527_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3096__A _3096_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5492_ _4803_/X _5433_/A _5490_/X _5491_/X _6123_/Q VGND VGND VPWR VPWR _5493_/A
+ sky130_fd_sc_hd__a32o_1
X_4512_ _6126_/Q _4511_/X _4224_/A VGND VGND VPWR VPWR _4512_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4137__B1 _4152_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4443_ _4728_/A _4860_/B VGND VGND VPWR VPWR _4884_/A sky130_fd_sc_hd__nand2_2
XANTENNA__5885__B1 _5884_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4374_ _5240_/C VGND VGND VPWR VPWR _4374_/X sky130_fd_sc_hd__buf_4
XFILLER_98_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3896__C1 _3410_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6158__CLK _6201_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3325_ _3621_/D VGND VGND VPWR VPWR _3528_/A sky130_fd_sc_hd__buf_2
XANTENNA__3543__B _3543_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6113_ _6123_/CLK _6113_/D VGND VGND VPWR VPWR _6113_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _3386_/A VGND VGND VPWR VPWR _3462_/B sky130_fd_sc_hd__buf_2
XANTENNA__5101__A2 _5099_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_86_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3035__S _3043_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _6202_/CLK _6044_/D VGND VGND VPWR VPWR _6044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3112__A1 _6089_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3187_ _4004_/B VGND VGND VPWR VPWR _3195_/A sky130_fd_sc_hd__buf_2
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5404__A3 _4232_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4612__A1 _4273_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5486__A _5486_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3820__C1 _3819_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5828_ _4360_/X _5826_/X _5732_/B _5827_/X VGND VGND VPWR VPWR _5828_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5168__A2 _4290_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5759_ _5756_/X _5757_/X _5758_/Y _5739_/Y VGND VGND VPWR VPWR _5759_/Y sky130_fd_sc_hd__a22oi_2
XANTENNA__4915__A2 _4629_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3437__C _3437_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5876__B1 _5858_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3887__C1 _3886_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4626__A2_N _4571_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5891__A3 _5903_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3351__B2 _3347_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3351__A1 _3342_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3103__A1 _6085_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4565__A _4565_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4851__B2 _4850_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4603__A1 _4329_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5800__B1 _4488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4064__C1 _3508_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3709__A3 _3911_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3628__B _3748_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4906__A2 _4227_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3590__A1 _3862_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4119__B1 _3680_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5335__S _5339_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3878__C1 _3241_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3110_ _6059_/Q _6088_/Q _3116_/S VGND VGND VPWR VPWR _3111_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5619__A0 _6168_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4090_ _3299_/A _4089_/Y _3482_/X _3510_/X _3218_/X VGND VGND VPWR VPWR _4090_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5095__A1 _5089_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4842__A1 _4950_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3041_ _6038_/Q _6170_/Q _3043_/S VGND VGND VPWR VPWR _3042_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4194__B input7/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_15_0_CLK clkbuf_3_7_0_CLK/X VGND VGND VPWR VPWR _6146_/CLK sky130_fd_sc_hd__clkbuf_2
X_4992_ _5438_/C _4227_/A input9/X _5042_/A VGND VGND VPWR VPWR _4992_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4070__A2 _3975_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3943_ _3286_/X _3930_/Y _3935_/X _3941_/Y _3942_/X VGND VGND VPWR VPWR _3943_/X
+ sky130_fd_sc_hd__o32a_1
X_3874_ _3410_/B _3254_/X _3512_/A _3873_/X VGND VGND VPWR VPWR _3874_/X sky130_fd_sc_hd__o211a_1
X_5613_ _5613_/A VGND VGND VPWR VPWR _6165_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3030__A0 _6033_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5544_ _5544_/A VGND VGND VPWR VPWR _6139_/D sky130_fd_sc_hd__clkbuf_1
X_5475_ _5475_/A _5501_/B VGND VGND VPWR VPWR _5476_/A sky130_fd_sc_hd__and2_1
X_4426_ _4759_/C VGND VGND VPWR VPWR _4860_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__5858__B1 _5982_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4125__A3 _3654_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4369__B _5188_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3273__B _3773_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3869__C1 _3868_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4357_ _4738_/A VGND VGND VPWR VPWR _4865_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4088__C _4088_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4288_ _4527_/A _4298_/A _4358_/A _4354_/D VGND VGND VPWR VPWR _4578_/A sky130_fd_sc_hd__nand4_4
XFILLER_58_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3308_ _3308_/A VGND VGND VPWR VPWR _3308_/X sky130_fd_sc_hd__clkbuf_4
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5086__B2 _5085_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4385__A _4385_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3239_ _3218_/X _3223_/X _3230_/X _3238_/X VGND VGND VPWR VPWR _3239_/X sky130_fd_sc_hd__a31o_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6027_ _6197_/CLK _6027_/D VGND VGND VPWR VPWR _6027_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3097__A0 _6054_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4833__A1 _5899_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5389__A2 _4985_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4046__C1 _4045_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3939__A3 _3904_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5010__A1 _5008_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5944__A _5944_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3021__A0 _6029_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5561__A2 _5529_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3464__A _3574_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5849__B1 _5848_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3324__A1 _3305_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6197__D _6197_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5864__A3 _4953_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3875__A2 _3588_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5077__A1 _4945_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5496__A1_N _6124_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4295__A _4860_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3911__B _3911_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3088__A0 _6186_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4824__A1 _4483_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4824__B2 _5188_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4726__C _5018_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3627__A2 _3342_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4037__C1 _3673_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output111_A _3126_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4588__B1 _4696_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4052__A2 _3666_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6015__A _6015_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_4_0_CLK clkbuf_3_5_0_CLK/A VGND VGND VPWR VPWR clkbuf_4_9_0_CLK/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5434__A1_N _6108_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5001__A1 _5944_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3590_ _3862_/A _4116_/B _3588_/X _4128_/A VGND VGND VPWR VPWR _3590_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5552__A2 _4218_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5260_ _5260_/A VGND VGND VPWR VPWR _5260_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4211_ _4211_/A VGND VGND VPWR VPWR _5648_/S sky130_fd_sc_hd__buf_2
XANTENNA__4512__B1 _4224_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5191_ _5191_/A VGND VGND VPWR VPWR _5899_/A sky130_fd_sc_hd__buf_2
XFILLER_68_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4917__B _5761_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4142_ _3406_/A _4073_/C _3631_/A _3841_/B _4149_/A VGND VGND VPWR VPWR _4143_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4073_ _4073_/A _4073_/B _4073_/C _4073_/D VGND VGND VPWR VPWR _4073_/X sky130_fd_sc_hd__or4_4
XFILLER_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3079__A0 _6182_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3024_ _6030_/Q _6162_/Q _3032_/S VGND VGND VPWR VPWR _3025_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4028__C1 _4048_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4975_ _4975_/A VGND VGND VPWR VPWR _4975_/X sky130_fd_sc_hd__buf_2
X_3926_ _4048_/A VGND VGND VPWR VPWR _3926_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__4043__A2 _4042_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3549__A _3549_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4594__A3 _5029_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3268__B _3359_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3857_ _3666_/X _3830_/D _3342_/X _3653_/B _3447_/X VGND VGND VPWR VPWR _3857_/Y
+ sky130_fd_sc_hd__a41oi_2
XANTENNA__4658__A1_N _4297_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3788_ _3777_/Y _3638_/Y _3778_/X _3785_/X _3787_/X VGND VGND VPWR VPWR _3788_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4751__B1 _4956_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5527_ _4801_/X _4268_/B _5092_/X _5504_/A _4277_/Y VGND VGND VPWR VPWR _5528_/A
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3554__B2 _3553_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3554__A1 _3549_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5458_ input21/X _5437_/A _5439_/A input13/X VGND VGND VPWR VPWR _5767_/C sky130_fd_sc_hd__a22o_1
X_4409_ _4404_/X _4405_/X _4864_/C _4864_/D _4369_/C VGND VGND VPWR VPWR _4409_/X
+ sky130_fd_sc_hd__o221a_4
XFILLER_59_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5389_ _4246_/A _4985_/A _4246_/C _4859_/D VGND VGND VPWR VPWR _5432_/A sky130_fd_sc_hd__o31a_2
XANTENNA__3857__A2 _3830_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5059__A1 _5058_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3731__B _3873_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5004__A _5004_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4806__A1 _4716_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6008__B1 _6011_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4843__A _4843_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3490__B1 _3488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5231__A1 _5018_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3459__A _3983_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3178__B _3468_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3793__A1 _3673_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5674__A _5674_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4990__B1 _4976_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input72_A memory_dmem_request_put[98] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3194__A _4089_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5570__A_N _6200_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5298__A1 _6065_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3848__A2 _3881_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4456__C _4780_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5470__A1 input24/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4753__A _5211_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5470__B2 _5431_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5568__B _5568_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4025__A2 _3457_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3369__A _4042_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _4876_/A VGND VGND VPWR VPWR _4956_/D sky130_fd_sc_hd__buf_4
XANTENNA__4430__C1 _4955_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4576__A3 _4852_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5773__A2 _4721_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4691_ _4686_/X _5755_/D _5829_/C _4690_/Y VGND VGND VPWR VPWR _4691_/X sky130_fd_sc_hd__o211a_1
X_3711_ _3711_/A _3711_/B _3746_/A VGND VGND VPWR VPWR _3711_/X sky130_fd_sc_hd__or3b_4
XANTENNA__3784__A1 _3783_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5584__A _5584_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4981__B1 _4224_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3642_ _3642_/A _3648_/B VGND VGND VPWR VPWR _3938_/C sky130_fd_sc_hd__nor2_8
XANTENNA__3816__B _3816_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3573_ _3895_/A VGND VGND VPWR VPWR _3573_/X sky130_fd_sc_hd__buf_2
X_5312_ _5312_/A VGND VGND VPWR VPWR _6071_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5289__A1 _5285_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5243_ _4855_/A _5971_/A _4917_/A _5179_/A _5829_/A VGND VGND VPWR VPWR _5243_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4928__A _4928_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5174_ _5168_/Y _5169_/Y _5172_/Y _5173_/X VGND VGND VPWR VPWR _5174_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__3832__A _3832_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3839__A2 _3636_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4125_ _3178_/X _3767_/B _3654_/X _3359_/B _3904_/D VGND VGND VPWR VPWR _4126_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_96_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3043__S _3043_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4056_ _3603_/B _3300_/X _3580_/X _4055_/X _3302_/X VGND VGND VPWR VPWR _4056_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_83_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3007_ _3007_/A VGND VGND VPWR VPWR _3007_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5749__C1 _5748_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5213__A1 _4580_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3279__A _3279_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4016__A2 _3829_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4958_ _4954_/X _4956_/Y _4957_/X VGND VGND VPWR VPWR _4958_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5764__A2 _5763_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4889_ _4886_/Y _5732_/B _4888_/X _4420_/A VGND VGND VPWR VPWR _4889_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4972__B1 _5125_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3775__B2 _3764_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3775__A1 _3815_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3909_ _3286_/X _3899_/X _4088_/D _3909_/D VGND VGND VPWR VPWR _3909_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__5494__A _5494_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5516__A2 _5433_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4724__B1 _5048_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5921__C1 _5920_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5909__A1_N _6192_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3461__B _3461_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4255__A2 _4244_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5452__A1 _4977_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3463__B1 _3460_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5452__B2 _6111_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5388__B _5388_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3189__A _3344_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4007__A2 _3720_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5204__A1 _5201_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4963__B1 _4962_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3766__A1 _3764_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3766__B2 _3815_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5608__S _5616_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5507__A2 _4632_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5912__C1 _4956_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6041__CLK _6202_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6191__CLK _6196_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5570__C _5570_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5691__B2 _5690_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3802__D _3802_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4483__A _4483_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5930_ _5926_/X _5927_/Y _5929_/Y VGND VGND VPWR VPWR _5930_/X sky130_fd_sc_hd__o21a_1
XFILLER_34_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5994__A2 _5998_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3454__B1 _6018_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5861_ _5706_/B _5706_/C _5032_/Y _5068_/X _4765_/A VGND VGND VPWR VPWR _5861_/Y
+ sky130_fd_sc_hd__a41oi_1
XFILLER_34_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4812_ _4843_/A _4843_/C _5078_/A _5761_/B VGND VGND VPWR VPWR _4812_/X sky130_fd_sc_hd__o211a_2
X_5792_ _4927_/X _5712_/A _5782_/X _5720_/A _5752_/Y VGND VGND VPWR VPWR _5792_/Y
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA__4954__B1 _4953_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4743_ _4739_/X _4740_/X _4931_/A _4742_/X VGND VGND VPWR VPWR _4743_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__3757__A1 _3689_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5745__C _5745_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4674_ _5067_/A VGND VGND VPWR VPWR _4675_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5708__A2_N _5706_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3625_ _3613_/X _3623_/X _3624_/X VGND VGND VPWR VPWR _3625_/X sky130_fd_sc_hd__a21o_1
X_3556_ _4105_/B VGND VGND VPWR VPWR _3628_/A sky130_fd_sc_hd__buf_2
XANTENNA__5761__B _5761_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3487_ _4073_/B VGND VGND VPWR VPWR _4044_/A sky130_fd_sc_hd__buf_2
XANTENNA__3562__A _3562_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5226_ _6124_/Q _4807_/X _5013_/X VGND VGND VPWR VPWR _5226_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5682__A1 _4345_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5157_ _5150_/Y _5156_/X _4767_/X VGND VGND VPWR VPWR _5157_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_69_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3693__B1 _3429_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4108_ _4105_/X _4107_/X _3242_/X VGND VGND VPWR VPWR _4108_/Y sky130_fd_sc_hd__a21oi_1
X_5088_ _5093_/A VGND VGND VPWR VPWR _5256_/A sky130_fd_sc_hd__buf_2
XFILLER_71_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4393__A _4685_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4039_ _4039_/A _4039_/B VGND VGND VPWR VPWR _4039_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5434__B2 _5433_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3445__B1 _3588_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3996__B2 _3849_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5737__A2 _4604_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6064__CLK _6201_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5370__B1 _5381_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4568__A _4767_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3920__A1 _3477_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5122__B1 _5121_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3472__A _3647_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5658__D1 _4965_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4287__B _4287_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3684__B1 _3580_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input35_A memory_dmem_request_put[61] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4881__C1 _4880_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4228__A2 _4717_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3987__A1 _3357_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5189__B1 _4582_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5728__A2 _4511_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3647__A _3647_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3366__B _3440_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4427__A1_N _4313_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4390_ _4243_/A _4985_/A _4986_/A _6140_/Q VGND VGND VPWR VPWR _4390_/X sky130_fd_sc_hd__o31a_4
X_3410_ _3410_/A _3410_/B VGND VGND VPWR VPWR _3934_/D sky130_fd_sc_hd__nor2_1
XANTENNA__5361__A0 _6050_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4164__B2 _3891_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4164__A1 _4157_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3341_ _3468_/B VGND VGND VPWR VPWR _3515_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__5900__A2 _5026_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4478__A _4788_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3382__A _3841_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3272_ _3272_/A _3330_/A VGND VGND VPWR VPWR _3773_/B sky130_fd_sc_hd__or2b_4
XANTENNA__5113__B1 _4746_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5664__A1 _4644_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4197__B _4227_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6060_ _6207_/CLK _6060_/D VGND VGND VPWR VPWR _6060_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _4644_/X _4642_/X _5010_/X _4584_/X VGND VGND VPWR VPWR _5011_/X sky130_fd_sc_hd__o31a_2
XANTENNA__3675__B1 _3724_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5416__A1 input12/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5102__A _5102_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5967__A2 _4799_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3978__A1 _4089_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5913_ _4332_/X _5080_/X _5098_/X _4931_/A VGND VGND VPWR VPWR _5913_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6087__CLK _6176_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5719__A2 _4582_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5844_ _5235_/X _4927_/X _5712_/A _4420_/X VGND VGND VPWR VPWR _5844_/X sky130_fd_sc_hd__a31o_1
X_5775_ _5761_/D _5878_/B _5118_/D VGND VGND VPWR VPWR _5775_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3557__A _3557_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2987_ _2987_/A VGND VGND VPWR VPWR _2987_/X sky130_fd_sc_hd__clkbuf_1
X_4726_ _4726_/A _5148_/C _5018_/D VGND VGND VPWR VPWR _4732_/A sky130_fd_sc_hd__and3_1
XFILLER_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4657_ _4657_/A VGND VGND VPWR VPWR _4657_/X sky130_fd_sc_hd__buf_2
X_3608_ _3756_/A _3779_/C _4042_/A VGND VGND VPWR VPWR _3608_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4155__A1 _3666_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput80 memory_imem_request_put[6] VGND VGND VPWR VPWR _3275_/B sky130_fd_sc_hd__buf_4
XANTENNA__5772__A _5772_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4588_ _4404_/X _4405_/X _4696_/A VGND VGND VPWR VPWR _4589_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__3363__C1 _4004_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3292__A _3366_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3539_ _3535_/X _3536_/X _3537_/X _3816_/A VGND VGND VPWR VPWR _3539_/X sky130_fd_sc_hd__o31a_1
XFILLER_89_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5104__B1 _4584_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5655__A1 _4459_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5209_ _5207_/X _5208_/X _4859_/X _4858_/Y VGND VGND VPWR VPWR _5209_/X sky130_fd_sc_hd__o2bb2a_1
X_6189_ _6205_/CLK _6189_/D VGND VGND VPWR VPWR _6189_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4863__C1 _5721_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3681__A3 _3679_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5407__A1 _5640_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5407__B2 _4800_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5958__A2 _4975_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3969__A1 _3967_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4091__B1 _3293_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3467__A _4065_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3197__A2 _3142_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5894__A1 _5882_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4729__C _4926_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4298__A _4298_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4449__A2 _4423_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output141_A _3055_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5621__S _5627_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5949__A2 _5955_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4237__S _4633_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4082__B1 _4124_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4761__A _4946_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3890_ _3357_/X _6033_/Q _3880_/Y _3889_/X VGND VGND VPWR VPWR _6033_/D sky130_fd_sc_hd__a211o_1
XANTENNA__4366__A1_N _4527_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4480__B _4725_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5560_ _5437_/A _5439_/A _4976_/A VGND VGND VPWR VPWR _5560_/X sky130_fd_sc_hd__o21a_1
X_4511_ _5772_/A VGND VGND VPWR VPWR _4511_/X sky130_fd_sc_hd__clkbuf_2
X_5491_ _5499_/A VGND VGND VPWR VPWR _5491_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4442_ _4442_/A VGND VGND VPWR VPWR _4728_/A sky130_fd_sc_hd__buf_2
XANTENNA__4137__B2 _4061_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4137__A1 _3835_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5885__A1 _4870_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4373_ _4643_/A VGND VGND VPWR VPWR _5240_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__3896__B1 _3403_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3324_ _3305_/X _3308_/X _3314_/Y _3320_/Y _4146_/A VGND VGND VPWR VPWR _3324_/X
+ sky130_fd_sc_hd__a311o_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6112_ _6123_/CLK _6112_/D VGND VGND VPWR VPWR _6112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4936__A _4936_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3255_ _3461_/A _3272_/A VGND VGND VPWR VPWR _3386_/A sky130_fd_sc_hd__nand2_1
XFILLER_86_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _6045_/CLK _6043_/D VGND VGND VPWR VPWR _6043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _3447_/C VGND VGND VPWR VPWR _4004_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_26_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4671__A _5003_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4612__A2 _4211_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5767__A _5805_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5486__B _5501_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3820__B1 _3763_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5827_ _5152_/A _5971_/C _4953_/X _5721_/C VGND VGND VPWR VPWR _5827_/X sky130_fd_sc_hd__a211o_1
X_5758_ _4422_/X _4423_/X _4822_/X _5033_/Y VGND VGND VPWR VPWR _5758_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__4915__A3 _4630_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4709_ _4702_/A _5152_/A _4891_/A _4708_/D VGND VGND VPWR VPWR _4709_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3584__C1 _3583_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5689_ _5757_/B _5013_/S _4882_/X _4652_/A _5756_/A VGND VGND VPWR VPWR _5690_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__6102__CLK _6146_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3887__B1 _3476_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5876__B2 _5875_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3351__A2 _3343_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5089__C1 _4987_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3639__B1 _3638_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4581__A _5034_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4603__A2 _4330_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5800__A1 _4317_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5800__B2 _5240_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4064__B1 _3699_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5261__C1 _4804_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5677__A _5772_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3811__B1 _6029_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3709__A4 _4065_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3628__C _3628_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5564__B1 _4987_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3575__C1 _3574_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4119__A1 _3314_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5616__S _5616_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3590__A2 _4116_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3878__B1 _3877_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5619__A1 _6036_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3660__A _3841_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_67_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5095__A2 _4991_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3040_ _3040_/A VGND VGND VPWR VPWR _3040_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4842__A2 _4841_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4194__C _5438_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5252__C1 _4950_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4055__B1 _4052_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4991_ _5715_/A _5968_/B _4990_/X _5924_/A VGND VGND VPWR VPWR _4991_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5587__A _5587_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3942_ _3940_/X _3492_/X _3806_/A VGND VGND VPWR VPWR _3942_/X sky130_fd_sc_hd__a21bo_1
X_3873_ _3983_/A _3873_/B _3966_/C VGND VGND VPWR VPWR _3873_/X sky130_fd_sc_hd__or3_1
X_5612_ _6165_/Q _6033_/Q _5616_/S VGND VGND VPWR VPWR _5613_/A sky130_fd_sc_hd__mux2_1
X_5543_ _5543_/A _5568_/B VGND VGND VPWR VPWR _5544_/A sky130_fd_sc_hd__and2_1
XANTENNA__6125__CLK _6147_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3835__A _3835_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3030__A1 _6165_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5858__A1 _5734_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5474_ _5508_/A VGND VGND VPWR VPWR _5501_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4425_ _4566_/A VGND VGND VPWR VPWR _4640_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3869__B1 _3603_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3046__S _3054_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4369__C _4369_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4356_ _4369_/D VGND VGND VPWR VPWR _5140_/B sky130_fd_sc_hd__buf_2
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3307_ _3797_/A VGND VGND VPWR VPWR _3308_/A sky130_fd_sc_hd__buf_2
XANTENNA__4088__D _4088_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4666__A _4666_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4287_ _4301_/A _4287_/B _4405_/C _4405_/D VGND VGND VPWR VPWR _4354_/D sky130_fd_sc_hd__nand4_4
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4294__B1 _4234_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3238_ _3509_/A _3557_/A _3549_/A _3847_/B VGND VGND VPWR VPWR _3238_/X sky130_fd_sc_hd__and4b_1
XFILLER_39_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ _6045_/CLK _6026_/D VGND VGND VPWR VPWR _6026_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3097__A1 _6082_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4833__A2 _4843_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3169_ _3278_/A VGND VGND VPWR VPWR _4065_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5389__A3 _4246_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4046__B1 _3838_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5794__B1 _5721_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5546__B1 _6140_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5010__A2 _5009_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5944__B _5944_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4826__A1_N _4821_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5561__A3 _5560_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3021__A1 _6161_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5849__A1 _6190_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3324__A2 _3308_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3480__A _3480_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5077__A2 _5076_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3911__C _3911_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3088__A1 _6078_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4824__A2 _4485_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5234__C1 _4652_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4037__B1 _3882_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5785__B1 _4924_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4588__A1 _4404_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output104_A _3113_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6148__CLK _6197_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4052__A3 _3844_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5001__A2 _5971_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5552__A3 _5260_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5346__S _5350_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4210_ _5818_/S VGND VGND VPWR VPWR _4211_/A sky130_fd_sc_hd__buf_4
XFILLER_5_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4512__A1 _6126_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5190_ _4347_/A _4673_/B _4960_/A _5022_/A VGND VGND VPWR VPWR _5190_/X sky130_fd_sc_hd__a31o_2
XANTENNA__4486__A _4738_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3390__A _3522_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4141_ _4134_/X _4140_/Y _3290_/X _6044_/Q _3891_/X VGND VGND VPWR VPWR _6044_/D
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4917__C _5878_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4072_ _4064_/Y _4071_/X _3624_/X VGND VGND VPWR VPWR _4072_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3079__A1 _6074_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3023_ _3056_/S VGND VGND VPWR VPWR _3032_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_64_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4028__B1 _3444_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5225__C1 _5260_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5776__B1 _5017_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4974_ _4974_/A _4974_/B _4974_/C VGND VGND VPWR VPWR _4974_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__4043__A3 _3279_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3925_ _3195_/B _3831_/X _3342_/X _3653_/B _3924_/X VGND VGND VPWR VPWR _3925_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__4594__A4 _5021_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3856_ _3840_/Y _3855_/X _3821_/X _6032_/Q _3822_/X VGND VGND VPWR VPWR _6032_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_118_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3565__A _3858_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3787_ _4088_/D VGND VGND VPWR VPWR _3787_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4751__A1 _4488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3554__A2 _3767_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5526_ _5526_/A VGND VGND VPWR VPWR _6133_/D sky130_fd_sc_hd__clkbuf_1
X_5457_ _5444_/X _5445_/X _5455_/X _5447_/X _5456_/X VGND VGND VPWR VPWR _6112_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4408_ _4533_/A VGND VGND VPWR VPWR _4864_/D sky130_fd_sc_hd__buf_2
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5700__B1 _5679_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5388_ _5388_/A _5388_/B VGND VGND VPWR VPWR _6100_/D sky130_fd_sc_hd__nor2_1
XANTENNA__4396__A _4734_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4339_ _5687_/A _5687_/B _4328_/X _4332_/X _5179_/A VGND VGND VPWR VPWR _4339_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_101_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3857__A3 _3342_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3731__C _3966_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5059__A2 _5944_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5004__B _5731_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4806__A2 _4513_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6009_ _6009_/A _6013_/B _5293_/X VGND VGND VPWR VPWR _6011_/A sky130_fd_sc_hd__or3b_1
XANTENNA__6008__A1 _6143_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4843__B _4843_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5216__C1 _5215_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4019__B1 _3520_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3490__A1 _3536_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5231__A2 _5021_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5020__A _5020_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5955__A _5955_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3793__A2 _3293_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4990__A1 _4804_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5674__B _5674_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3950__C1 _3949_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input65_A memory_dmem_request_put[91] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5690__A _5690_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_4_14_0_CLK clkbuf_3_7_0_CLK/X VGND VGND VPWR VPWR _6145_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_111_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3848__A3 _3195_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4456__D _4623_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5470__A2 _5437_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3982__B_N _3976_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5758__B1 _4822_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3369__B _3686_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4430__B1 _4640_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3710_ _3998_/A _3719_/B _3710_/C _3611_/A VGND VGND VPWR VPWR _3710_/X sky130_fd_sc_hd__or4b_1
X_4690_ _5745_/C _5667_/B _4581_/C VGND VGND VPWR VPWR _4690_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3784__A2 _3734_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2992__A0 _6017_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4981__A1 _6132_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3641_ _4149_/B VGND VGND VPWR VPWR _4135_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3385__A _3686_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3572_ _3572_/A VGND VGND VPWR VPWR _3910_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__5930__B1 _5929_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3816__C _3816_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5311_ _6195_/Q _6071_/Q _5317_/S VGND VGND VPWR VPWR _5312_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5289__A2 _5286_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5242_ _5239_/X _5240_/X _5241_/X _4836_/X VGND VGND VPWR VPWR _5242_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4497__B1 _4390_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5173_ _4673_/Y _4398_/X _5102_/D _4959_/X _5140_/C VGND VGND VPWR VPWR _5173_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_68_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3839__A3 _3249_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4124_ _4124_/A _4124_/B _4124_/C _4124_/D VGND VGND VPWR VPWR _4124_/X sky130_fd_sc_hd__or4_1
XFILLER_29_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4249__B1 _6139_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput1 EN_memory_dmem_request_put VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__buf_6
X_4055_ _4126_/B _4049_/Y _4051_/X _4052_/Y _4054_/X VGND VGND VPWR VPWR _4055_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__5997__B1 _6201_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3006_ _6022_/Q _6154_/Q _3010_/S VGND VGND VPWR VPWR _3007_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5749__B1 _5673_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5213__A2 _4878_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4957_ _4957_/A VGND VGND VPWR VPWR _4957_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4888_ _4488_/X _4887_/X _5761_/B _5687_/C _5240_/C VGND VGND VPWR VPWR _4888_/X
+ sky130_fd_sc_hd__a221o_1
X_3908_ _3340_/X _3901_/Y _3903_/Y _3695_/B _3907_/Y VGND VGND VPWR VPWR _3909_/D
+ sky130_fd_sc_hd__a311o_2
XANTENNA__4972__A1 _4524_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3775__A2 _3765_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3839_ _3536_/X _3636_/X _3249_/X _3838_/X VGND VGND VPWR VPWR _3839_/X sky130_fd_sc_hd__o31a_2
XFILLER_20_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3295__A _3983_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4724__A1 _4692_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5921__B1 _4964_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5198__B1_N _5015_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5509_ _5509_/A _5531_/B VGND VGND VPWR VPWR _5510_/A sky130_fd_sc_hd__and2_1
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5015__A _5015_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_3_0_CLK clkbuf_3_3_0_CLK/A VGND VGND VPWR VPWR clkbuf_4_7_0_CLK/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4854__A _4854_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3463__A1 _3543_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4255__A3 _4264_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5452__A2 _5412_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4660__B1 _4580_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3463__B2 _3761_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5204__A2 _5202_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4963__A1 _4487_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3766__A2 _3634_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5507__A3 _5498_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5912__B1 _4345_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4764__A _4875_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5979__B1 _5063_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3454__A1 _3396_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5860_ _4890_/A _5018_/B _4761_/X _5123_/B VGND VGND VPWR VPWR _5860_/X sky130_fd_sc_hd__o211a_1
XFILLER_34_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3454__B2 _3357_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4811_ _4811_/A VGND VGND VPWR VPWR _5761_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_92_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5791_ _6187_/Q VGND VGND VPWR VPWR _5791_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5595__A _5595_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4954__A1 _4680_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4742_ _4742_/A VGND VGND VPWR VPWR _4742_/X sky130_fd_sc_hd__buf_2
XANTENNA__3757__A2 _3663_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4673_ _4673_/A _4673_/B VGND VGND VPWR VPWR _4673_/Y sky130_fd_sc_hd__nand2_4
X_3624_ _3806_/A VGND VGND VPWR VPWR _3624_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__4004__A _4004_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3555_ _3687_/B VGND VGND VPWR VPWR _4105_/B sky130_fd_sc_hd__buf_2
XANTENNA__5761__C _5761_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3486_ _3871_/B VGND VGND VPWR VPWR _3975_/B sky130_fd_sc_hd__buf_2
X_5225_ _5201_/X _5224_/Y _5968_/C _5260_/A VGND VGND VPWR VPWR _5225_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5682__A2 _5213_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3054__S _3054_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5156_ _5151_/Y _5154_/X _5155_/Y VGND VGND VPWR VPWR _5156_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3693__A1 _3659_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4674__A _5067_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4107_ _3537_/B _4106_/X _3509_/Y _4040_/X VGND VGND VPWR VPWR _4107_/X sky130_fd_sc_hd__o22a_1
X_5087_ _5757_/A VGND VGND VPWR VPWR _5093_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3445__A1 _3719_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4038_ _3583_/A _4037_/X _3990_/X _4014_/X VGND VGND VPWR VPWR _4039_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5198__A1 _5196_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5989_ _5989_/A VGND VGND VPWR VPWR _6197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3507__B1_N _4088_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5370__A1 _4189_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3920__A2 _3831_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5658__C1 _4672_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5122__B2 _4744_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4287__C _4405_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4881__B1 _4875_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3684__A1 _3681_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4584__A _4584_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input28_A memory_dmem_request_put[54] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4633__A0 _4632_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3987__A2 _6037_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5189__A1 _4374_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5619__S _5627_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4759__A _4759_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output96_A _3098_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5361__A1 _6094_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4164__A2 _4163_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5900__A3 _5899_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3663__A _3663_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3340_ _3546_/A VGND VGND VPWR VPWR _3340_/X sky130_fd_sc_hd__buf_2
XANTENNA__5113__A1 _4836_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3382__B _4149_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5649__C1 _5163_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5010_ _5008_/X _5009_/X _4353_/A _5711_/B VGND VGND VPWR VPWR _5010_/X sky130_fd_sc_hd__a211o_1
X_3271_ _3271_/A VGND VGND VPWR VPWR _3359_/B sky130_fd_sc_hd__buf_2
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5664__A2 _4642_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3675__A1 _3673_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4494__A _5140_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5416__A2 _5395_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5102__B _5102_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5821__C1 _5820_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3978__A2 _3512_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5912_ _4672_/X _5167_/X _4345_/X _4956_/Y VGND VGND VPWR VPWR _5912_/Y sky130_fd_sc_hd__o211ai_2
X_5843_ _5176_/X _4971_/X _4793_/X _5842_/X _5031_/X VGND VGND VPWR VPWR _5843_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_61_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5719__A3 _5717_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3838__A _3838_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5774_ _5676_/X _5773_/X _5769_/X VGND VGND VPWR VPWR _5774_/Y sky130_fd_sc_hd__a21oi_1
X_2986_ _5640_/D _2986_/B _2986_/C VGND VGND VPWR VPWR _2987_/A sky130_fd_sc_hd__and3b_4
X_4725_ _4725_/A VGND VGND VPWR VPWR _5018_/D sky130_fd_sc_hd__buf_4
X_4656_ _4656_/A VGND VGND VPWR VPWR _4657_/A sky130_fd_sc_hd__clkbuf_2
X_4587_ _4811_/A VGND VGND VPWR VPWR _4996_/A sky130_fd_sc_hd__clkbuf_4
X_3607_ _3781_/C _3609_/B _3781_/A _3781_/B VGND VGND VPWR VPWR _3607_/X sky130_fd_sc_hd__and4bb_2
XANTENNA__4155__A2 _3308_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput81 memory_imem_request_put[7] VGND VGND VPWR VPWR _3754_/B sky130_fd_sc_hd__buf_6
Xinput70 memory_dmem_request_put[96] VGND VGND VPWR VPWR _4219_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__5772__B _5772_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3573__A _3895_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3363__B1 _3382_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3538_ _3538_/A VGND VGND VPWR VPWR _3816_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3292__B _3432_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5104__A1 _4998_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3469_ _3609_/B VGND VGND VPWR VPWR _3611_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5655__A2 _4461_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5208_ _4882_/X _4461_/X _4931_/A _4785_/X VGND VGND VPWR VPWR _5208_/X sky130_fd_sc_hd__a31o_1
XFILLER_57_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6188_ _6205_/CLK _6188_/D VGND VGND VPWR VPWR _6188_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__4863__B1 _5240_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5139_ _4859_/D _4333_/A _4518_/A _4786_/X _5118_/A VGND VGND VPWR VPWR _5140_/D
+ sky130_fd_sc_hd__a311o_4
XFILLER_57_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5407__A2 _2986_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4615__B1 _4728_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6031__CLK _6197_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3969__A2 _3444_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4091__A1 _3194_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4091__B2 _3975_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3743__A1_N _3734_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3748__A _3748_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3467__B _4042_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6181__CLK _6196_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3197__A3 _3157_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4579__A _4878_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5879__C1 _5782_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5894__A2 _5886_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5203__A _5203_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output134_A _3042_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4606__B1 _4395_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4082__A1 _3831_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4480__C _4480_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4790__C1 _4789_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5490_ input31/X _4978_/X _5042_/X _4906_/X VGND VGND VPWR VPWR _5490_/X sky130_fd_sc_hd__a22o_1
X_4510_ _5648_/S VGND VGND VPWR VPWR _5772_/A sky130_fd_sc_hd__clkbuf_2
X_4441_ _4769_/A _4769_/C VGND VGND VPWR VPWR _4549_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4489__A _4769_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4137__A2 _3305_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5885__A2 _5859_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3896__A1 _3895_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4372_ _4415_/A VGND VGND VPWR VPWR _4643_/A sky130_fd_sc_hd__clkbuf_4
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ _6123_/CLK _6111_/D VGND VGND VPWR VPWR _6111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3323_ _3992_/A VGND VGND VPWR VPWR _4146_/A sky130_fd_sc_hd__buf_2
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3254_ _3847_/A VGND VGND VPWR VPWR _3254_/X sky130_fd_sc_hd__buf_2
XFILLER_39_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ _6045_/CLK _6042_/D VGND VGND VPWR VPWR _6042_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4845__B1 _4696_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6054__CLK _6205_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3185_ _3442_/B _3440_/A VGND VGND VPWR VPWR _3447_/C sky130_fd_sc_hd__or2b_2
XFILLER_81_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4952__A _4952_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5767__B _5805_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3820__A1 _3760_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5826_ _4843_/A _5899_/C _4945_/A _4565_/A _4879_/A VGND VGND VPWR VPWR _5826_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5757_ _5757_/A _5757_/B _5757_/C _5757_/D VGND VGND VPWR VPWR _5757_/X sky130_fd_sc_hd__or4_4
XFILLER_108_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4708_ _4708_/A _5152_/A _4891_/A _4708_/D VGND VGND VPWR VPWR _4708_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__3584__B1 _3548_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5688_ _5653_/Y _5687_/X _5235_/X VGND VGND VPWR VPWR _5690_/C sky130_fd_sc_hd__o21ai_2
X_4639_ _4929_/B VGND VGND VPWR VPWR _5745_/A sky130_fd_sc_hd__buf_2
XANTENNA__3887__A1 _3717_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5089__B1 _6119_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3639__A1 _3628_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4862__A _4862_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4064__A1 _4058_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5800__A2 _4363_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4064__B2 _4063_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5261__B1 _4718_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5677__B _5772_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4581__B _5711_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3811__A1 _3806_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3811__B2 _3728_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5013__A0 _4990_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3909__C _4088_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5564__A1 _5256_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5564__B2 _5482_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3575__B1 _3573_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4119__A2 _3654_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3590__A3 _3588_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4102__A _4102_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3878__A1 _3548_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6077__CLK _6203_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5632__S _5638_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3660__B _3660_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4772__A _4772_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4055__A1 _4126_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5252__B1 _5251_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4055__B2 _4054_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4990_ _4804_/A _5042_/A _4976_/A VGND VGND VPWR VPWR _4990_/X sky130_fd_sc_hd__o21a_2
XANTENNA__3388__A _3582_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3941_ _3562_/X _3359_/B _3482_/X _3940_/X VGND VGND VPWR VPWR _3941_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3872_ _4083_/C _3460_/X _3161_/A _3871_/X VGND VGND VPWR VPWR _3872_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5555__A1 _2986_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5611_ _5611_/A VGND VGND VPWR VPWR _6164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5542_ _5523_/X _5757_/B _5529_/X _5491_/X _6139_/Q VGND VGND VPWR VPWR _5543_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5473_ _4994_/X _5405_/A _5503_/A _6117_/Q VGND VGND VPWR VPWR _5475_/A sky130_fd_sc_hd__a2bb2o_1
X_4424_ _4860_/B VGND VGND VPWR VPWR _4926_/C sky130_fd_sc_hd__buf_2
XANTENNA__3869__A1 _3867_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5858__A2 _5856_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4355_ _4729_/B VGND VGND VPWR VPWR _4369_/D sky130_fd_sc_hd__buf_4
XANTENNA__4369__D _4369_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3306_ _3687_/A VGND VGND VPWR VPWR _3797_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4818__B1 _4817_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4286_ _4293_/A _4246_/A _4308_/A _4246_/C _6133_/Q VGND VGND VPWR VPWR _4358_/A
+ sky130_fd_sc_hd__o41ai_4
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _3983_/B VGND VGND VPWR VPWR _3847_/B sky130_fd_sc_hd__buf_2
XFILLER_73_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4294__B2 _6133_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4294__A1 _4313_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ _6045_/CLK _6025_/D VGND VGND VPWR VPWR _6025_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4833__A3 _5118_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3168_ _3632_/A VGND VGND VPWR VPWR _3648_/A sky130_fd_sc_hd__buf_2
XFILLER_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5243__B1 _5179_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4046__A1 _3962_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3099_ _6055_/Q _6083_/Q _3105_/S VGND VGND VPWR VPWR _3100_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5794__B2 _5793_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3298__A _3353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5546__A1 _5093_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5546__B2 _5482_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5809_ _5045_/A _5470_/X _5403_/X _5163_/X VGND VGND VPWR VPWR _5809_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5944__C _5944_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5018__A _5018_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5849__A2 _4629_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3324__A3 _3314_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3761__A _3761_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5739__A1_N _4665_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4809__B1 _4808_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4995__A1_N _4988_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4592__A _4614_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input10_A memory_dmem_request_put[36] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5234__B1 _4945_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4037__A1 _3475_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4037__B2 _3902_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5785__A1 _5102_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4588__A2 _4405_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3001__A _3056_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3796__B1 _6028_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4745__C1 _4744_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5001__A3 _5944_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5627__S _5627_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4767__A _4767_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4512__A2 _4511_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4140_ _3760_/X _3919_/X _3142_/X _4139_/X _3828_/X VGND VGND VPWR VPWR _4140_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_122_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4917__D _5079_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4071_ _4067_/Y _3546_/X _3695_/B _4069_/X _4070_/X VGND VGND VPWR VPWR _4071_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_83_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3022_ _3022_/A VGND VGND VPWR VPWR _3022_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5473__B1 _5503_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5598__A _5598_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4028__B2 _3902_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4028__A1 _3679_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5225__B1 _5968_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5776__A1 _4353_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4973_ _4973_/A _4973_/B VGND VGND VPWR VPWR _4974_/B sky130_fd_sc_hd__nand2_1
X_3924_ _3581_/A _3882_/C _3674_/C _3860_/A VGND VGND VPWR VPWR _3924_/X sky130_fd_sc_hd__a31o_1
XFILLER_51_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3855_ _3846_/X _3854_/X _3142_/X VGND VGND VPWR VPWR _3855_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3539__B1 _3816_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3786_ _3786_/A VGND VGND VPWR VPWR _4088_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4751__A2 _5021_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3554__A3 _3499_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5525_ _5525_/A _5531_/B VGND VGND VPWR VPWR _5526_/A sky130_fd_sc_hd__and2_1
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5456_ _6112_/Q _5222_/X _5256_/X _5260_/X VGND VGND VPWR VPWR _5456_/X sky130_fd_sc_hd__o22a_1
XFILLER_105_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4407_ _4926_/B VGND VGND VPWR VPWR _4864_/C sky130_fd_sc_hd__buf_2
XANTENNA__3581__A _3581_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5700__B2 _5699_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5387_ _5387_/A VGND VGND VPWR VPWR _6099_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4338_ _4742_/A VGND VGND VPWR VPWR _5179_/A sky130_fd_sc_hd__buf_2
XFILLER_59_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3857__A4 _3653_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3731__D _3731_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_86_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4269_ _4313_/A _4268_/Y _4234_/A _6134_/Q VGND VGND VPWR VPWR _4759_/A sky130_fd_sc_hd__a22oi_4
XANTENNA__5059__A3 _4420_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input2_A EN_memory_dmem_response_get VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5004__C _5973_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6008_ _6143_/Q _4975_/X _5367_/Y _6011_/B _4715_/X VGND VGND VPWR VPWR _6205_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__5464__B1 _5256_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4806__A3 input38/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6008__A2 _4975_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4843__C _4843_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5216__B1 _4964_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4019__B2 _4135_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4019__A1 _3183_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3490__A2 _3975_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5301__A _5301_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5231__A3 _5028_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5955__B _5955_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3756__A _3756_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5033__A1_N _4786_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4990__A2 _5042_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5674__C _5725_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3475__B _3674_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5971__A _5971_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3950__B1 _4146_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5690__B _5746_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input58_A memory_dmem_request_put[84] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4587__A _4811_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3491__A _3491_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5455__B1 _5439_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6115__CLK _6123_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3466__C1 _3465_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5211__A _5211_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5207__B1 _4345_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5758__A1 _4422_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5758__B2 _5033_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3369__C _3756_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3769__B1 _3492_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4242__A1_N _4224_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4430__A1 _4738_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3666__A _3666_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5357__S _5361_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4981__A2 _4807_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3640_ _3625_/X _3639_/X _3453_/X _6021_/Q _3541_/X VGND VGND VPWR VPWR _6021_/D
+ sky130_fd_sc_hd__a32o_1
XANTENNA__2992__A1 _6148_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5930__A1 _5926_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3571_ _3571_/A _3571_/B _3571_/C VGND VGND VPWR VPWR _3571_/X sky130_fd_sc_hd__or3_1
XANTENNA__3816__D _3816_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5310_ _5310_/A VGND VGND VPWR VPWR _6070_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3941__B1 _3940_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5241_ _4610_/X _5048_/X _4618_/X _4824_/X VGND VGND VPWR VPWR _5241_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5694__B1 _5692_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4497__A1 _4859_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5172_ _5973_/B _5171_/X _4420_/X VGND VGND VPWR VPWR _5172_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4123_ _3773_/C _3571_/B _3954_/X _3501_/Y VGND VGND VPWR VPWR _4123_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_110_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4054_ _4053_/X _3926_/X _3748_/A VGND VGND VPWR VPWR _4054_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4249__A1 _4520_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput2 EN_memory_dmem_response_get VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__buf_4
XANTENNA__5446__B1 _5439_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5997__A1 _5998_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3005_ _3005_/A VGND VGND VPWR VPWR _3005_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5749__A1 _4952_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5213__A3 _4815_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4960__A _4960_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4956_ _4956_/A _5971_/B _5944_/B _4956_/D VGND VGND VPWR VPWR _4956_/Y sky130_fd_sc_hd__nand4_4
X_4887_ _5188_/B VGND VGND VPWR VPWR _4887_/X sky130_fd_sc_hd__buf_2
X_3907_ _3904_/X _3464_/X _3711_/X _3906_/Y _4036_/A VGND VGND VPWR VPWR _3907_/Y
+ sky130_fd_sc_hd__a311oi_4
XANTENNA__3576__A _3934_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4972__A2 _4971_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3838_ _3838_/A VGND VGND VPWR VPWR _3838_/X sky130_fd_sc_hd__buf_2
XFILLER_20_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4724__A2 _4350_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5921__A1 _4665_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6102__D _6102_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3769_ _3766_/Y _3768_/Y _3492_/X VGND VGND VPWR VPWR _3769_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5791__A _6187_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5508_ _5508_/A VGND VGND VPWR VPWR _5531_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5439_ _5439_/A VGND VGND VPWR VPWR _5439_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5685__B1 _4665_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6138__CLK _6146_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3696__C1 _3695_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4645__D1 _4644_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4660__A1 _5188_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3463__A2 _4042_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3999__B1 _3633_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5031__A _5140_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4255__A4 _4245_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5452__A3 _5701_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4870__A _5018_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4963__A2 _4959_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3486__A _3871_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5912__A1 _4672_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5373__C1 _5369_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3923__B1 _3495_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5979__B2 _4898_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5979__A1 _5061_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4100__B1 _3900_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3454__A2 _3452_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4810_ _5188_/D VGND VGND VPWR VPWR _4843_/A sky130_fd_sc_hd__buf_2
XANTENNA__4780__A _4780_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5790_ _6186_/Q _5646_/X _5774_/Y _5789_/Y VGND VGND VPWR VPWR _6186_/D sky130_fd_sc_hd__a2bb2oi_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _4738_/A _4729_/B _5016_/A _4604_/A VGND VGND VPWR VPWR _4931_/A sky130_fd_sc_hd__o211ai_4
XANTENNA__4954__A2 _4668_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3396__A _3806_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4672_ _4672_/A VGND VGND VPWR VPWR _4672_/X sky130_fd_sc_hd__buf_4
XFILLER_119_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3623_ _3959_/D _3623_/B _3623_/C _3622_/X VGND VGND VPWR VPWR _3623_/X sky130_fd_sc_hd__or4b_1
XANTENNA__3914__B1 _4073_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4004__B _4004_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3554_ _3549_/X _3767_/D _3499_/X _3910_/A _3553_/X VGND VGND VPWR VPWR _3554_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5116__C1 _5115_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5761__D _5761_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3485_ _3873_/B VGND VGND VPWR VPWR _3871_/B sky130_fd_sc_hd__buf_4
X_5224_ input32/X _4978_/X _5223_/X VGND VGND VPWR VPWR _5224_/Y sky130_fd_sc_hd__a21oi_2
X_5155_ _5140_/D _5153_/Y _5152_/Y _4582_/X _4794_/X VGND VGND VPWR VPWR _5155_/Y
+ sky130_fd_sc_hd__a41oi_1
XANTENNA__4955__A _4955_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5682__A3 _5681_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3693__A2 _3673_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5419__B1 _5528_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4106_ _3572_/A _3797_/A _3911_/C _3157_/C _3932_/B VGND VGND VPWR VPWR _4106_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_56_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5086_ _6054_/Q _5040_/X _5047_/X _5085_/Y VGND VGND VPWR VPWR _6054_/D sky130_fd_sc_hd__a2bb2oi_1
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4037_ _3475_/D _3205_/X _3882_/B _3902_/A _3673_/A VGND VGND VPWR VPWR _4037_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3070__S _3072_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3445__A2 _3444_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5198__A2 _5197_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_13_0_CLK clkbuf_3_6_0_CLK/X VGND VGND VPWR VPWR _6196_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_40_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5988_ _5988_/A _5988_/B VGND VGND VPWR VPWR _5989_/A sky130_fd_sc_hd__or2_1
X_4939_ _4680_/X _4935_/X _4750_/Y VGND VGND VPWR VPWR _4939_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4158__B1 _3628_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5370__A2 _5369_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3920__A3 _3359_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5658__B1 _4665_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4287__D _4405_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4881__A1 _4870_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4865__A _4865_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3684__A2 _3683_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5830__B1 _5237_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4094__C1 _3414_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4633__A1 _6127_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5189__A2 _4378_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4105__A _4105_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5897__B1 _4387_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4759__B _4860_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4164__A3 _3290_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3663__B _3711_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output89_A _3082_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3382__C _3779_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3270_ _4074_/C VGND VGND VPWR VPWR _3271_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5649__B1 _5403_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5113__A2 _5105_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5664__A3 _4961_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3675__A2 _3593_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2994__S _2998_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5102__C _5102_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5911_ _5712_/A _5102_/D _4610_/X _5782_/X VGND VGND VPWR VPWR _5911_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5821__B1 _5905_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5842_ _5018_/C _5098_/X _4740_/X _5029_/X _4948_/A VGND VGND VPWR VPWR _5842_/X
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__4388__B1 _4387_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5773_ _6114_/Q _4721_/X _5772_/X VGND VGND VPWR VPWR _5773_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4724_ _4692_/A _4350_/A _4707_/C _5048_/A VGND VGND VPWR VPWR _4726_/A sky130_fd_sc_hd__a31o_4
X_2985_ _5382_/B _6060_/Q VGND VGND VPWR VPWR _2986_/C sky130_fd_sc_hd__or2b_1
XANTENNA__3060__A0 _6190_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4655_ _4333_/A _5818_/S _5061_/A _4835_/A VGND VGND VPWR VPWR _4656_/A sky130_fd_sc_hd__a211o_1
Xclkbuf_3_2_0_CLK clkbuf_3_3_0_CLK/A VGND VGND VPWR VPWR clkbuf_4_5_0_CLK/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5888__B1 _5020_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3606_ _3606_/A VGND VGND VPWR VPWR _3781_/C sky130_fd_sc_hd__clkbuf_2
X_4586_ _4879_/A VGND VGND VPWR VPWR _4666_/A sky130_fd_sc_hd__buf_2
XANTENNA__4155__A3 _4152_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3899__C1 _3838_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput82 memory_imem_request_put[8] VGND VGND VPWR VPWR _3353_/A sky130_fd_sc_hd__buf_2
Xinput60 memory_dmem_request_put[86] VGND VGND VPWR VPWR _4174_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__5772__C _5772_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput71 memory_dmem_request_put[97] VGND VGND VPWR VPWR _4219_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__3363__A1 _3847_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3363__B2 _3362_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3537_ _3537_/A _3537_/B _3491_/A VGND VGND VPWR VPWR _3537_/X sky130_fd_sc_hd__or3b_4
XFILLER_107_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3468_ _3468_/A _3468_/B _3621_/A VGND VGND VPWR VPWR _3468_/X sky130_fd_sc_hd__and3_1
XANTENNA__5104__A2 _5102_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4863__A1 _5745_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3399_ _3841_/B _3847_/A _3653_/A VGND VGND VPWR VPWR _3807_/A sky130_fd_sc_hd__o21ai_4
X_5207_ _5148_/C _4409_/X _5018_/D _4345_/A VGND VGND VPWR VPWR _5207_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4312__B1 _6138_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4685__A _4685_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6187_ _6204_/CLK _6187_/D VGND VGND VPWR VPWR _6187_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4863__B2 _5079_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5138_ _4403_/X _5102_/C _4574_/X _5732_/B _5137_/X VGND VGND VPWR VPWR _5138_/Y
+ sky130_fd_sc_hd__o311ai_4
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4615__A1 _4329_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5069_ _4931_/X _4871_/Y _5068_/X _4387_/X VGND VGND VPWR VPWR _5069_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5812__B1 _4657_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4091__A2 _3834_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3748__B _3748_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3467__C _4074_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3764__A _3938_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5879__B1 _5878_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input40_A memory_dmem_request_put[66] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4606__A1 _4600_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5803__B1 _5716_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output127_A _3029_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4082__A2 _4124_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4480__D _4960_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4790__B1 _4785_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5365__S _5365_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4440_ _4754_/A _4942_/A _4551_/A _5211_/A VGND VGND VPWR VPWR _4440_/Y sky130_fd_sc_hd__nand4_4
XANTENNA__3674__A _3767_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5876__A2_N _4715_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4542__B1 _4541_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5885__A3 _5883_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3896__A2 _3457_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4371_ _4307_/A _4362_/A _4308_/X _4309_/X _4364_/A VGND VGND VPWR VPWR _4415_/A
+ sky130_fd_sc_hd__o41ai_1
X_6110_ _6204_/CLK _6110_/D VGND VGND VPWR VPWR _6110_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6200__D _6200_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3322_ _3589_/B VGND VGND VPWR VPWR _3992_/A sky130_fd_sc_hd__buf_2
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3253_ _3858_/A VGND VGND VPWR VPWR _3847_/A sky130_fd_sc_hd__buf_2
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6202_/CLK _6041_/D VGND VGND VPWR VPWR _6041_/Q sky130_fd_sc_hd__dfxtp_1
X_3184_ _3443_/B VGND VGND VPWR VPWR _3440_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4845__A1 _4614_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4952__B _4952_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5767__C _5767_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5825_ _4829_/Y _4316_/X _5823_/X _5824_/Y _4875_/X VGND VGND VPWR VPWR _5825_/Y
+ sky130_fd_sc_hd__a32oi_4
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3820__A2 _3457_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5756_ _5756_/A VGND VGND VPWR VPWR _5756_/X sky130_fd_sc_hd__buf_2
XFILLER_22_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5687_ _5687_/A _5687_/B _5687_/C VGND VGND VPWR VPWR _5687_/X sky130_fd_sc_hd__and3_1
X_4707_ _4865_/D _4862_/A _4707_/C _4707_/D VGND VGND VPWR VPWR _4708_/D sky130_fd_sc_hd__nand4_1
XANTENNA__4781__B1 _5006_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3584__A1 _4124_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4638_ _4759_/A VGND VGND VPWR VPWR _4929_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_108_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3887__A2 _3883_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4569_ _4746_/A _4563_/X _5755_/A _4956_/A _4568_/X VGND VGND VPWR VPWR _4569_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_1_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6110__D _6110_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5089__A1 _5256_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3639__A2 _3635_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4064__A2 _4060_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3759__A _4002_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5261__B2 input20/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5261__A1 input12/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5677__C _5677_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4581__C _4581_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3811__A2 _3810_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5013__A1 _6146_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3909__D _3909_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5564__A2 _5968_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3024__A0 _6030_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3575__B2 _3520_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3575__A1 _3910_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4102__B _4102_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3878__A2 _3874_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6020__D _6020_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3660__C _4092_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5252__A1 _4765_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3940_ _3936_/X _3699_/A _3937_/X _3939_/X VGND VGND VPWR VPWR _3940_/X sky130_fd_sc_hd__a31o_2
XANTENNA__4055__A2 _4049_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3388__B _3802_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3871_ _3871_/A _3871_/B _3904_/D VGND VGND VPWR VPWR _3871_/X sky130_fd_sc_hd__or3_1
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5555__A2 _5640_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3015__A0 _6026_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5610_ _6164_/Q _6032_/Q _5616_/S VGND VGND VPWR VPWR _5611_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4763__B1 _4757_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5541_ _5541_/A VGND VGND VPWR VPWR _6138_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3608__S _4042_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5472_ _5444_/X _5433_/X _5470_/X _5540_/A _5471_/X VGND VGND VPWR VPWR _6116_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_99_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4423_ _4699_/A VGND VGND VPWR VPWR _4423_/X sky130_fd_sc_hd__buf_4
XANTENNA__3869__A2 _3910_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6021__CLK _6155_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4354_ _4354_/A _4354_/B _4358_/A _4354_/D VGND VGND VPWR VPWR _4729_/B sky130_fd_sc_hd__nand4_4
XFILLER_113_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3305_ _3305_/A _3343_/A _3475_/D VGND VGND VPWR VPWR _3305_/X sky130_fd_sc_hd__or3b_1
XANTENNA__5124__A _5124_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_86_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4818__A1 _5140_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4285_ _4301_/A _4285_/B _4301_/C _4405_/D VGND VGND VPWR VPWR _4298_/A sky130_fd_sc_hd__nand4_4
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6171__CLK _6203_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6024_ _6045_/CLK _6024_/D VGND VGND VPWR VPWR _6024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3236_ _3446_/B VGND VGND VPWR VPWR _3983_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__4294__A2 _4293_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3167_ _3437_/A VGND VGND VPWR VPWR _3632_/A sky130_fd_sc_hd__buf_2
X_3098_ _3098_/A VGND VGND VPWR VPWR _3098_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5243__A1 _4855_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5243__B2 _5829_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4046__A2 _4041_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4451__C1 _4450_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5546__A2 _5715_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5808_ _5791_/Y _5166_/A _5804_/Y _5807_/Y VGND VGND VPWR VPWR _6187_/D sky130_fd_sc_hd__a22oi_1
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3006__A0 _6022_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6105__D _6105_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5739_ _4665_/A _5737_/Y _5738_/Y _4793_/X VGND VGND VPWR VPWR _5739_/Y sky130_fd_sc_hd__a2bb2oi_2
XFILLER_10_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5944__D _5944_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4203__A input1/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5018__B _5018_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5849__A3 _4630_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5034__A _5971_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4809__A1 _4801_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4809__B2 _4189_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4873__A _4873_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5234__A1 _5018_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5234__B2 _5829_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4037__A2 _3205_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3489__A _3648_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5785__A2 _4935_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4993__B1 _4992_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3796__B2 _3728_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3796__A1 _3792_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4745__B1 _4743_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6044__CLK _6202_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6194__CLK _6196_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4070_ _3967_/X _3975_/B _3962_/A _3648_/Y _3230_/X VGND VGND VPWR VPWR _4070_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4783__A _4864_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3021_ _6029_/Q _6161_/Q _3021_/S VGND VGND VPWR VPWR _3022_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5473__B2 _6117_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4028__A2 _4042_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5225__A1 _5201_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5776__A2 _5775_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4972_ _4524_/X _4971_/X _4456_/X _5125_/A VGND VGND VPWR VPWR _4973_/B sky130_fd_sc_hd__o31a_1
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3923_ _4004_/C _3543_/B _3495_/X VGND VGND VPWR VPWR _3923_/Y sky130_fd_sc_hd__o21ai_4
X_3854_ _3701_/X _3241_/X _3848_/X _3853_/X VGND VGND VPWR VPWR _3854_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5818__S _5818_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4736__B1 _4621_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3539__A1 _3535_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5933__C1 _4957_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3785_ _3139_/X _3577_/X _4116_/A _3784_/Y VGND VGND VPWR VPWR _3785_/X sky130_fd_sc_hd__a31o_1
XFILLER_118_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5524_ _5523_/X _4287_/B _5498_/X _5491_/X _6133_/Q VGND VGND VPWR VPWR _5525_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_105_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5455_ input20/X _5437_/X _5439_/X input12/X VGND VGND VPWR VPWR _5455_/X sky130_fd_sc_hd__a22o_1
X_4406_ _4860_/A VGND VGND VPWR VPWR _4926_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3862__A _3862_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5161__B1 _5042_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5386_ _5383_/X _5386_/B _6014_/B VGND VGND VPWR VPWR _5387_/A sky130_fd_sc_hd__and3b_1
XFILLER_113_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4337_ _5067_/A VGND VGND VPWR VPWR _4742_/A sky130_fd_sc_hd__buf_2
XFILLER_59_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5059__A4 _4563_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4268_ _4268_/A _4268_/B VGND VGND VPWR VPWR _4268_/Y sky130_fd_sc_hd__nor2_2
XFILLER_101_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4693__A _5188_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3219_ _3387_/B VGND VGND VPWR VPWR _3461_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5004__D _5004_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6007_ _5291_/X _5294_/X _6013_/C _5410_/X VGND VGND VPWR VPWR _6204_/D sky130_fd_sc_hd__o31a_1
XANTENNA__5464__B2 _5260_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5464__A1 _6114_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6008__A3 _5367_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4199_ _4717_/A _4718_/A _4804_/A VGND VGND VPWR VPWR _4199_/X sky130_fd_sc_hd__or3_2
XANTENNA__5216__A1 _5006_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4019__A2 _3835_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3490__A3 _3359_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3102__A _3102_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6067__CLK _6074_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5955__C _5955_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3756__B _3799_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5029__A _5029_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3475__C _3871_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5971__B _5971_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3950__A1 _3948_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3772__A _3781_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5690__C _5690_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5455__B2 input12/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5455__A1 input20/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3466__B1 _3241_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4663__C1 _5756_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5207__A1 _5148_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5758__A2 _4423_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3012__A _3056_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4966__B1 _4965_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3769__A1 _3766_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4430__A2 _4926_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5638__S _5638_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5915__C1 _5914_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3570_ _3592_/A _3956_/B _3600_/A VGND VGND VPWR VPWR _3571_/B sky130_fd_sc_hd__o21a_4
XANTENNA__5930__A2 _5927_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5391__B1 _4225_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4778__A _4778_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3941__A1 _3562_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5240_ _5240_/A _5240_/B _5240_/C _5240_/D VGND VGND VPWR VPWR _5240_/X sky130_fd_sc_hd__or4_2
XANTENNA__5143__B1 _4420_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5694__A1 _4858_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4497__A2 _5715_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5171_ _5170_/X _5971_/D _5018_/B _4661_/X _5029_/X VGND VGND VPWR VPWR _5171_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5694__B2 _5693_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5291__A_N input2/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4859__A_N _5757_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4122_ _3357_/X _6043_/Q _4121_/X _3453_/X VGND VGND VPWR VPWR _6043_/D sky130_fd_sc_hd__a22o_1
XFILLER_96_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4053_ _3910_/C _3362_/Y _3571_/B _3588_/X VGND VGND VPWR VPWR _4053_/X sky130_fd_sc_hd__a31o_1
XFILLER_56_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4249__A2 _4859_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5446__A1 input18/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5446__B2 input10/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5402__A _5402_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5997__A2 _5998_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput3 EN_memory_imem_request_put VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_2
X_3004_ _6021_/Q _6153_/Q _3010_/S VGND VGND VPWR VPWR _3005_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5749__A2 _5736_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4955_ _4955_/A VGND VGND VPWR VPWR _5944_/B sky130_fd_sc_hd__buf_4
XFILLER_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3906_ _3666_/A _3567_/X _3205_/X _4152_/B _4105_/A VGND VGND VPWR VPWR _3906_/Y
+ sky130_fd_sc_hd__a221oi_2
X_4886_ _4672_/X _4332_/X _4882_/X _4885_/Y VGND VGND VPWR VPWR _4886_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__3576__B _3576_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4972__A3 _4456_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4709__B1 _4708_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3837_ _3830_/X _3517_/X _3833_/X _4124_/C _3836_/X VGND VGND VPWR VPWR _3837_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__5906__C1 _5403_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3068__S _3072_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4724__A3 _4707_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5921__A2 _4956_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3768_ _3674_/X _3748_/C _3767_/X _3695_/A VGND VGND VPWR VPWR _3768_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_118_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4688__A _4869_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3393__C1 _3692_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5507_ _5495_/X _4632_/X _5498_/X _6127_/Q _5499_/X VGND VGND VPWR VPWR _5509_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_106_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3592__A _3592_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3699_ _3699_/A VGND VGND VPWR VPWR _3699_/X sky130_fd_sc_hd__buf_6
XFILLER_10_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5685__A1 _5026_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5438_ _5392_/C _4227_/A _5438_/C _5438_/D VGND VGND VPWR VPWR _5439_/A sky130_fd_sc_hd__and4bb_2
XFILLER_121_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3696__B1 _3539_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5369_ _4520_/A _4859_/B _4859_/C _5367_/Y _6143_/Q VGND VGND VPWR VPWR _5369_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__4200__B _4200_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4645__C1 _4642_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5842__D1 _4948_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3448__B1 _3571_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5312__A _5312_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3999__A1 _3998_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3999__B2 _3708_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4660__A2 _4929_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5070__C1 _5152_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4963__A3 _4891_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5982__A _5982_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5373__B1 _5381_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3923__A1 _4004_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5912__A2 _5167_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input70_A memory_dmem_request_put[96] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4598__A _4832_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3007__A _3007_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3439__B1 _3438_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4100__A1 _3653_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5979__A2 _5062_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5222__A _5643_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3454__A3 _3453_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4939__B1 _4750_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4954__A3 _4852_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4740_ _4707_/D _4350_/A _4707_/C _4697_/A VGND VGND VPWR VPWR _4740_/X sky130_fd_sc_hd__a31o_4
XFILLER_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4671_ _5003_/C VGND VGND VPWR VPWR _4671_/X sky130_fd_sc_hd__buf_2
XANTENNA__3396__B _3396_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3622_ _3157_/X _3621_/X _3281_/A VGND VGND VPWR VPWR _3622_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6203__D _6203_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3914__A1 _3780_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4004__C _4004_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3553_ _3553_/A VGND VGND VPWR VPWR _3553_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5116__B1 _4742_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4301__A _4301_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3484_ _3871_/A VGND VGND VPWR VPWR _3536_/A sky130_fd_sc_hd__buf_2
XANTENNA__3678__B1 _6022_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5223_ _4716_/A _4513_/A _5431_/A _5042_/A VGND VGND VPWR VPWR _5223_/X sky130_fd_sc_hd__o211a_1
X_5154_ _5018_/C _4840_/X _5152_/Y _5153_/Y VGND VGND VPWR VPWR _5154_/X sky130_fd_sc_hd__o211a_1
XFILLER_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4105_ _4105_/A _4105_/B _4105_/C VGND VGND VPWR VPWR _4105_/X sky130_fd_sc_hd__or3_1
XFILLER_57_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5419__A1 _5416_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5085_ _5057_/Y _5059_/X _5220_/C _5084_/Y VGND VGND VPWR VPWR _5085_/Y sky130_fd_sc_hd__o211ai_4
XANTENNA__4627__C1 _4626_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4036_ _4036_/A _4036_/B _4036_/C _4036_/D VGND VGND VPWR VPWR _4036_/X sky130_fd_sc_hd__or4_1
XFILLER_37_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3850__B1 _3849_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5047__A1_N _5041_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5052__C1 _4665_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5987_ _5984_/Y _5985_/Y _5986_/Y _5570_/X _5998_/C VGND VGND VPWR VPWR _5988_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4938_ _4398_/X _4935_/X _5712_/C _4937_/Y VGND VGND VPWR VPWR _4938_/X sky130_fd_sc_hd__o211a_1
X_4869_ _4869_/A VGND VGND VPWR VPWR _5018_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__4158__A1 _3558_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5355__A0 _6048_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6113__D _6113_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6105__CLK _6145_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5307__A _5307_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4211__A _4211_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5658__A1 _4783_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3920__A4 _3919_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3669__B1 _4092_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4881__A2 _4871_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4865__B _5048_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5042__A _5042_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4094__B1 _3868_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5830__A1 _4875_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5189__A3 _5706_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5594__A0 _6157_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4105__B _4105_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6023__D _6023_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5346__A0 _6180_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5897__A1 _5896_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4759__C _4759_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3663__C _3663_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3382__D _3382_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5649__A1 _5045_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__A3 _5108_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3675__A3 _3674_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3465__A1_N _3457_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4609__C1 _4364_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5910_ _5020_/X _4378_/Y _4852_/Y _4744_/X VGND VGND VPWR VPWR _5910_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4085__B1 _3649_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5821__A1 _6101_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5282__C1 _5279_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5102__D _5102_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3798__B1_N _4105_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5841_ _6189_/Q _4629_/X _4630_/X _5822_/X _5840_/X VGND VGND VPWR VPWR _6189_/D
+ sky130_fd_sc_hd__o32a_1
XANTENNA__4388__A1 _4374_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5772_ _5772_/A _5772_/B _5772_/C VGND VGND VPWR VPWR _5772_/X sky130_fd_sc_hd__and3_1
XANTENNA__6128__CLK _6147_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2984_ _5381_/B VGND VGND VPWR VPWR _5382_/B sky130_fd_sc_hd__clkbuf_2
X_4723_ _4720_/X _4721_/X _4189_/A _4722_/Y VGND VGND VPWR VPWR _4723_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3060__A1 _6066_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5337__A0 _6055_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5888__A1 _5211_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4654_ _4654_/A VGND VGND VPWR VPWR _5757_/B sky130_fd_sc_hd__buf_2
XFILLER_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4585_ _4585_/A VGND VGND VPWR VPWR _4879_/A sky130_fd_sc_hd__buf_2
X_3605_ _3496_/Y _3601_/X _3308_/A _3604_/X _3281_/A VGND VGND VPWR VPWR _3613_/A
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3899__B1 _3898_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput50 memory_dmem_request_put[76] VGND VGND VPWR VPWR _4654_/A sky130_fd_sc_hd__clkbuf_4
Xinput61 memory_dmem_request_put[87] VGND VGND VPWR VPWR _4174_/A sky130_fd_sc_hd__clkbuf_1
Xinput72 memory_dmem_request_put[98] VGND VGND VPWR VPWR _4169_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__5127__A _5127_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3363__A2 _3557_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3536_ _3536_/A VGND VGND VPWR VPWR _3536_/X sky130_fd_sc_hd__clkbuf_4
Xinput83 memory_imem_request_put[9] VGND VGND VPWR VPWR _3301_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5104__A3 _5103_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3870__A _3870_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3467_ _4065_/A _4042_/D _4074_/C VGND VGND VPWR VPWR _3476_/A sky130_fd_sc_hd__and3_1
XANTENNA__4312__A1 _4482_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5206_ _4629_/A _4630_/A _5204_/X _5205_/Y VGND VGND VPWR VPWR _5206_/X sky130_fd_sc_hd__o22a_1
X_3398_ _3657_/C VGND VGND VPWR VPWR _3653_/A sky130_fd_sc_hd__buf_2
XFILLER_69_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6186_ _6204_/CLK _6186_/D VGND VGND VPWR VPWR _6186_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4863__A2 _5034_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5137_ _4702_/A _4891_/A _4693_/X _5721_/C VGND VGND VPWR VPWR _5137_/X sky130_fd_sc_hd__a211o_1
XFILLER_57_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3195__C_N _3194_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3081__S _3083_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5068_ _5152_/D VGND VGND VPWR VPWR _5068_/X sky130_fd_sc_hd__buf_2
XANTENNA__4615__A2 _4330_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5812__A1 _5097_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4019_ _3183_/X _3835_/X _3520_/X _4135_/A VGND VGND VPWR VPWR _4019_/X sky130_fd_sc_hd__o22a_1
XFILLER_44_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4076__B1 _3838_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6108__D _6108_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3823__B1 _6030_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4206__A _4283_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3748__C _3748_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5328__A0 _6187_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5879__A1 _5877_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4000__B1 _3999_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4876__A _4876_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3780__A _3780_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5500__B1 _6125_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input33_A memory_dmem_request_put[59] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4606__A2 _4605_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5803__B2 _5802_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5803__A1 _5715_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6018__D _6018_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4082__A3 _3249_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4116__A _4116_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5567__B1 _5499_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3578__C1 _3577_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3020__A _3020_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4775__D1 _4673_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4790__A1 _4680_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3674__B _3674_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4542__A1 _4532_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4370_ _4362_/X _5263_/A _4364_/X _4369_/Y VGND VGND VPWR VPWR _4370_/X sky130_fd_sc_hd__o211a_2
X_3321_ _3754_/B VGND VGND VPWR VPWR _3589_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4786__A _5061_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3252_ _3956_/A _3687_/A VGND VGND VPWR VPWR _3998_/C sky130_fd_sc_hd__nand2_4
Xclkbuf_4_12_0_CLK clkbuf_3_6_0_CLK/X VGND VGND VPWR VPWR _6205_/CLK sky130_fd_sc_hd__clkbuf_2
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _6202_/CLK _6040_/D VGND VGND VPWR VPWR _6040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4845__A2 _4738_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3183_ _4004_/C VGND VGND VPWR VPWR _3183_/X sky130_fd_sc_hd__clkbuf_4
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4058__B1 _3546_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3805__B1 _3804_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4952__C _4952_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5410__A _5422_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5007__C1 _5006_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5824_ _4960_/X _4840_/X _5971_/C _4855_/Y VGND VGND VPWR VPWR _5824_/Y sky130_fd_sc_hd__o31ai_2
XFILLER_62_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3820__A3 _3762_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5755_ _5755_/A _5755_/B _5755_/C _5755_/D VGND VGND VPWR VPWR _5755_/X sky130_fd_sc_hd__or4_2
X_4706_ _4772_/A VGND VGND VPWR VPWR _4707_/C sky130_fd_sc_hd__buf_2
XANTENNA__4781__A1 _5829_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5686_ _5706_/A _5706_/B _5706_/C _4656_/A VGND VGND VPWR VPWR _5746_/A sky130_fd_sc_hd__a31o_1
XANTENNA__3584__A2 _3525_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5983__A2_N _5982_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4637_ _5191_/A VGND VGND VPWR VPWR _4855_/D sky130_fd_sc_hd__buf_2
XANTENNA__5730__B1 _4657_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4568_ _4767_/A VGND VGND VPWR VPWR _4568_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4696__A _4696_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3519_ _4092_/B VGND VGND VPWR VPWR _3519_/X sky130_fd_sc_hd__buf_2
X_4499_ _5079_/A _4456_/X _4495_/Y _4498_/X VGND VGND VPWR VPWR _4504_/B sky130_fd_sc_hd__o211ai_1
XANTENNA__5089__A2 _5757_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3639__A3 _3637_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6169_ _6197_/CLK _6169_/D VGND VGND VPWR VPWR _6169_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4049__B1 _4048_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5797__B1 _5796_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3759__B _3759_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5261__A2 _4717_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4581__D _5078_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5549__B1 _5499_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3811__A3 _3727_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5564__A3 _4990_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3024__A1 _6162_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3575__A2 _3519_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3980__C1 _3979_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4102__C _4102_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3660__D _4152_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_1_0_CLK clkbuf_3_1_0_CLK/A VGND VGND VPWR VPWR clkbuf_4_3_0_CLK/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5788__B1 _4498_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5252__A2 _5249_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4055__A3 _4051_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4460__B1 _4734_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3870_ _3870_/A _3870_/B VGND VGND VPWR VPWR _3904_/D sky130_fd_sc_hd__nor2_4
XFILLER_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3685__A _3959_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3015__A1 _6158_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4763__B2 _4762_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4763__A1 _4755_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3365__B_N _3272_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5960__B1 _5782_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5540_ _5540_/A _5540_/B VGND VGND VPWR VPWR _5541_/A sky130_fd_sc_hd__or2_1
XANTENNA__3971__C1 _3970_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5471_ _6116_/Q _5222_/X _5256_/X _5260_/X VGND VGND VPWR VPWR _5471_/X sky130_fd_sc_hd__o22a_1
XFILLER_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4422_ _4422_/A VGND VGND VPWR VPWR _4422_/X sky130_fd_sc_hd__buf_4
XFILLER_98_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4353_ _4353_/A VGND VGND VPWR VPWR _4353_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3869__A3 _3773_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3304_ _3780_/C VGND VGND VPWR VPWR _3475_/D sky130_fd_sc_hd__clkbuf_2
X_4284_ _4293_/A _4246_/A _4308_/A _4246_/C _6135_/Q VGND VGND VPWR VPWR _4527_/A
+ sky130_fd_sc_hd__o41ai_4
XANTENNA__5405__A _5405_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5124__B _5124_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3235_ _3904_/A VGND VGND VPWR VPWR _3549_/A sky130_fd_sc_hd__buf_2
XANTENNA__4818__A2 _5976_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6023_ _6155_/CLK _6023_/D VGND VGND VPWR VPWR _6023_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3166_ _3461_/A VGND VGND VPWR VPWR _3437_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5779__B1 _4843_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3097_ _6054_/Q _6082_/Q _3105_/S VGND VGND VPWR VPWR _3098_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5243__A2 _5971_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5140__A _5140_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4451__B1 _4393_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3999_ _3998_/D _3572_/A _3911_/C _3633_/A _3708_/A VGND VGND VPWR VPWR _3999_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5546__A3 _4802_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5807_ _5676_/X _5806_/X _5769_/X VGND VGND VPWR VPWR _5807_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3006__A1 _6154_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5738_ _5903_/D _5170_/X _4385_/A _5680_/C VGND VGND VPWR VPWR _5738_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__5951__B1 _5721_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5669_ _5190_/X _5667_/X _4642_/X _5668_/X VGND VGND VPWR VPWR _5669_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__6121__D _6121_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5018__C _5018_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5703__B1 _5811_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3714__C1 _3713_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5034__B _5034_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4809__A2 _4802_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4690__B1 _4581_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5234__A2 _5755_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3489__B _4074_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5785__A3 _5097_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5985__A _5985_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4993__A1 input25/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3796__A2 _3795_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4745__A1 _5712_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5942__B1 _4773_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3953__C1 _3934_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6031__D _6031_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3020_ _3020_/A VGND VGND VPWR VPWR _3020_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4681__B1 _4605_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5225__A2 _5224_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4971_ _4297_/X _4536_/X _4404_/X _4405_/X VGND VGND VPWR VPWR _4971_/X sky130_fd_sc_hd__o2bb2a_4
XFILLER_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6206__D _6206_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3922_ _6034_/Q _3891_/X _3909_/X _3921_/Y VGND VGND VPWR VPWR _6034_/D sky130_fd_sc_hd__a211o_1
X_3853_ _3850_/X _3851_/Y _3680_/X _3852_/Y VGND VGND VPWR VPWR _3853_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4736__A1 _4369_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3539__A2 _3536_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5933__B1 _4771_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3784_ _3783_/X _3734_/Y _3695_/B VGND VGND VPWR VPWR _3784_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5523_ _5715_/A VGND VGND VPWR VPWR _5523_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5454_ _5454_/A VGND VGND VPWR VPWR _6111_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4405_ _4405_/A _4405_/B _4405_/C _4405_/D VGND VGND VPWR VPWR _4405_/X sky130_fd_sc_hd__and4_2
XANTENNA__5161__B2 input13/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5161__A1 input29/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5385_ _6098_/Q _5382_/B _5383_/B _5383_/C _5384_/Y VGND VGND VPWR VPWR _5386_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_87_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4336_ _4432_/A VGND VGND VPWR VPWR _5067_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5449__C1 _5448_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4267_ _4405_/B VGND VGND VPWR VPWR _4268_/B sky130_fd_sc_hd__inv_2
XANTENNA__4974__A _4974_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3218_ _3700_/A VGND VGND VPWR VPWR _3218_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4198_ _4515_/A VGND VGND VPWR VPWR _4804_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_6006_ _6206_/Q _5382_/B _5292_/Y VGND VGND VPWR VPWR _6013_/C sky130_fd_sc_hd__a21oi_2
XANTENNA__5464__A2 _5222_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3149_ _3165_/A VGND VGND VPWR VPWR _3443_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5216__A2 _4855_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3880__D1 _3879_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6116__D _6116_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3756__C _3756_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5955__D _5955_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4214__A _4243_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3475__D _3475_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3935__C1 _3577_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5971__C _5971_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3950__A2 _3868_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3772__B _3966_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5690__D _5690_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4360__C1 _4668_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5045__A _5045_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4884__A _4884_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3466__A1 _3178_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5455__A2 _5437_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5860__C1 _5123_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4663__B1 _4657_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5207__A2 _4409_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4966__A1 _4524_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3769__A2 _3768_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output102_A _3109_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6026__D _6026_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5122__A2_N _5119_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5915__B1 _5237_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4124__A _4124_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6161__CLK _6201_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5391__A1 _5438_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3941__A2 _3359_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5143__A1 _5097_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5694__A2 _4859_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4497__A3 _4518_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5170_ _5170_/A VGND VGND VPWR VPWR _5170_/X sky130_fd_sc_hd__buf_4
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4794__A _4819_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4121_ _3828_/X _4109_/X _4120_/X VGND VGND VPWR VPWR _4121_/X sky130_fd_sc_hd__a21bo_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4249__A3 _4859_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4052_ _3919_/X _3666_/X _3844_/X _3934_/B _3621_/C VGND VGND VPWR VPWR _4052_/Y
+ sky130_fd_sc_hd__a311oi_1
XANTENNA__5446__A2 _5437_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5851__C1 _4957_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5997__A3 _5998_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3003_ _3003_/A VGND VGND VPWR VPWR _3003_/X sky130_fd_sc_hd__clkbuf_1
Xinput4 EN_memory_imem_response_get VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3203__A _3344_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4331__A2_N _4527_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4954_ _4680_/A _4668_/B _4852_/C _4953_/X VGND VGND VPWR VPWR _4954_/X sky130_fd_sc_hd__a31o_2
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3905_ _4092_/D VGND VGND VPWR VPWR _4152_/B sky130_fd_sc_hd__buf_4
XFILLER_51_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4885_ _5878_/C _5118_/C _5079_/B _5240_/B VGND VGND VPWR VPWR _4885_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__4709__A1 _4702_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4034__A _4034_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3836_ _4135_/A _3834_/X _3835_/X _3347_/X _3975_/D VGND VGND VPWR VPWR _3836_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__5906__B1 _5529_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3767_ _3308_/A _3767_/B _3867_/A _3767_/D VGND VGND VPWR VPWR _3767_/X sky130_fd_sc_hd__and4b_1
XANTENNA__3917__C1 _3916_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3873__A _3983_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5921__A3 _5917_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3393__B1 _3392_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5506_ _6126_/Q _5504_/X _5388_/A _5505_/Y VGND VGND VPWR VPWR _6126_/D sky130_fd_sc_hd__a211o_1
XFILLER_106_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3698_ _3749_/B VGND VGND VPWR VPWR _3699_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5437_ _5437_/A VGND VGND VPWR VPWR _5437_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5685__A2 _5680_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3696__A1 _3580_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5368_ _6143_/Q _4211_/A _5367_/Y input2/X _4188_/A VGND VGND VPWR VPWR _5368_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_114_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4319_ _4482_/B _4234_/A _4318_/Y VGND VGND VPWR VPWR _4566_/A sky130_fd_sc_hd__o21ai_4
X_5299_ _5299_/A VGND VGND VPWR VPWR _6065_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4645__B1 _5004_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5842__C1 _5029_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3448__A1 _3338_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5200__A1_N _6057_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6034__CLK _6202_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3999__A2 _3572_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4209__A _4209_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3113__A _3113_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5070__B1 _4843_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3767__B _3767_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6184__CLK _6207_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4963__A4 _4961_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4879__A _4879_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3908__C1 _3907_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5982__B _5982_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5373__A1 _4238_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3923__A2 _3543_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input63_A memory_dmem_request_put[89] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5503__A _5503_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3439__A1 _4149_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4100__A2 _3293_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3023__A _3056_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4939__A1 _4680_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5691__A2_N _4571_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4670_ _4955_/A VGND VGND VPWR VPWR _5003_/C sky130_fd_sc_hd__clkbuf_4
X_3621_ _3621_/A _3679_/A _3621_/C _3621_/D VGND VGND VPWR VPWR _3621_/X sky130_fd_sc_hd__or4_2
X_3552_ _3956_/B _3500_/A _3600_/A VGND VGND VPWR VPWR _3553_/A sky130_fd_sc_hd__o21a_1
XANTENNA__3914__A2 _4092_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5116__A1 _4661_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4301__B _4405_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3483_ _3621_/C _3230_/X _3482_/X _3374_/X VGND VGND VPWR VPWR _3483_/Y sky130_fd_sc_hd__a211oi_1
XANTENNA__3127__A0 _6052_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3678__A1 _3665_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5222_ _5643_/B VGND VGND VPWR VPWR _5222_/X sky130_fd_sc_hd__clkbuf_2
X_5153_ _4855_/A _5034_/C _5240_/D _5240_/B _5152_/C VGND VGND VPWR VPWR _5153_/Y
+ sky130_fd_sc_hd__a32oi_4
XANTENNA__3678__B2 _3541_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6057__CLK _6203_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5419__A2 _5417_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4104_ _6042_/Q _3891_/X _4088_/X _4103_/X VGND VGND VPWR VPWR _6042_/D sky130_fd_sc_hd__a211o_1
XFILLER_111_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5084_ _5066_/X _5072_/Y _4393_/X _5083_/Y VGND VGND VPWR VPWR _5084_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__4627__B1 _4974_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4035_ _3350_/A _4061_/A _4035_/C VGND VGND VPWR VPWR _4036_/D sky130_fd_sc_hd__and3b_1
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3850__A1 _3525_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3868__A _3868_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5052__B1 _5020_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5986_ _6201_/Q _6198_/Q VGND VGND VPWR VPWR _5986_/Y sky130_fd_sc_hd__xnor2_1
X_4937_ _4937_/A _4937_/B _4999_/A _4937_/D VGND VGND VPWR VPWR _4937_/Y sky130_fd_sc_hd__nand4_4
XANTENNA__3602__A1 _3366_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3079__S _3083_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4868_ _4857_/Y _4867_/Y _4698_/X VGND VGND VPWR VPWR _4868_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4699__A _4699_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4158__A2 _3716_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3819_ _3818_/Y _3775_/Y _3492_/X VGND VGND VPWR VPWR _3819_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5355__A1 _6091_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4799_ _5646_/A VGND VGND VPWR VPWR _4799_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3669__A1 _3447_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5658__A2 _4398_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4866__B1 _5006_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4865__C _4865_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5323__A _5323_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4881__A3 _4874_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4094__A1 _3762_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5830__A2 _5018_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3778__A _3828_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5043__B1 _5042_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5594__A1 _6025_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4105__C _4105_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5346__A1 _6087_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5897__A2 _5068_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4554__C1 _4744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4402__A _5003_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3663__D _3938_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4306__C1 _4305_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3018__A _3018_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5649__A2 _5440_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4857__B1 _5732_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4609__B1 _4864_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4085__A1 _4084_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5821__A2 _4807_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5282__B1 _5272_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5840_ _4498_/X _5831_/Y _5982_/C _5839_/Y VGND VGND VPWR VPWR _5840_/X sky130_fd_sc_hd__o211a_1
XFILLER_22_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4388__A2 _4378_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5771_ _5751_/Y _5166_/A _5766_/Y _5770_/Y VGND VGND VPWR VPWR _6185_/D sky130_fd_sc_hd__a22oi_1
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2983_ input2/X VGND VGND VPWR VPWR _5381_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__3596__B1 _3724_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4722_ _6129_/Q _4975_/A _4224_/A VGND VGND VPWR VPWR _4722_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5337__A1 _6083_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4653_ _4648_/X _4581_/Y _4650_/X _4652_/X VGND VGND VPWR VPWR _4664_/B sky130_fd_sc_hd__a31o_1
XANTENNA__5408__A _5482_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput40 memory_dmem_request_put[66] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5888__A2 _5761_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4584_ _4584_/A VGND VGND VPWR VPWR _4584_/X sky130_fd_sc_hd__clkbuf_4
X_3604_ _3549_/A _4004_/B _3686_/A _3603_/X VGND VGND VPWR VPWR _3604_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3899__A1 _3546_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput51 memory_dmem_request_put[77] VGND VGND VPWR VPWR _5715_/B sky130_fd_sc_hd__clkbuf_4
Xinput62 memory_dmem_request_put[88] VGND VGND VPWR VPWR _4217_/D sky130_fd_sc_hd__clkbuf_1
Xinput73 memory_dmem_request_put[99] VGND VGND VPWR VPWR _4169_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__5127__B _5127_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3535_ _3830_/C _3533_/X _3534_/X _3830_/D VGND VGND VPWR VPWR _3535_/X sky130_fd_sc_hd__o22a_2
XFILLER_107_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3466_ _3178_/X _3157_/C _3241_/X _3465_/X VGND VGND VPWR VPWR _3466_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3870__B _3870_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4848__B1 _4568_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5205_ _6122_/Q _4807_/X _5013_/X VGND VGND VPWR VPWR _5205_/Y sky130_fd_sc_hd__o21ai_1
X_3397_ _3397_/A VGND VGND VPWR VPWR _3841_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_69_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4312__A2 _4308_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6185_ _6204_/CLK _6185_/D VGND VGND VPWR VPWR _6185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5136_ _5102_/A _4708_/A _5148_/B _5148_/A _5135_/Y VGND VGND VPWR VPWR _5136_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_57_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5067_ _5067_/A VGND VGND VPWR VPWR _5152_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__4076__A1 _4073_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5812__A2 _5944_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4018_ _3699_/X _4013_/X _4015_/Y _4017_/X _3580_/X VGND VGND VPWR VPWR _4018_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5273__B1 _5272_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3284__C1 _3283_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3823__A1 _3816_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3823__B2 _3822_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5025__B1 _5003_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3748__D _3748_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5969_ _6108_/Q _4807_/X _5905_/X VGND VGND VPWR VPWR _5969_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3587__B1 _3278_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4784__C1 _4364_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6124__D _6124_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5328__A1 _6079_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5318__A _5318_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4000__B2 _3962_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5879__A2 _4931_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4839__B1 _4697_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3780__B _4073_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5500__A1 _5495_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5500__B2 _5499_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5988__A _5988_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input26_A memory_dmem_request_put[52] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5803__A2 _4390_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3301__A _3301_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4116__B _4116_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5567__A1 _4199_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5567__B2 _6147_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4775__C1 _4259_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3578__B1 _3571_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6034__D _6034_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5228__A _5228_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4790__A2 _4783_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3674__C _3674_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4542__A2 _4539_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output94_A _3093_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3320_ _4089_/B _3814_/A _3319_/X VGND VGND VPWR VPWR _3320_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__3750__B1 _3816_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3251_ _3275_/B VGND VGND VPWR VPWR _3687_/A sky130_fd_sc_hd__buf_2
XFILLER_79_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4845__A3 _4772_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3182_ _3870_/B VGND VGND VPWR VPWR _4004_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_78_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3502__B1 _3428_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4058__A1 _3338_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5255__B1 _5227_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3266__C1 _3299_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3805__A1 _3934_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5007__B1 _4644_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4307__A _4307_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5823_ _4754_/X _5745_/B _5761_/D _5687_/A VGND VGND VPWR VPWR _5823_/X sky130_fd_sc_hd__a31o_1
XFILLER_34_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3569__B1 _3208_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5754_ _5752_/Y _5753_/X _4964_/A VGND VGND VPWR VPWR _5754_/Y sky130_fd_sc_hd__a21oi_4
X_4705_ _4705_/A VGND VGND VPWR VPWR _4772_/A sky130_fd_sc_hd__buf_2
XANTENNA__4781__A2 _4967_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5685_ _5026_/X _5680_/C _4779_/Y _4665_/A VGND VGND VPWR VPWR _5690_/A sky130_fd_sc_hd__a31o_1
XFILLER_118_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4636_ _4860_/C VGND VGND VPWR VPWR _5191_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__4042__A _4042_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5730__A1 _4398_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4977__A _5772_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4567_ _4929_/C _5744_/A _4580_/A VGND VGND VPWR VPWR _4956_/A sky130_fd_sc_hd__a21oi_4
XFILLER_89_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3741__B1 _3282_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3881__A _3881_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3518_ _4034_/B VGND VGND VPWR VPWR _4092_/B sky130_fd_sc_hd__clkbuf_2
X_4498_ _5125_/A VGND VGND VPWR VPWR _4498_/X sky130_fd_sc_hd__clkbuf_2
X_3449_ _3161_/A _3439_/X _3448_/Y _3815_/A VGND VGND VPWR VPWR _3449_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__3092__S _3094_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5089__A3 _5757_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6203_/CLK _6168_/D VGND VGND VPWR VPWR _6168_/Q sky130_fd_sc_hd__dfxtp_1
X_5119_ _5117_/Y _5118_/Y _4582_/X VGND VGND VPWR VPWR _5119_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6119__D _6119_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5246__B1 _5829_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4049__A1 _3347_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6099_ _6207_/CLK _6099_/D VGND VGND VPWR VPWR _6099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5797__A1 _5754_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3759__C _3816_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4217__A _4217_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5549__A1 _5523_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5549__B2 _6141_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5048__A _5048_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3980__B1 _3546_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4887__A _5188_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5485__B1 _5451_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6118__CLK _6147_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6029__D _6029_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output132_A _3038_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5788__A1 _5716_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4460__A1 _4860_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3031__A _3031_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3966__A _4042_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4763__A2 _5829_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5960__A1 _4750_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3971__B1 _3964_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5470_ input24/X _5437_/X _5439_/X _5431_/A VGND VGND VPWR VPWR _5470_/X sky130_fd_sc_hd__a22o_1
XFILLER_8_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5173__C1 _5140_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4421_ _4421_/A VGND VGND VPWR VPWR _4422_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__4797__A _4797_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4352_ _4832_/A VGND VGND VPWR VPWR _4353_/A sky130_fd_sc_hd__buf_4
XANTENNA__3723__B1 _3673_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3303_ _4073_/C VGND VGND VPWR VPWR _3305_/A sky130_fd_sc_hd__clkbuf_4
X_4283_ _4283_/A VGND VGND VPWR VPWR _4308_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3234_ _3582_/C VGND VGND VPWR VPWR _3904_/A sky130_fd_sc_hd__buf_2
XANTENNA__3206__A _3275_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4818__A3 _4456_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6022_ _6155_/CLK _6022_/D VGND VGND VPWR VPWR _6022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3165_ _3165_/A VGND VGND VPWR VPWR _3461_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_94_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5779__A1 _5078_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3096_ _3096_/A VGND VGND VPWR VPWR _3105_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__5243__A3 _4917_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5140__B _5140_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4451__A1 _4252_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3876__A _3876_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3998_ _3998_/A _4092_/B _3998_/C _3998_/D VGND VGND VPWR VPWR _3998_/X sky130_fd_sc_hd__or4_1
XFILLER_10_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5806_ _6115_/Q _5643_/A _5805_/X VGND VGND VPWR VPWR _5806_/X sky130_fd_sc_hd__a21o_1
XFILLER_22_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5737_ _4686_/X _4604_/X _4864_/Y _5018_/A VGND VGND VPWR VPWR _5737_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__5951__A1 _4459_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5951__B2 _4619_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5668_ _5078_/B _5687_/C _5003_/C _4887_/X _4827_/A VGND VGND VPWR VPWR _5668_/X
+ sky130_fd_sc_hd__a41o_1
X_4619_ _5188_/A _4619_/B _4852_/A VGND VGND VPWR VPWR _4619_/X sky130_fd_sc_hd__and3_4
XANTENNA__5018__D _5018_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5703__A1 _5676_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5599_ _6159_/Q _6027_/Q _5605_/S VGND VGND VPWR VPWR _5600_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5164__C1 _4984_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3714__B1 _3538_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4500__A _6142_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5034__C _5034_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5467__B1 _5451_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4809__A3 _4806_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4690__A1 _5745_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5219__B1 _4767_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3489__C _4135_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5985__B _5985_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4993__A2 _4978_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3796__A3 _3727_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3786__A _3786_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_4_11_0_CLK clkbuf_3_5_0_CLK/X VGND VGND VPWR VPWR _6147_/CLK sky130_fd_sc_hd__clkbuf_2
XANTENNA__4745__A2 _4737_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5942__A1 _5167_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3953__B1 _3338_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3705__B1 _3704_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5458__B1 _5439_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4681__A1 _4680_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4130__B1 _3700_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6090__CLK _6176_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4969__C1 _4836_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4970_ _4958_/Y _4963_/X _4964_/X _4969_/Y VGND VGND VPWR VPWR _4973_/A sky130_fd_sc_hd__o211ai_2
XFILLER_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5630__A0 _6173_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3921_ _3508_/X _3917_/X _3918_/X _3920_/Y VGND VGND VPWR VPWR _3921_/Y sky130_fd_sc_hd__a211oi_1
X_3852_ _4128_/A _3722_/X _3731_/D _3301_/A VGND VGND VPWR VPWR _3852_/Y sky130_fd_sc_hd__o31ai_1
XANTENNA__4736__A2 _4296_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5933__A1 _4360_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3539__A3 _3537_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3783_ _3157_/X _3780_/X _3782_/X _3537_/B VGND VGND VPWR VPWR _3783_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3944__B1 _5388_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5522_ _6132_/Q _5504_/X _5447_/X _5521_/Y VGND VGND VPWR VPWR _6132_/D sky130_fd_sc_hd__a211o_1
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5146__C1 _5145_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5453_ _5453_/A _5468_/B VGND VGND VPWR VPWR _5454_/A sky130_fd_sc_hd__and2_1
XANTENNA__4320__A _4566_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5697__B1 _5696_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4404_ _4482_/A _4308_/X _4309_/X _6134_/Q VGND VGND VPWR VPWR _4404_/X sky130_fd_sc_hd__o31a_2
XANTENNA__5161__A2 _4804_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5384_ _5373_/Y _5371_/Y _5376_/Y VGND VGND VPWR VPWR _5384_/Y sky130_fd_sc_hd__a21oi_1
X_4335_ _4307_/A _4362_/A _4246_/B _4309_/X _4364_/A VGND VGND VPWR VPWR _4432_/A
+ sky130_fd_sc_hd__o41a_2
XFILLER_5_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2981__A_N _6099_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5449__B1 _5447_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4266_ _4266_/A VGND VGND VPWR VPWR _4313_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__4974__B _4974_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3217_ _3621_/D VGND VGND VPWR VPWR _3700_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_39_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4197_ _4225_/A _4227_/A VGND VGND VPWR VPWR _4515_/A sky130_fd_sc_hd__nor2_1
X_6005_ _6203_/Q _5293_/X _6004_/Y VGND VGND VPWR VPWR _6203_/D sky130_fd_sc_hd__a21oi_1
X_3148_ _3446_/B VGND VGND VPWR VPWR _3278_/A sky130_fd_sc_hd__buf_2
XFILLER_55_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5216__A3 _5212_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3880__C1 _3866_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3079_ _6182_/Q _6074_/Q _3083_/S VGND VGND VPWR VPWR _3080_/A sky130_fd_sc_hd__mux2_2
XANTENNA__5621__A0 _6169_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5385__C1 _5384_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3935__B1 _3934_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6132__D _6132_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5971__D _5971_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5137__C1 _5721_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_3_0_0_CLK clkbuf_3_1_0_CLK/A VGND VGND VPWR VPWR clkbuf_4_1_0_CLK/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5688__B1 _5235_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4230__A _4230_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4360__B1 _4865_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4112__B1 _3648_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5860__B1 _4761_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3466__A2 _3157_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5061__A _5061_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4663__B2 _4662_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4663__A1 _5757_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5207__A3 _5018_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5612__A0 _6165_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4966__A2 _4431_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4405__A _4405_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5915__A1 _5910_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4124__B _4124_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6042__D _6042_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5391__A2 input7/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3941__A3 _3482_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5143__A2 _4459_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5679__B1 _5811_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4120_ _3707_/X _4115_/X _4117_/Y _4119_/X _3806_/A VGND VGND VPWR VPWR _4120_/X
+ sky130_fd_sc_hd__a221o_1
X_4051_ _3536_/A _3844_/X _3717_/X _4050_/X VGND VGND VPWR VPWR _4051_/X sky130_fd_sc_hd__o211a_1
XFILLER_110_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5851__B1 _5880_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput5 RST_N VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__buf_6
X_3002_ _6020_/Q _6152_/Q _3010_/S VGND VGND VPWR VPWR _3003_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5603__A0 _6161_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4953_ _5182_/A VGND VGND VPWR VPWR _4953_/X sky130_fd_sc_hd__buf_2
X_3904_ _3904_/A _3904_/B _3904_/C _3904_/D VGND VGND VPWR VPWR _3904_/X sky130_fd_sc_hd__or4_4
XANTENNA__3090__A0 _6187_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4884_ _4884_/A VGND VGND VPWR VPWR _5118_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_32_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4034__B _4034_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3835_ _3835_/A VGND VGND VPWR VPWR _3835_/X sky130_fd_sc_hd__buf_2
XANTENNA__4709__A2 _5152_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5906__A1 input12/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3917__B1 _4036_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3766_ _3764_/X _3634_/X _3765_/X _3815_/B VGND VGND VPWR VPWR _3766_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_20_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4590__B1 _5680_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3873__B _3873_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3393__A1 _3218_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5505_ _4522_/A _5433_/X _5504_/X VGND VGND VPWR VPWR _5505_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3697_ _3691_/X _3290_/X _3696_/Y _6023_/Q _3541_/X VGND VGND VPWR VPWR _6023_/D
+ sky130_fd_sc_hd__a32o_1
X_5436_ _5436_/A VGND VGND VPWR VPWR _5437_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_121_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4342__B1 _4341_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5685__A3 _4779_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4985__A _4985_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5367_ _6147_/Q _6146_/Q _6145_/Q _6144_/Q VGND VGND VPWR VPWR _5367_/Y sky130_fd_sc_hd__nor4_4
XANTENNA__3696__A2 _3596_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4318_ _4293_/A _4246_/A _4246_/B _4246_/C _6136_/Q VGND VGND VPWR VPWR _4318_/Y
+ sky130_fd_sc_hd__o41ai_4
X_5298_ _6189_/Q _6065_/Q _5306_/S VGND VGND VPWR VPWR _5299_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4249_ _4520_/A _4859_/B _4859_/C _6139_/Q VGND VGND VPWR VPWR _5756_/A sky130_fd_sc_hd__a31o_2
XFILLER_101_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4645__A1 _4612_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5842__B1 _4740_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3448__A2 _3571_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3999__A3 _3911_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6127__D _6127_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3605__C1 _3281_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5070__A1 _5096_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3767__C _3867_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3081__A0 _6183_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4225__A _4225_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4030__C1 _3562_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3908__B1 _3695_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5982__C _5982_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5373__A2 _5805_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3246__C_N _3746_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4895__A _4895_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input56_A memory_dmem_request_put[82] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3396__C_N _4002_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3439__A2 _3660_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4097__C1 _3470_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3304__A _3780_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5833__B1 _5761_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4100__A3 _3965_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6037__D _6037_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4939__A2 _4935_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4135__A _4135_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3072__A0 _6195_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3620_ _3781_/D _4034_/A VGND VGND VPWR VPWR _3679_/A sky130_fd_sc_hd__nor2_1
XANTENNA__4021__C1 _4020_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3551_ _3551_/A VGND VGND VPWR VPWR _3910_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3914__A3 _3382_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5116__A2 _4464_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3482_ _3482_/A VGND VGND VPWR VPWR _3482_/X sky130_fd_sc_hd__buf_2
XANTENNA__4301__C _4301_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3127__A1 _6096_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4324__B1 _4527_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3678__A2 _3290_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5221_ _6058_/Q _5040_/X _5206_/X _5220_/Y VGND VGND VPWR VPWR _6058_/D sky130_fd_sc_hd__a2bb2oi_1
X_5152_ _5152_/A _5152_/B _5152_/C _5152_/D VGND VGND VPWR VPWR _5152_/Y sky130_fd_sc_hd__nand4_2
XFILLER_69_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4103_ _3286_/X _4096_/X _4103_/C _4103_/D VGND VGND VPWR VPWR _4103_/X sky130_fd_sc_hd__and4bb_1
XFILLER_111_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5824__B1 _4855_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5083_ _5075_/Y _5077_/Y _4746_/A _5082_/Y VGND VGND VPWR VPWR _5083_/Y sky130_fd_sc_hd__o211ai_4
XANTENNA__3214__A _4034_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4627__A1 _4558_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4034_ _4034_/A _4034_/B _3397_/A VGND VGND VPWR VPWR _4061_/A sky130_fd_sc_hd__or3b_1
XFILLER_49_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3850__A2 _3631_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5052__B2 _5051_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5052__A1 _5049_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5985_ _5985_/A _5985_/B VGND VGND VPWR VPWR _5985_/Y sky130_fd_sc_hd__nand2_1
X_4936_ _4936_/A VGND VGND VPWR VPWR _4999_/A sky130_fd_sc_hd__buf_4
XANTENNA__3602__A2 _3432_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4867_ _4858_/Y _4859_/X _4863_/X _4866_/X VGND VGND VPWR VPWR _4867_/Y sky130_fd_sc_hd__o22ai_1
XANTENNA__5575__S _5583_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3884__A _3956_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4158__A3 _3868_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3818_ _3807_/X _3767_/X _3817_/Y _3695_/A VGND VGND VPWR VPWR _3818_/Y sky130_fd_sc_hd__o31ai_1
X_4798_ _4715_/X _6049_/Q _4723_/X _4797_/Y VGND VGND VPWR VPWR _6049_/D sky130_fd_sc_hd__a2bb2oi_1
X_3749_ _4044_/A _3749_/B _3749_/C _3749_/D VGND VGND VPWR VPWR _3749_/X sky130_fd_sc_hd__or4_1
XFILLER_21_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4315__B1 _4421_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5419_ _5416_/Y _5417_/Y _5528_/B VGND VGND VPWR VPWR _6104_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__5512__C1 _5511_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3669__A2 _3527_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4866__A1 _5829_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5604__A _5604_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4865__D _4865_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4079__C1 _4078_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5815__B1 _4393_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3124__A _3124_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4094__A2 _3254_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6151__CLK _6197_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3826__C1 _3787_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5830__A3 _5829_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3778__B _3792_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3054__A0 _6044_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5043__B2 input10/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5043__A1 input26/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4554__B1 _4551_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4003__C1 _3934_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5897__A3 _4773_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4306__B1 _4290_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4857__A1 _4581_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5514__A _5514_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4609__A1 _4243_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5806__B1 _5805_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3034__A _3056_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3817__C1 _3464_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4085__A2 _3208_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5282__A1 _5985_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4388__A3 _5102_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5770_ _5676_/X _5768_/X _5769_/X VGND VGND VPWR VPWR _5770_/Y sky130_fd_sc_hd__a21oi_1
X_2982_ _4186_/A VGND VGND VPWR VPWR _2986_/B sky130_fd_sc_hd__buf_2
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _5263_/A VGND VGND VPWR VPWR _4721_/X sky130_fd_sc_hd__buf_2
XANTENNA__3596__A1 _3593_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4652_ _4652_/A VGND VGND VPWR VPWR _4652_/X sky130_fd_sc_hd__buf_4
XFILLER_30_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3603_ _3603_/A _3603_/B _3612_/D _3603_/D VGND VGND VPWR VPWR _3603_/X sky130_fd_sc_hd__and4_4
Xinput30 memory_dmem_request_put[56] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5888__A3 _4839_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4583_ _4574_/X _4576_/X _4581_/Y _4582_/X VGND VGND VPWR VPWR _4583_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__3209__A _3754_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3899__A2 _3892_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput41 memory_dmem_request_put[67] VGND VGND VPWR VPWR _4200_/B sky130_fd_sc_hd__clkbuf_1
Xinput52 memory_dmem_request_put[78] VGND VGND VPWR VPWR _4218_/D sky130_fd_sc_hd__clkbuf_2
Xinput63 memory_dmem_request_put[89] VGND VGND VPWR VPWR _4217_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__6024__CLK _6045_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5127__C _5220_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3534_ _3756_/C VGND VGND VPWR VPWR _3534_/X sky130_fd_sc_hd__clkbuf_4
Xinput74 memory_imem_request_put[10] VGND VGND VPWR VPWR _3918_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3465_ _3457_/X _3674_/B _3463_/X _3464_/X VGND VGND VPWR VPWR _3465_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_6_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4848__A1 _4842_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6174__CLK _6201_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5204_ _5201_/X _5202_/Y _5968_/C _5260_/A VGND VGND VPWR VPWR _5204_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4312__A3 _4986_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3396_ _3806_/B _3396_/B _4002_/A VGND VGND VPWR VPWR _3396_/X sky130_fd_sc_hd__or3b_1
X_6184_ _6207_/CLK _6184_/D VGND VGND VPWR VPWR _6184_/Q sky130_fd_sc_hd__dfxtp_1
X_5135_ _5006_/A _4878_/Y _4852_/Y _5743_/B VGND VGND VPWR VPWR _5135_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_84_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5066_ _4422_/X _4423_/X _5060_/X _5065_/X VGND VGND VPWR VPWR _5066_/X sky130_fd_sc_hd__o22a_2
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5812__A3 _4671_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4017_ _3990_/X _4016_/X _3161_/X VGND VGND VPWR VPWR _4017_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4076__A2 _4075_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5273__A1 _5286_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3569__A2_N _3815_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3284__B1 _3674_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3823__A2 _3820_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5025__A1 _4707_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5968_ _5968_/A _5968_/B _5968_/C VGND VGND VPWR VPWR _5968_/X sky130_fd_sc_hd__and3_1
XFILLER_25_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4919_ _5745_/C _5078_/B _4675_/A _4744_/A VGND VGND VPWR VPWR _4919_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__3587__A1 _3956_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4784__B1 _4815_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5981__C1 _4767_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5899_ _5899_/A _5899_/B _5899_/C VGND VGND VPWR VPWR _5899_/X sky130_fd_sc_hd__or3_2
XANTENNA__4503__A _4503_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6140__D _6140_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4839__A1 _4754_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3780__C _3780_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5334__A _5334_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5500__A2 _4229_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5988__B _5988_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input19_A memory_dmem_request_put[45] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3909__B_N _3899_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5567__A2 _5433_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4775__B1 _4937_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3578__B2 _3576_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3578__A1 _4126_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5972__C1 _5971_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6047__CLK _6205_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5509__A _5509_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4413__A _4574_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4790__A3 _5761_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6050__D _6050_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3029__A _3029_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6197__CLK _6197_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3750__A1 _3537_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output87_A _2979_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3440_/A _3366_/A _3440_/B VGND VGND VPWR VPWR _3612_/D sky130_fd_sc_hd__nand3_4
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _3330_/A _3442_/B VGND VGND VPWR VPWR _3870_/B sky130_fd_sc_hd__or2b_4
XFILLER_78_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3502__A1 _4083_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3699__A _3699_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4058__A2 _3564_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5255__B2 _5254_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3266__B1 _4048_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3805__A2 _3798_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5007__A1 _4878_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5822_ _5822_/A _5822_/B VGND VGND VPWR VPWR _5822_/X sky130_fd_sc_hd__or2_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4766__B1 _4763_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5753_ _4328_/X _5020_/A _4708_/A _4891_/A _4345_/A VGND VGND VPWR VPWR _5753_/X
+ sky130_fd_sc_hd__a41o_2
XANTENNA__3569__B2 _3568_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4704_ _4483_/A _4485_/A _5188_/D VGND VGND VPWR VPWR _4891_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__5963__C1 _4541_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4323__A _4354_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4781__A3 _4928_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5684_ _4556_/X _5680_/X _5682_/X _5683_/Y VGND VGND VPWR VPWR _5684_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_30_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4635_ _4864_/D _5188_/C _4955_/A _4472_/X VGND VGND VPWR VPWR _5721_/A sky130_fd_sc_hd__o211ai_4
XANTENNA__4042__B _4073_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4566_ _4566_/A VGND VGND VPWR VPWR _4580_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3741__A1 _3509_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5730__A2 _4671_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3517_ _3748_/A VGND VGND VPWR VPWR _3517_/X sky130_fd_sc_hd__buf_2
XANTENNA__3881__B _3881_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4497_ _4859_/D _5715_/B _4518_/A _4390_/X VGND VGND VPWR VPWR _5125_/A sky130_fd_sc_hd__a31o_2
X_3448_ _3338_/Y _3571_/C _3447_/X _3571_/A VGND VGND VPWR VPWR _3448_/Y sky130_fd_sc_hd__o31ai_1
X_3379_ _3606_/A _3432_/B VGND VGND VPWR VPWR _3904_/C sky130_fd_sc_hd__and2_2
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _6197_/CLK _6167_/D VGND VGND VPWR VPWR _6167_/Q sky130_fd_sc_hd__dfxtp_1
X_5118_ _5118_/A _5118_/B _5118_/C _5118_/D VGND VGND VPWR VPWR _5118_/Y sky130_fd_sc_hd__nand4_4
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5246__A1 _5687_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4049__A2 _3553_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6098_ _6207_/CLK _6098_/D VGND VGND VPWR VPWR _6098_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3402__A _3876_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5049_ _4552_/X _4783_/X _4890_/A _5048_/X _4935_/X VGND VGND VPWR VPWR _5049_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5797__A2 _5792_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4217__B _4217_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6135__D _6135_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5549__A2 _4218_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4757__B1 _4882_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5329__A _5329_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4233__A _4233_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3980__A1 _3338_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3496__B1 _3495_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5999__A _5999_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5485__B2 _6121_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5485__A1 _4803_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3312__A _3383_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4408__A _4533_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5788__A2 _5787_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output125_A _3025_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4460__A2 _4462_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6045__D _6045_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4748__B1 _5022_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3966__B _3966_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5945__C1 _4964_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4143__A _4143_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5960__A2 _5899_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3971__A1 _3962_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4420_ _4420_/A VGND VGND VPWR VPWR _4420_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5173__B1 _4959_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4797__B _4974_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3723__A1 _3701_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4351_ _4566_/A VGND VGND VPWR VPWR _4832_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3261__B_N _3311_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4920__B1 _4919_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3723__B2 _3524_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4282_ _4282_/A VGND VGND VPWR VPWR _4293_/A sky130_fd_sc_hd__clkbuf_4
X_3302_ _3806_/A VGND VGND VPWR VPWR _3302_/X sky130_fd_sc_hd__buf_2
XFILLER_113_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3233_ _3233_/A VGND VGND VPWR VPWR _3582_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6021_ _6155_/CLK _6021_/D VGND VGND VPWR VPWR _6021_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3164_ _3876_/B VGND VGND VPWR VPWR _4004_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5779__A2 _5745_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3222__A _3648_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3239__B1 _3238_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3095_ _3095_/A VGND VGND VPWR VPWR _3095_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5140__C _5140_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4451__A2 _4346_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3876__B _3876_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3997_ _3781_/B _3781_/C _3781_/D VGND VGND VPWR VPWR _3998_/D sky130_fd_sc_hd__o21a_1
XANTENNA__5936__C1 _4823_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5805_ _5805_/A _5805_/B _5805_/C VGND VGND VPWR VPWR _5805_/X sky130_fd_sc_hd__and3_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5951__A2 _4918_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5736_ _5733_/Y _5734_/X _5735_/X VGND VGND VPWR VPWR _5736_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5667_ _5667_/A _5667_/B _5899_/A VGND VGND VPWR VPWR _5667_/X sky130_fd_sc_hd__and3_1
X_4618_ _4742_/A VGND VGND VPWR VPWR _4618_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5164__B1 _5163_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5583__S _5583_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3714__A1 _3613_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5598_ _5598_/A VGND VGND VPWR VPWR _6158_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5703__A2 _5702_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4549_ _4549_/A VGND VGND VPWR VPWR _4680_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4500__B _6141_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4911__B1 _4984_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5467__A1 _4977_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5467__B2 _6115_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3478__B1 _3477_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4690__A2 _5667_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_85_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5219__A1 _5216_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3132__A input3/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5675__A1_N _6181_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5942__A2 _5880_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3953__A1 _3867_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5155__B1 _4794_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4902__B1 _4901_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3705__A1 _3343_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3307__A _3797_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5458__B2 input13/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5458__A1 input21/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4130__A1 _3583_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4681__A2 _4551_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4418__C1 _4369_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4969__B1 _4968_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3042__A _3042_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3920_ _3477_/X _3831_/X _3359_/B _3919_/X _3917_/X VGND VGND VPWR VPWR _3920_/Y
+ sky130_fd_sc_hd__a41oi_1
XANTENNA__5630__A1 _6041_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5918__C1 _5880_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3851_ _4135_/B _3659_/D _3215_/X _3868_/A VGND VGND VPWR VPWR _3851_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_20_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3782_ _3781_/X _3380_/X _3528_/A VGND VGND VPWR VPWR _3782_/X sky130_fd_sc_hd__a21o_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4736__A3 _5867_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5933__A2 _4740_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3944__B2 _6035_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5521_ _4980_/Y _5433_/X _5504_/A VGND VGND VPWR VPWR _5521_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4601__A _4601_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5146__B1 _4668_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5697__A1 _4870_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5452_ _4977_/X _5412_/X _5701_/C _5451_/X _6111_/Q VGND VGND VPWR VPWR _5453_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4403_ _5240_/C VGND VGND VPWR VPWR _4403_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5697__B2 _4679_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5383_ _5383_/A _5383_/B _5383_/C VGND VGND VPWR VPWR _5383_/X sky130_fd_sc_hd__and3_1
XFILLER_99_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3217__A _3621_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4334_ _4293_/A _4244_/A _4308_/A _4245_/A _6137_/Q VGND VGND VPWR VPWR _4364_/A
+ sky130_fd_sc_hd__o41ai_4
XFILLER_101_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5449__A1 _5444_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4265_ _4265_/A _4283_/A _4265_/C VGND VGND VPWR VPWR _4266_/A sky130_fd_sc_hd__nor3_4
XANTENNA__4974__C _4974_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4121__A1 _3828_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6004_ _6203_/Q _5293_/X _5288_/X VGND VGND VPWR VPWR _6004_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5432__A _5432_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3216_ _3275_/B VGND VGND VPWR VPWR _3621_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_86_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4196_ input7/X VGND VGND VPWR VPWR _4227_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3147_ _3272_/A VGND VGND VPWR VPWR _3446_/B sky130_fd_sc_hd__buf_2
XANTENNA__4409__C1 _4369_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4048__A _4048_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3880__B1 _3624_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5082__C1 _5081_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3078_ _3078_/A VGND VGND VPWR VPWR _3078_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5621__A1 _6037_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5385__B1 _5383_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3935__A1 _3695_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6108__CLK _6145_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5719_ _4666_/A _4582_/X _5717_/Y _5955_/D VGND VGND VPWR VPWR _5719_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5607__A _5618_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5137__B1 _4693_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5688__A1 _5653_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4511__A _5772_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4230__B _4230_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4360__A1 _4243_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4112__B2 _4152_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4112__A1 _3557_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5860__A1 _4890_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4663__A2 _5263_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3797__A _3797_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5612__A1 _6033_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4405__B _4405_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5915__A2 _5911_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4124__C _4124_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4421__A _4421_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5128__B1 _5095_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5679__A1 _5676_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5143__A3 _5743_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4050_ _3626_/X _3832_/A _4089_/A _3520_/X VGND VGND VPWR VPWR _4050_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5300__A0 _6190_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5851__A1 _4360_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5851__B2 _5025_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput6 memory_dmem_request_put[32] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3001_ _3056_/S VGND VGND VPWR VPWR _3010_/S sky130_fd_sc_hd__buf_2
XFILLER_91_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5603__A1 _6029_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3500__A _3500_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4952_ _4952_/A _4952_/B _4952_/C VGND VGND VPWR VPWR _4974_/A sky130_fd_sc_hd__nand3_1
XFILLER_51_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4883_ _4883_/A VGND VGND VPWR VPWR _5878_/C sky130_fd_sc_hd__clkbuf_4
X_3903_ _3830_/C _3834_/X _3902_/X _3488_/X VGND VGND VPWR VPWR _3903_/Y sky130_fd_sc_hd__o31ai_1
XANTENNA__3090__A1 _6079_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3200__A2_N _3197_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3834_ _4135_/B VGND VGND VPWR VPWR _3834_/X sky130_fd_sc_hd__buf_2
XANTENNA__4709__A3 _4891_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3917__A1 _3815_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5906__A2 _5395_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3765_ _3867_/A _3767_/D _3882_/B _3749_/C VGND VGND VPWR VPWR _3765_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3917__B2 _3628_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5119__B1 _4582_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4590__A1 _4673_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4590__B2 _4574_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3873__C _3966_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3393__A2 _3380_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3696_ _3580_/X _3596_/Y _3539_/X _3695_/X VGND VGND VPWR VPWR _3696_/Y sky130_fd_sc_hd__o211ai_1
X_5504_ _5504_/A VGND VGND VPWR VPWR _5504_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5435_ _5435_/A _5528_/B VGND VGND VPWR VPWR _6108_/D sky130_fd_sc_hd__nand2_1
XANTENNA__4342__A1 _4340_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5366_ _5366_/A VGND VGND VPWR VPWR _6096_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4317_ _4317_/A VGND VGND VPWR VPWR _4482_/B sky130_fd_sc_hd__inv_2
XANTENNA__5162__A _5162_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5297_ _5365_/S VGND VGND VPWR VPWR _5306_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_101_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4248_ _4405_/C VGND VGND VPWR VPWR _4859_/B sky130_fd_sc_hd__clkbuf_4
Xclkbuf_4_10_0_CLK clkbuf_3_5_0_CLK/X VGND VGND VPWR VPWR _6123_/CLK sky130_fd_sc_hd__clkbuf_2
XANTENNA__4645__A2 _5721_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5842__A1 _5018_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3448__A3 _3447_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3853__B1 _3852_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4179_ _4218_/C _4218_/D VGND VGND VPWR VPWR _4231_/B sky130_fd_sc_hd__nor2_1
XFILLER_28_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3605__B1 _3308_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4506__A _5643_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5070__A2 _4369_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3410__A _3410_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3081__A1 _6075_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3767__D _3767_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6143__D _6143_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4030__B1 _4029_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3908__A1 _3340_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6080__CLK _6176_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4241__A _4807_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5530__B1 _5491_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input49_A memory_dmem_request_put[75] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3439__A3 _4092_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4097__B1 _3573_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5833__B2 _4328_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5833__A1 _4332_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4100__A4 _4083_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4416__A _4585_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5597__A0 _6158_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3072__A1 _6071_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4135__B _4135_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6053__D _6053_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6010__A1 _3060_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4021__B1 _3161_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3550_ _3397_/A _3592_/A _3657_/C _3582_/B VGND VGND VPWR VPWR _3551_/A sky130_fd_sc_hd__a22o_2
XFILLER_6_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4324__A1 _4527_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3481_ _3876_/A _3588_/C VGND VGND VPWR VPWR _3482_/A sky130_fd_sc_hd__nor2_1
XANTENNA__4301__D _4301_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5220_ _5220_/A _5220_/B _5220_/C VGND VGND VPWR VPWR _5220_/Y sky130_fd_sc_hd__nand3_2
XFILLER_102_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4324__B2 _4527_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5521__B1 _5504_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5151_ _5755_/B _4524_/X _4829_/Y _4574_/X _4316_/X VGND VGND VPWR VPWR _5151_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_96_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5194__B1_N _5193_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3678__A3 _3677_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5082_ _4644_/X _5078_/X _5079_/X _4345_/X _5081_/Y VGND VGND VPWR VPWR _5082_/Y
+ sky130_fd_sc_hd__o311ai_4
XFILLER_96_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4102_ _4102_/A _4102_/B _4102_/C VGND VGND VPWR VPWR _4103_/D sky130_fd_sc_hd__or3_2
XFILLER_110_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5824__A1 _4960_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3214__B _3746_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4627__A2 _4569_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4033_ _4018_/X _4024_/Y _4032_/X VGND VGND VPWR VPWR _6039_/D sky130_fd_sc_hd__a21o_1
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5710__A _5710_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5037__C1 _5036_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4326__A _4354_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3850__A3 _3571_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5588__A0 _6154_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5052__A2 _4748_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3230__A _3882_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5984_ _6197_/Q _5998_/B VGND VGND VPWR VPWR _5984_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4935_ _5118_/C VGND VGND VPWR VPWR _4935_/X sky130_fd_sc_hd__clkbuf_2
X_4866_ _5829_/C _4864_/Y _4865_/Y _5006_/A VGND VGND VPWR VPWR _4866_/X sky130_fd_sc_hd__a31o_1
XFILLER_33_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4797_ _4797_/A _4974_/C _4797_/C VGND VGND VPWR VPWR _4797_/Y sky130_fd_sc_hd__nand3_1
X_3817_ _3668_/X _3910_/A _3536_/A _3464_/X VGND VGND VPWR VPWR _3817_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4061__A _4061_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5760__B1 _5759_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3748_ _3748_/A _3748_/B _3748_/C _3748_/D VGND VGND VPWR VPWR _3748_/X sky130_fd_sc_hd__or4_1
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4996__A _4996_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3679_ _3679_/A VGND VGND VPWR VPWR _3679_/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__4315__A1 _5061_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4315__B2 _4699_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5418_ _5422_/B VGND VGND VPWR VPWR _5528_/B sky130_fd_sc_hd__clkbuf_4
Xoutput140 _2997_/X VGND VGND VPWR VPWR memory_imem_response_get[2] sky130_fd_sc_hd__buf_2
XFILLER_0_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5512__B1 _5447_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3669__A3 _3278_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4866__A2 _4864_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5349_ _5349_/A VGND VGND VPWR VPWR _6088_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3405__A _3781_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4079__B1 _3517_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5815__A1 _5754_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6138__D _6138_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5620__A _5620_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3826__B1 _3816_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4094__A3 _3549_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4236__A _5013_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5579__A0 _6150_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3140__A _3353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5043__A2 _4978_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3054__A1 _6176_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4038__A1_N _3583_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4003__B1 _3512_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4554__A1 _4680_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5067__A _5067_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4554__B2 _4552_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4306__A1 _4890_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4857__A2 _4852_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5514__B _5531_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3315__A _3315_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4609__A2 _4362_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5806__A1 _6115_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6048__D _6048_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3817__B1 _3536_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5282__A2 _3822_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5019__C1 _5018_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4146__A _4146_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2981_ _6099_/Q _6098_/Q _6097_/Q VGND VGND VPWR VPWR _4186_/A sky130_fd_sc_hd__nand3b_1
XANTENNA__4242__B1 _4239_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3596__A2 _3595_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5990__B1 _5288_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4720_ _4716_/X _4513_/X input37/X _5805_/B _4719_/X VGND VGND VPWR VPWR _4720_/X
+ sky130_fd_sc_hd__o311a_4
X_4651_ _4780_/A VGND VGND VPWR VPWR _4652_/A sky130_fd_sc_hd__clkbuf_4
X_3602_ _3366_/A _3432_/B _3330_/A VGND VGND VPWR VPWR _3603_/B sky130_fd_sc_hd__o21bai_4
Xinput31 memory_dmem_request_put[57] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_1
Xinput20 memory_dmem_request_put[46] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5742__B1 _4353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4582_ _4875_/A VGND VGND VPWR VPWR _4582_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3899__A3 _3894_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput53 memory_dmem_request_put[79] VGND VGND VPWR VPWR _4218_/C sky130_fd_sc_hd__clkbuf_2
Xinput42 memory_dmem_request_put[68] VGND VGND VPWR VPWR _5392_/C sky130_fd_sc_hd__clkbuf_1
Xinput64 memory_dmem_request_put[90] VGND VGND VPWR VPWR _4170_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_0_CLK_A CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3533_ _3911_/C VGND VGND VPWR VPWR _3533_/X sky130_fd_sc_hd__clkbuf_4
Xinput75 memory_imem_request_put[11] VGND VGND VPWR VPWR _3918_/A sky130_fd_sc_hd__clkbuf_2
X_3464_ _3574_/A VGND VGND VPWR VPWR _3464_/X sky130_fd_sc_hd__buf_4
XANTENNA__4848__A2 _4847_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5203_ _5203_/A VGND VGND VPWR VPWR _5260_/A sky130_fd_sc_hd__buf_2
XANTENNA__3505__C1 _3504_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6183_ _6204_/CLK _6183_/D VGND VGND VPWR VPWR _6183_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3225__A _3440_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5134_ _5235_/A VGND VGND VPWR VPWR _5743_/B sky130_fd_sc_hd__clkbuf_4
X_3395_ _3377_/Y _3393_/X _3580_/A VGND VGND VPWR VPWR _3396_/B sky130_fd_sc_hd__a21oi_1
XFILLER_69_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5065_ _5061_/X _5062_/X _5063_/X _5064_/X VGND VGND VPWR VPWR _5065_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3808__B1 _3724_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_4_9_0_CLK_A clkbuf_4_9_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5812__A4 _5944_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4016_ _3343_/X _3829_/X _3194_/X _3533_/X _4124_/A VGND VGND VPWR VPWR _4016_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4076__A3 _3479_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3284__A1 _3359_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5273__A2 input3/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3284__B2 _3359_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3823__A3 _3821_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5025__A2 _4619_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3895__A _3895_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5967_ _6195_/Q _4799_/X _5958_/Y _5966_/Y VGND VGND VPWR VPWR _6195_/D sky130_fd_sc_hd__o22a_1
XANTENNA__5586__S _5594_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3587__A2 _3983_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4918_ _4918_/A VGND VGND VPWR VPWR _5148_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__4784__A1 _4243_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5981__B1 _5237_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5898_ _4353_/X _5021_/X _5192_/X _5878_/Y _4403_/X VGND VGND VPWR VPWR _5898_/X
+ sky130_fd_sc_hd__o311a_1
X_4849_ _4685_/X _4818_/X _4837_/X _4848_/Y VGND VGND VPWR VPWR _4850_/A sky130_fd_sc_hd__o22ai_4
XFILLER_32_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5615__A _5615_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4839__A2 _4437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5497__C1 _5496_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3135__A _3754_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5500__A3 _5498_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5567__A3 _4803_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4775__A1 _4692_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5972__B1 _5720_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3578__A2 _3569_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5509__B _5531_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5724__B1 _5716_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5525__A _5525_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3750__A2 _3716_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3045__A _5985_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3180_ _3226_/A VGND VGND VPWR VPWR _3442_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3502__A2 _3457_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4160__C1 _3717_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5260__A _5260_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4463__B1 _4815_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5660__C1 _4675_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3266__B2 _3882_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3266__A1 _3254_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3805__A3 _3800_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5007__A2 _5118_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5821_ _6101_/Q _4807_/A _5905_/A _5820_/X VGND VGND VPWR VPWR _5822_/B sky130_fd_sc_hd__o211a_1
XANTENNA__4604__A _4604_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4766__A1 _4749_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4766__B2 _4765_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5963__B1 _4870_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5752_ _5743_/A _5743_/B _5706_/Y _5145_/A VGND VGND VPWR VPWR _5752_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_34_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4703_ _5003_/B VGND VGND VPWR VPWR _5152_/A sky130_fd_sc_hd__buf_4
XANTENNA__4781__A4 _4779_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5683_ _4422_/A _4699_/X _5060_/X _5033_/Y VGND VGND VPWR VPWR _5683_/Y sky130_fd_sc_hd__o22ai_4
XANTENNA__4042__C _4042_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6141__CLK _6145_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5750__A2_N _5646_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4634_ _4239_/X _4630_/A _4224_/X _4633_/X VGND VGND VPWR VPWR _4634_/X sky130_fd_sc_hd__a2bb2o_1
X_4565_ _4565_/A VGND VGND VPWR VPWR _5755_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3726__C1 _3302_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4034__C_N _3397_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3741__A2 _3740_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3516_ _3512_/X _3410_/B _3320_/Y _3748_/B VGND VGND VPWR VPWR _3516_/Y sky130_fd_sc_hd__a31oi_1
XANTENNA__5730__A3 _5944_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5435__A _5435_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4496_ _4520_/A VGND VGND VPWR VPWR _4859_/D sky130_fd_sc_hd__buf_2
XFILLER_103_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3447_ _3621_/C _3527_/C _3447_/C VGND VGND VPWR VPWR _3447_/X sky130_fd_sc_hd__and3_2
XFILLER_97_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3378_ _3436_/B VGND VGND VPWR VPWR _4034_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__4151__C1 _3862_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6203_/CLK _6166_/D VGND VGND VPWR VPWR _6166_/Q sky130_fd_sc_hd__dfxtp_1
X_5117_ _4551_/Y _4996_/A _4887_/X _5721_/C VGND VGND VPWR VPWR _5117_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ _6207_/CLK _6097_/D VGND VGND VPWR VPWR _6097_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5246__A2 _4604_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5170__A _5170_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5048_ _5048_/A VGND VGND VPWR VPWR _5048_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4217__C _4217_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4757__A1 _4369_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5549__A3 _5529_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4514__A _4976_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5954__B1 _4657_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6151__D _6151_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3980__A2 _3978_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5890__A1_N _4824_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5345__A _5345_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3496__A1 _3968_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4142__C1 _4149_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5999__B _5999_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5485__A2 _5161_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input31_A memory_dmem_request_put[57] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output118_A _3078_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4460__A3 _4769_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4424__A _4860_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4748__A1 _5899_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3966__C _3966_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5945__B1 _5944_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6164__CLK _6203_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4143__B _4143_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5960__A3 _4965_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6061__D _6061_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3971__A2 _3963_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5173__A1 _4673_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4350_ _4350_/A VGND VGND VPWR VPWR _5018_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__4797__C _4797_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4920__A1 _5148_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3723__A2 _3512_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3301_ _3301_/A VGND VGND VPWR VPWR _3806_/A sky130_fd_sc_hd__clkbuf_2
X_4281_ _4738_/B VGND VGND VPWR VPWR _4815_/C sky130_fd_sc_hd__buf_2
XFILLER_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3232_ _3667_/B VGND VGND VPWR VPWR _3557_/A sky130_fd_sc_hd__clkbuf_2
X_6020_ _6155_/CLK _6020_/D VGND VGND VPWR VPWR _6020_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ _3513_/A VGND VGND VPWR VPWR _3876_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__5881__C1 _5004_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3503__A _3537_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3239__A1 _3218_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3094_ _6053_/Q _6081_/Q _3094_/S VGND VGND VPWR VPWR _3095_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5140__D _5140_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4451__A3 _4389_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2998__A0 _6019_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5804_ _5175_/X _5797_/Y _5803_/Y _5673_/A VGND VGND VPWR VPWR _5804_/Y sky130_fd_sc_hd__o211ai_4
X_3996_ _3645_/A _3994_/X _4044_/C _3849_/X VGND VGND VPWR VPWR _3996_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__5936__B1 _4708_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5735_ _5712_/A _4556_/X _5050_/Y _4950_/A VGND VGND VPWR VPWR _5735_/X sky130_fd_sc_hd__o31a_2
XANTENNA__3947__C1 _3799_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5666_ _5782_/A _4773_/Y _4965_/Y _4730_/Y _5731_/A VGND VGND VPWR VPWR _5666_/Y
+ sky130_fd_sc_hd__a32oi_1
XANTENNA__5951__A3 _5098_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4617_ _4707_/D _4619_/B _5034_/C _4946_/A VGND VGND VPWR VPWR _4617_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__5164__A1 _5161_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5597_ _6158_/Q _6026_/Q _5605_/S VGND VGND VPWR VPWR _5598_/A sky130_fd_sc_hd__mux2_1
X_4548_ _5976_/B _5971_/B _4547_/Y VGND VGND VPWR VPWR _4548_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3714__A2 _3707_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4911__B2 _5162_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4479_ _4543_/A VGND VGND VPWR VPWR _4960_/A sky130_fd_sc_hd__buf_2
XFILLER_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3478__A1 _3466_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5467__A2 _5433_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6037__CLK _6045_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5872__C1 _4984_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3413__A _3642_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5219__A2 _5218_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3830__A_N _3829_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4509__A _4975_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6149_ _6197_/CLK _6149_/D VGND VGND VPWR VPWR _6149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4427__B1 _4261_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_3_6_0_CLK_A clkbuf_3_7_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6146__D _6146_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6187__CLK _6204_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5927__B1 _4563_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4244__A _4244_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3953__A2 _3975_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5155__A1 _5140_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input79_A memory_imem_request_put[5] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4902__A1 _4403_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3705__A2 _3893_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5458__A2 _5437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4419__A _4584_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3323__A _3992_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4130__A2 _3515_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4681__A3 _5079_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4418__B1 _4957_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4851__A2_N _6050_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4969__A1 _4957_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6056__D _6056_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5918__B1 _5068_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3850_ _3525_/X _3631_/X _3571_/B _3849_/X VGND VGND VPWR VPWR _3850_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3929__C1 _3376_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3781_ _3781_/A _3781_/B _3781_/C _3781_/D VGND VGND VPWR VPWR _3781_/X sky130_fd_sc_hd__or4_4
XFILLER_20_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5520_ _5520_/A VGND VGND VPWR VPWR _6131_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5146__A1 _5680_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5146__B2 _4726_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5451_ _5499_/A VGND VGND VPWR VPWR _5451_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4402_ _5003_/B VGND VGND VPWR VPWR _5944_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5697__A2 _4440_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5382_ _6099_/Q _5382_/B VGND VGND VPWR VPWR _5383_/C sky130_fd_sc_hd__nand2_1
XFILLER_99_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4333_ _4333_/A VGND VGND VPWR VPWR _4362_/A sky130_fd_sc_hd__clkinv_2
X_4264_ _4268_/A _4293_/B _4264_/C _4309_/A VGND VGND VPWR VPWR _4602_/A sky130_fd_sc_hd__nor4_4
XFILLER_5_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5449__A2 _5445_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5854__C1 _4928_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_86_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3215_ _3710_/C VGND VGND VPWR VPWR _3215_/X sky130_fd_sc_hd__buf_4
X_6003_ _3060_/S _5291_/X _6009_/A _5540_/A _6002_/X VGND VGND VPWR VPWR _6202_/D
+ sky130_fd_sc_hd__a311o_1
XANTENNA__4329__A _4601_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3233__A _3233_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4121__A2 _4109_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4195_ _4195_/A VGND VGND VPWR VPWR _4718_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3146_ _3387_/B VGND VGND VPWR VPWR _3272_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4409__B1 _4864_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4048__B _4048_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3880__A1 _3863_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3077_ _6181_/Q _6073_/Q _3083_/S VGND VGND VPWR VPWR _3078_/A sky130_fd_sc_hd__mux2_2
XFILLER_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5082__B1 _4345_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5909__B1 _5894_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4999__A _4999_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5385__B2 _5383_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5385__A1 _6098_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5718_ _5761_/D _4996_/A _4887_/X _4924_/A VGND VGND VPWR VPWR _5955_/D sky130_fd_sc_hd__a31o_2
X_3979_ _3660_/B _4004_/A _3495_/X _4116_/A VGND VGND VPWR VPWR _3979_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3935__A2 _3931_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5594__S _5594_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5137__A1 _4702_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5649_ _5045_/A _5440_/X _5403_/X _5163_/X VGND VGND VPWR VPWR _5649_/X sky130_fd_sc_hd__a211o_1
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5688__A2 _5687_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4230__C _4230_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4360__A2 _4293_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4648__B1 _5148_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3143__A _3226_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4112__A2 _4042_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4239__A _5643_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5860__A2 _5018_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3320__B1 _3319_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2982__A _4186_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4820__B1 _4942_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4405__C _4405_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4124__D _4124_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4702__A _4702_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6202__CLK _6202_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5128__B2 _5127_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3318__A _3586_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5679__A2 _5678_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5143__A4 _4945_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4149__A _4149_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3053__A _3053_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5300__A1 _6066_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_83_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5851__A2 _4960_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput7 memory_dmem_request_put[33] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_2
X_3000_ _5985_/B VGND VGND VPWR VPWR _3056_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_37_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5064__B1 _4621_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4951_ _4938_/X _4941_/Y _4949_/Y _4950_/X VGND VGND VPWR VPWR _4952_/C sky130_fd_sc_hd__o211ai_4
XFILLER_45_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4882_ _4882_/A VGND VGND VPWR VPWR _4882_/X sky130_fd_sc_hd__buf_4
X_3902_ _3902_/A _4074_/A VGND VGND VPWR VPWR _3902_/X sky130_fd_sc_hd__and2_1
XFILLER_51_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3833_ _3831_/X _3975_/A _3488_/X _3439_/X VGND VGND VPWR VPWR _3833_/X sky130_fd_sc_hd__o22a_1
XFILLER_32_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3764_ _3938_/B VGND VGND VPWR VPWR _3764_/X sky130_fd_sc_hd__buf_4
XANTENNA__3917__A2 _3910_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5119__A1 _5117_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4590__A2 _4996_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3393__A3 _3382_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3695_ _3695_/A _3695_/B _3695_/C _3694_/X VGND VGND VPWR VPWR _3695_/X sky130_fd_sc_hd__or4b_1
X_5503_ _5503_/A VGND VGND VPWR VPWR _5504_/A sky130_fd_sc_hd__buf_2
XANTENNA__3228__A _3621_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5434_ _6108_/Q _5425_/B _5968_/A _5433_/X VGND VGND VPWR VPWR _5435_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__4342__A2 _5818_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3550__B1 _3657_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5365_ _6052_/Q _6096_/Q _5365_/S VGND VGND VPWR VPWR _5366_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5443__A _5443_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5827__C1 _5721_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4316_ _5235_/A VGND VGND VPWR VPWR _4316_/X sky130_fd_sc_hd__buf_4
X_5296_ _5352_/A VGND VGND VPWR VPWR _5365_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4247_ _4247_/A VGND VGND VPWR VPWR _4910_/A sky130_fd_sc_hd__buf_2
XANTENNA__5992__B1_N _5985_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5842__A2 _5098_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4178_ _4218_/A _4218_/B VGND VGND VPWR VPWR _4231_/A sky130_fd_sc_hd__nor2_1
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3853__A1 _3850_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5055__B1 _4793_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3129_ _6064_/Q _6063_/Q _6062_/Q VGND VGND VPWR VPWR _3129_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_28_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3605__A1 _3496_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3605__B2 _3604_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3410__B _3410_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5618__A _5618_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4030__A1 _3376_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3908__A2 _3901_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4522__A _4522_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3138__A _4044_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3129__A_N _6064_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5530__B2 _6135_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5530__A1 _5523_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2977__A _6199_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4097__A1 _3512_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3439__A4 _3732_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4097__B2 _3873_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5833__A2 _5018_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_3_0_CLK_A clkbuf_2_3_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5597__A1 _6026_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output100_A _3104_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3780__D_N _3611_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4135__C _4135_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5528__A _5528_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6010__A2 _5291_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4432__A _4432_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4021__A1 _4019_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3480_ _3480_/A VGND VGND VPWR VPWR _3588_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5473__A2_N _5405_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4324__A2 _4536_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5263__A _5263_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5521__A1 _4980_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5150_ _5150_/A _5150_/B _5150_/C VGND VGND VPWR VPWR _5150_/Y sky130_fd_sc_hd__nor3_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5081_ _4661_/X _4464_/X _5080_/X _5021_/X _4957_/A VGND VGND VPWR VPWR _5081_/Y
+ sky130_fd_sc_hd__o221ai_4
X_4101_ _4099_/X _4100_/X _3862_/A VGND VGND VPWR VPWR _4102_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__5809__C1 _5163_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5824__A2 _4840_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4032_ _4031_/X _3787_/X _3763_/X _6039_/Q _3891_/A VGND VGND VPWR VPWR _4032_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5488__A2_N _4239_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3511__A _3841_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5037__B1 _4685_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5983_ _5970_/X _5982_/Y _4190_/X _6196_/Q VGND VGND VPWR VPWR _6196_/D sky130_fd_sc_hd__o2bb2a_1
XANTENNA__5588__A1 _6022_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3733__B1_N _3528_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4934_ _4934_/A _4934_/B VGND VGND VPWR VPWR _4952_/A sky130_fd_sc_hd__nand2_1
XFILLER_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3599__B1 _6020_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4865_ _4865_/A _5048_/A _4865_/C _4865_/D VGND VGND VPWR VPWR _4865_/Y sky130_fd_sc_hd__nand4_2
XFILLER_32_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4796_ _4782_/X _4790_/X _4795_/X _4568_/X VGND VGND VPWR VPWR _4797_/C sky130_fd_sc_hd__a31o_1
XANTENNA__4012__A1 _3525_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3816_ _3816_/A _3816_/B _3816_/C _3816_/D VGND VGND VPWR VPWR _3816_/X sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_4_5_0_CLK_A clkbuf_4_5_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3747_ _3299_/A _3319_/X _3968_/C _3593_/X VGND VGND VPWR VPWR _3748_/D sky130_fd_sc_hd__a31o_1
XANTENNA__5760__A1 _5754_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3771__B1 _6026_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3678_ _3665_/X _3290_/X _3677_/Y _6022_/Q _3541_/X VGND VGND VPWR VPWR _6022_/D
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4315__A2 _4787_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5417_ _6104_/Q _5425_/B VGND VGND VPWR VPWR _5417_/Y sky130_fd_sc_hd__nor2_1
Xoutput130 _3036_/X VGND VGND VPWR VPWR memory_imem_response_get[19] sky130_fd_sc_hd__buf_2
Xoutput141 _3055_/X VGND VGND VPWR VPWR memory_imem_response_get[30] sky130_fd_sc_hd__buf_2
XANTENNA__5512__A1 _6128_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4866__A3 _4865_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5348_ _6059_/Q _6088_/Q _5350_/S VGND VGND VPWR VPWR _5349_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4720__C1 _4719_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4079__A1 _4124_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5815__A2 _5796_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5279_ _5285_/A _5279_/B VGND VGND VPWR VPWR _5279_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3826__A1 _3825_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3826__B2 _3778_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5579__A1 _6018_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6154__D _6154_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4252__A _4950_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4003__A1 _3867_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4554__A2 _5079_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3211__C1 _3692_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4003__B2 _4152_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5200__B1 _5166_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input61_A memory_dmem_request_put[87] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4306__A2 _5971_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3514__B1 _3600_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4857__A3 _4855_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4711__C1 _4710_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3315__B _3606_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4609__A3 _4910_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output148_A _3011_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5806__A2 _5643_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5811__A _5811_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3817__A1 _3668_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5019__B1 _4652_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3331__A _3802_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4146__B _4146_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6064__D _6064_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2980_ _6178_/Q VGND VGND VPWR VPWR _5640_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__4242__B2 _4241_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3450__C1 _3449_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5990__A1 _6198_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4650_ _4855_/D _5899_/B _5710_/A _4879_/A VGND VGND VPWR VPWR _4650_/X sky130_fd_sc_hd__or4_1
XANTENNA__5258__A _5545_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3601_ _3406_/A _3779_/C _3746_/B _4073_/D VGND VGND VPWR VPWR _3601_/X sky130_fd_sc_hd__o211a_1
Xinput10 memory_dmem_request_put[36] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_4
Xinput21 memory_dmem_request_put[47] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4581_ _5034_/B _5711_/B _4581_/C _5078_/A VGND VGND VPWR VPWR _4581_/Y sky130_fd_sc_hd__nand4_4
XANTENNA__5742__B2 _5741_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3753__B1 _3577_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput54 memory_dmem_request_put[80] VGND VGND VPWR VPWR _4218_/B sky130_fd_sc_hd__clkbuf_1
Xinput43 memory_dmem_request_put[69] VGND VGND VPWR VPWR _5438_/D sky130_fd_sc_hd__clkbuf_1
Xinput32 memory_dmem_request_put[58] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3532_ _4065_/A VGND VGND VPWR VPWR _3830_/C sky130_fd_sc_hd__buf_2
Xinput76 memory_imem_request_put[2] VGND VGND VPWR VPWR _3226_/A sky130_fd_sc_hd__buf_4
Xinput65 memory_dmem_request_put[91] VGND VGND VPWR VPWR _4170_/A sky130_fd_sc_hd__clkbuf_1
X_3463_ _3543_/B _4042_/D _3460_/X _3761_/A VGND VGND VPWR VPWR _3463_/X sky130_fd_sc_hd__o22a_1
XFILLER_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6182_ _6196_/CLK _6182_/D VGND VGND VPWR VPWR _6182_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3505__B1 _3492_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5202_ input30/X _4804_/X _5042_/X input14/X VGND VGND VPWR VPWR _5202_/Y sky130_fd_sc_hd__a22oi_4
XANTENNA__3506__A _3828_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3225__B _3366_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5133_ _5133_/A VGND VGND VPWR VPWR _5148_/A sky130_fd_sc_hd__buf_4
X_3394_ _3815_/A VGND VGND VPWR VPWR _3580_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5721__A _5721_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5064_ _4707_/C _4350_/A _4852_/A _4621_/A VGND VGND VPWR VPWR _5064_/X sky130_fd_sc_hd__o31a_1
XANTENNA__3808__A1 _3807_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4337__A _5067_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4015_ _3968_/X _4014_/X _3699_/X VGND VGND VPWR VPWR _4015_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__6070__CLK _6074_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3241__A _3476_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3284__A2 _3815_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5966_ _5734_/X _5962_/Y _5940_/X _5965_/Y VGND VGND VPWR VPWR _5966_/Y sky130_fd_sc_hd__a211oi_1
X_4917_ _4917_/A _5761_/B _5878_/C _5079_/C VGND VGND VPWR VPWR _4917_/X sky130_fd_sc_hd__and4_1
X_5897_ _5896_/Y _5068_/X _4773_/Y _4387_/X VGND VGND VPWR VPWR _5897_/X sky130_fd_sc_hd__a31o_1
XFILLER_80_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4784__A2 _4362_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5981__A1 _5708_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5981__B2 _5980_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4848_ _4842_/Y _4847_/X _4568_/X VGND VGND VPWR VPWR _4848_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4779_ _4777_/X _4778_/X _4369_/C _4369_/A VGND VGND VPWR VPWR _4779_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4800__A _4800_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3416__A _3680_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5497__B1 _5288_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6149__D _6149_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5249__B1 _5247_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5631__A _5631_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4247__A _4247_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3151__A _3315_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2990__A _6202_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5421__B1 _5398_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4775__A2 _4864_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5972__A1 _5061_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5078__A _5078_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5185__C1 _4652_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5724__B2 _5723_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5724__A1 _5715_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5525__B _5531_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3326__A _3528_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5488__B1 _4801_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4160__B1 _3482_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6093__CLK _6204_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6059__D _6059_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3502__A3 _3501_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5541__A _5541_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4463__A1 _4649_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5660__B1 _4440_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3266__A2 _3831_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3061__A _3061_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5820_ input9/X _5395_/A _5163_/A _4984_/A VGND VGND VPWR VPWR _5820_/X sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_1_0_0_CLK_A clkbuf_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4766__A2 _4752_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5963__A1 _4431_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5751_ _6185_/Q VGND VGND VPWR VPWR _5751_/Y sky130_fd_sc_hd__inv_2
X_4702_ _4702_/A VGND VGND VPWR VPWR _4708_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3974__B1 _3631_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5682_ _4345_/A _5213_/X _5681_/Y _5140_/C VGND VGND VPWR VPWR _5682_/X sky130_fd_sc_hd__o31a_1
XFILLER_8_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4042__D _4042_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4633_ _4632_/X _6127_/Q _4633_/S VGND VGND VPWR VPWR _4633_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4564_ _4788_/B VGND VGND VPWR VPWR _4565_/A sky130_fd_sc_hd__buf_4
XANTENNA__4620__A _4640_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3726__B1 _3142_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3515_ _4004_/C _3515_/B _3653_/C _3797_/A VGND VGND VPWR VPWR _3748_/B sky130_fd_sc_hd__and4_2
XFILLER_7_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5435__B _5528_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3236__A _3446_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4495_ _4469_/Y _4492_/X _4494_/X VGND VGND VPWR VPWR _4495_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5479__B1 _5451_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3446_ _3603_/D _3446_/B VGND VGND VPWR VPWR _3621_/C sky130_fd_sc_hd__and2_4
XFILLER_69_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3377_ _3361_/Y _3363_/X _3369_/X _3374_/X _3376_/X VGND VGND VPWR VPWR _3377_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__4151__B1 _4150_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6176_/CLK _6165_/D VGND VGND VPWR VPWR _6165_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5451__A _5499_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5116_ _4661_/X _4464_/X _4742_/X _5115_/Y VGND VGND VPWR VPWR _5116_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_85_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ _6204_/CLK _6096_/D VGND VGND VPWR VPWR _6096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5246__A3 _5079_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4067__A _4067_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5047_ _5041_/X _4991_/X _4241_/X _5046_/Y VGND VGND VPWR VPWR _5047_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_65_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5597__S _5605_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4217__D _4217_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4757__A2 _4619_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5954__A1 _4671_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5949_ _5946_/Y _5955_/A _5822_/A _5948_/X VGND VGND VPWR VPWR _5949_/X sky130_fd_sc_hd__a211o_1
XFILLER_41_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3965__B1 _4073_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4530__A _4661_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5626__A _5626_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_3_2_0_CLK_A clkbuf_3_3_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4390__B1 _6140_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3146__A _3387_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3496__A2 _3494_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4142__B1 _3631_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5999__C _6014_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2985__A _5382_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5485__A3 _5445_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5890__B1 _5107_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input24_A memory_dmem_request_put[50] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5642__B1 _5410_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4705__A _4705_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5300__S _5306_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4748__A2 _4621_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5945__A1 _4679_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_4_13_0_CLK_A clkbuf_3_6_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5945__B2 _4657_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5158__C1 _5157_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4440__A _4754_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5173__A2 _4398_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4905__C1 _4904_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5536__A input5/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3982__C _3982_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output92_A _3089_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4920__A2 _5148_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3723__A3 _3722_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3300_ _3881_/A VGND VGND VPWR VPWR _3300_/X sky130_fd_sc_hd__buf_2
X_4280_ _4860_/B VGND VGND VPWR VPWR _4738_/B sky130_fd_sc_hd__clkbuf_2
X_3231_ _3226_/A _3443_/B VGND VGND VPWR VPWR _3667_/B sky130_fd_sc_hd__and2b_1
XANTENNA__4133__B1 _4132_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ _3162_/A VGND VGND VPWR VPWR _3513_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5881__B1 _4930_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3892__C1 _3882_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3239__A2 _3223_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3093_ _3093_/A VGND VGND VPWR VPWR _3093_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2998__A1 _6151_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5803_ _5715_/X _4390_/X _5716_/X _5802_/Y VGND VGND VPWR VPWR _5803_/Y sky130_fd_sc_hd__o22ai_2
X_3995_ _3406_/A _3382_/D _3362_/Y _4073_/D VGND VGND VPWR VPWR _4044_/C sky130_fd_sc_hd__o211a_1
XANTENNA__5936__B2 _4610_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5936__A1 _5097_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3947__B1 _3548_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5734_ _5734_/A VGND VGND VPWR VPWR _5734_/X sky130_fd_sc_hd__clkbuf_2
X_5665_ _4873_/A _4864_/B _4864_/D _4869_/A _4589_/A VGND VGND VPWR VPWR _5731_/A
+ sky130_fd_sc_hd__o311a_1
X_4616_ _4937_/B VGND VGND VPWR VPWR _5034_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__4350__A _4350_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5164__A2 _5772_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5596_ _5618_/A VGND VGND VPWR VPWR _5605_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4547_ _4878_/A _4754_/A _4259_/A _5118_/B _4673_/B VGND VGND VPWR VPWR _4547_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_89_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4478_ _4788_/B VGND VGND VPWR VPWR _4480_/C sky130_fd_sc_hd__buf_2
XFILLER_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3429_ _3574_/A VGND VGND VPWR VPWR _3429_/X sky130_fd_sc_hd__buf_4
XANTENNA__5467__A3 _5805_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3478__A2 _3476_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6148_ _6197_/CLK _6148_/D VGND VGND VPWR VPWR _6148_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5872__B1 _5162_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4427__B2 _4209_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6079_ _6203_/CLK _6079_/D VGND VGND VPWR VPWR _6079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4525__A _4729_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5927__A1 _5118_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6162__D _6162_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3953__A3 _3567_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5155__A2 _5153_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4260__A _4268_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5356__A _5356_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4902__A2 _4894_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3705__A3 _3534_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4115__B1 _4114_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5863__B1 _4387_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5091__A _5162_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3874__C1 _3873_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4130__A3 _3551_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4418__A1 _5148_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output130_A _3036_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4969__A2 _4966_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6131__CLK _6145_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4435__A _4926_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5918__A1 _5021_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6072__D _6072_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3929__B1 _3928_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3780_ _3780_/A _4073_/C _3780_/C _3611_/A VGND VGND VPWR VPWR _3780_/X sky130_fd_sc_hd__or4b_1
XANTENNA__4051__C1 _4050_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5450_ input19/X _5437_/X _5439_/X input11/X VGND VGND VPWR VPWR _5701_/C sky130_fd_sc_hd__a22o_1
XANTENNA__4170__A _4170_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4401_ _4329_/X _4330_/X _4533_/A _4769_/A VGND VGND VPWR VPWR _5003_/B sky130_fd_sc_hd__o211ai_4
XANTENNA__5146__A2 _4739_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5697__A3 _4967_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5381_ _6099_/Q _5381_/B VGND VGND VPWR VPWR _5383_/B sky130_fd_sc_hd__or2_1
X_4332_ _4414_/A VGND VGND VPWR VPWR _4332_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_99_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4106__B1 _3157_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4263_ _4287_/B VGND VGND VPWR VPWR _4293_/B sky130_fd_sc_hd__clkinv_2
XFILLER_5_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5449__A3 _5677_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5854__B1 _4879_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3214_ _4034_/A _3746_/B VGND VGND VPWR VPWR _3710_/C sky130_fd_sc_hd__nand2_4
X_6002_ _3096_/A _5291_/X _5293_/X _6202_/Q VGND VGND VPWR VPWR _6002_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__3865__C1 _3508_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4194_ _4225_/A input7/X _5438_/D VGND VGND VPWR VPWR _4195_/A sky130_fd_sc_hd__and3b_1
X_3145_ _3437_/B VGND VGND VPWR VPWR _3858_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4409__B2 _4864_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4409__A1 _4404_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4048__C _4065_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_67_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3880__A2 _3865_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3076_ _3076_/A VGND VGND VPWR VPWR _3076_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5082__A1 _4644_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4345__A _4345_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4290__C1 _4725_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5909__B2 _5908_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3978_ _4089_/A _3512_/A _3470_/X VGND VGND VPWR VPWR _3978_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5385__A2 _5382_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4593__B1 _4929_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5717_ _4686_/X _5152_/B _5106_/X _4820_/Y VGND VGND VPWR VPWR _5717_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_50_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5176__A _5944_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3935__A3 _3933_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5137__A2 _4891_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5648_ _6145_/Q _5560_/X _5648_/S VGND VGND VPWR VPWR _5676_/A sky130_fd_sc_hd__mux2_4
XANTENNA__4911__A2_N _5640_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5579_ _6150_/Q _6018_/Q _5583_/S VGND VGND VPWR VPWR _5580_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4360__A3 _4910_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4648__A1 _4378_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3424__A _3802_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5845__B1 _5982_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6154__CLK _6155_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_85_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3320__A1 _4089_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6157__D _6157_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4820__A1 _4929_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4405__D _4405_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5781__C1 _4794_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3334__A _3876_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4149__B _4149_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 memory_dmem_request_put[34] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6067__D _6067_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4065__D_N _3495_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5064__A1 _4707_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3075__A0 _6196_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4950_ _4950_/A VGND VGND VPWR VPWR _4950_/X sky130_fd_sc_hd__buf_4
XANTENNA__4165__A input1/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4881_ _4870_/X _4871_/Y _4874_/X _4875_/X _4880_/Y VGND VGND VPWR VPWR _4881_/Y
+ sky130_fd_sc_hd__a311oi_4
X_3901_ _3834_/X _3895_/X _3215_/X _3900_/Y VGND VGND VPWR VPWR _3901_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_51_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3832_ _3832_/A VGND VGND VPWR VPWR _3975_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4024__C1 _3866_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3509__A _3509_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6027__CLK _6197_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5502_ _5502_/A VGND VGND VPWR VPWR _6125_/D sky130_fd_sc_hd__clkbuf_1
X_3763_ _3828_/A VGND VGND VPWR VPWR _3763_/X sky130_fd_sc_hd__buf_2
XANTENNA__5119__A2 _5118_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3694_ _3195_/A _3223_/X _3183_/X _3208_/X _3522_/X VGND VGND VPWR VPWR _3694_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_118_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3228__B _3500_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5433_ _5433_/A VGND VGND VPWR VPWR _5433_/X sky130_fd_sc_hd__buf_2
XANTENNA__6177__CLK _6201_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5364_ _5364_/A VGND VGND VPWR VPWR _6095_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3550__A1 _3397_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4315_ _5061_/A _4787_/A _4421_/A _4699_/A VGND VGND VPWR VPWR _5235_/A sky130_fd_sc_hd__o22a_1
XANTENNA__5827__B1 _4953_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3550__B2 _3582_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3244__A _3315_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5295_ _5291_/X _5292_/Y _5293_/X _5294_/X VGND VGND VPWR VPWR _5352_/A sky130_fd_sc_hd__a211oi_2
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4246_ _4246_/A _4246_/B _4246_/C VGND VGND VPWR VPWR _4247_/A sky130_fd_sc_hd__or3_1
XFILLER_19_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4177_ _4230_/A _4230_/B _4230_/C VGND VGND VPWR VPWR _4265_/A sky130_fd_sc_hd__nand3_4
XANTENNA_clkbuf_4_1_0_CLK_A clkbuf_4_1_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3853__A2 _3851_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3128_ _3128_/A VGND VGND VPWR VPWR _3128_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5055__A1 _5720_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3605__A2 _3601_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3059_ _3059_/A VGND VGND VPWR VPWR _3059_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3066__A0 _6192_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6004__B1 _5288_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4803__A _5044_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4030__A2 _4026_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3908__A3 _3903_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4522__B _5968_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4318__B1 _6136_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5530__A2 _4285_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3154__A _3233_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5818__A0 _6144_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4097__A2 _4152_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5833__A3 _5148_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2993__A _2993_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5796__A1_N _4858_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5528__B _5528_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4557__B1 _4554_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3329__A _4092_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4021__A2 _3139_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3444__A2_N _3437_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5506__C1 _5505_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5544__A _5544_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5521__A2 _5433_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4063__B1_N _4036_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5809__B1 _5403_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5080_ _4864_/D _5008_/A _5009_/X _4259_/A VGND VGND VPWR VPWR _5080_/X sky130_fd_sc_hd__a31o_4
X_4100_ _3653_/A _3293_/X _3965_/Y _4083_/B _3900_/Y VGND VGND VPWR VPWR _4100_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_111_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5824__A3 _5971_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4031_ _3685_/X _3962_/X _3414_/X _4030_/Y VGND VGND VPWR VPWR _4031_/X sky130_fd_sc_hd__a31o_1
XFILLER_110_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3511__B _3746_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5037__A1 _4964_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5982_ _5982_/A _5982_/B _5982_/C VGND VGND VPWR VPWR _5982_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__3048__A0 _6041_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4796__B1 _4568_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4933_ _4922_/X _4925_/Y _4932_/Y _4563_/X VGND VGND VPWR VPWR _4934_/B sky130_fd_sc_hd__a22oi_1
XANTENNA__3599__B2 _3541_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3599__A1 _3579_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4864_ _4864_/A _4864_/B _4864_/C _4864_/D VGND VGND VPWR VPWR _4864_/Y sky130_fd_sc_hd__nand4_2
XANTENNA__4623__A _4623_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4548__B1 _4547_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4795_ _4668_/X _5829_/A _4793_/X _4794_/X VGND VGND VPWR VPWR _4795_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4012__A2 _3170_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3815_ _3815_/A _3815_/B _3815_/C _3975_/D VGND VGND VPWR VPWR _3816_/C sky130_fd_sc_hd__and4_1
XFILLER_20_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3746_ _3746_/A _3746_/B VGND VGND VPWR VPWR _3968_/C sky130_fd_sc_hd__nor2_2
XANTENNA__5760__A2 _5755_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3771__A1 _3759_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3771__B2 _3728_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5416_ input12/X _5395_/X _5405_/X VGND VGND VPWR VPWR _5416_/Y sky130_fd_sc_hd__a21oi_1
X_3677_ _3508_/X _3676_/Y _3539_/X VGND VGND VPWR VPWR _3677_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5454__A _5454_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput131 _2995_/X VGND VGND VPWR VPWR memory_imem_response_get[1] sky130_fd_sc_hd__buf_2
Xoutput120 _2993_/X VGND VGND VPWR VPWR memory_imem_response_get[0] sky130_fd_sc_hd__buf_2
Xoutput142 _3057_/X VGND VGND VPWR VPWR memory_imem_response_get[31] sky130_fd_sc_hd__buf_2
XANTENNA__5512__A2 _5504_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5347_ _5347_/A VGND VGND VPWR VPWR _6087_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4720__B1 _5805_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5278_ _6063_/Q _5570_/C VGND VGND VPWR VPWR _5279_/B sky130_fd_sc_hd__or2_1
XANTENNA__4079__A2 _4077_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4229_ _4716_/A _4513_/A input33/X _5044_/A _4228_/X VGND VGND VPWR VPWR _4229_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__3702__A _3773_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3287__B1 _3286_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3826__A2 _3638_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3039__A0 _6037_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5629__A _5629_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4533__A _4533_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4539__B1 _4538_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4003__A2 _3831_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3149__A _3165_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3211__B1 _3208_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6170__D _6170_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5200__B2 _5199_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5364__A _5364_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2988__A _6204_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3514__A1 _3632_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4711__B1 _4698_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input54_A memory_dmem_request_put[80] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5811__B _5811_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4708__A _4708_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3612__A _3871_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3817__A2 _3910_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5019__A1 _4931_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4443__A _4728_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3450__B1 _3340_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5990__A2 _5570_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5727__C1 _5163_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4580_ _4580_/A VGND VGND VPWR VPWR _5078_/A sky130_fd_sc_hd__clkbuf_4
X_3600_ _3600_/A VGND VGND VPWR VPWR _4073_/D sky130_fd_sc_hd__buf_2
XANTENNA__3059__A _3059_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput22 memory_dmem_request_put[48] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__clkbuf_1
Xinput11 memory_dmem_request_put[37] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__6080__D _6080_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3531_ _3509_/Y _3510_/X _3516_/Y _3517_/X _3530_/Y VGND VGND VPWR VPWR _3531_/X
+ sky130_fd_sc_hd__o221a_2
XANTENNA__3753__A1 _3622_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput44 memory_dmem_request_put[70] VGND VGND VPWR VPWR _4287_/B sky130_fd_sc_hd__clkbuf_4
Xinput33 memory_dmem_request_put[59] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_1
Xinput55 memory_dmem_request_put[81] VGND VGND VPWR VPWR _4218_/A sky130_fd_sc_hd__clkbuf_1
Xinput77 memory_imem_request_put[3] VGND VGND VPWR VPWR _3165_/A sky130_fd_sc_hd__clkbuf_4
Xinput66 memory_dmem_request_put[92] VGND VGND VPWR VPWR _4171_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__5274__A input5/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3462_ _3480_/A _3462_/B VGND VGND VPWR VPWR _3761_/A sky130_fd_sc_hd__nand2_4
XFILLER_6_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3393_ _3218_/X _3380_/X _3382_/X _3392_/Y _3692_/A VGND VGND VPWR VPWR _3393_/X
+ sky130_fd_sc_hd__a311o_1
X_6181_ _6196_/CLK _6181_/D VGND VGND VPWR VPWR _6181_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3505__A1 _3479_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5201_ input6/X _4200_/B VGND VGND VPWR VPWR _5201_/X sky130_fd_sc_hd__or2b_2
XFILLER_111_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5132_ _5129_/X _4991_/X _4241_/X _5131_/Y VGND VGND VPWR VPWR _5132_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_111_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5721__B _5721_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4618__A _4742_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5063_ _4350_/A _4725_/A _4697_/A _5005_/A VGND VGND VPWR VPWR _5063_/X sky130_fd_sc_hd__o211a_2
XANTENNA__3522__A _3522_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3808__A2 _3748_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4014_ _3343_/A _3475_/D _3499_/X _3350_/A VGND VGND VPWR VPWR _4014_/X sky130_fd_sc_hd__o31a_1
XFILLER_37_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5965_ _5746_/B _5963_/X _5964_/X _5734_/X VGND VGND VPWR VPWR _5965_/Y sky130_fd_sc_hd__a31oi_1
XANTENNA__5966__C1 _5965_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4353__A _4353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5896_ _4754_/X _5903_/A _5903_/D _5118_/D VGND VGND VPWR VPWR _5896_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4916_ _5013_/S _6138_/Q _4699_/X _5034_/B VGND VGND VPWR VPWR _4916_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4784__A3 _4910_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5981__A2 _5978_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4847_ _4843_/X _4833_/X _5102_/A _4846_/X _4420_/A VGND VGND VPWR VPWR _4847_/X
+ sky130_fd_sc_hd__o221a_2
XANTENNA__3607__B_N _3609_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4778_ _4778_/A VGND VGND VPWR VPWR _4778_/X sky130_fd_sc_hd__buf_2
XFILLER_119_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4941__B1 _4939_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3729_ _3715_/X _3726_/Y _3727_/X _6024_/Q _3728_/X VGND VGND VPWR VPWR _6024_/D
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4664__A_N _4645_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5497__A1 _5201_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5249__B2 _5248_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6009__C_N _5293_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4528__A _5073_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6165__D _6165_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2990__B _6205_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5421__A1 input13/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5957__C1 _5956_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5972__A2 _5062_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4263__A _4287_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3794__B1_N _3766_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5421__B2 _6105_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5078__B _5078_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4194__A_N _4225_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5185__B1 _5184_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5724__A2 _4390_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3196__C1 _3195_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4932__B1 _4930_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5488__B2 _5092_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4160__A1 _3815_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5822__A _5822_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4160__B2 _3510_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4438__A _4769_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4448__C1 _5020_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3342__A _3515_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4463__A2 _5744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5660__A1 _4369_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6075__D _6075_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3671__B1 _3670_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5948__C1 _5947_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5269__A _5286_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5963__A2 _4937_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4173__A _4301_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5750_ _6184_/Q _5646_/X _5729_/Y _5749_/Y VGND VGND VPWR VPWR _6184_/D sky130_fd_sc_hd__a2bb2oi_1
X_5681_ _5761_/C _5118_/C _4661_/X VGND VGND VPWR VPWR _5681_/Y sky130_fd_sc_hd__a21oi_2
X_4701_ _5016_/A _5191_/A VGND VGND VPWR VPWR _4702_/A sky130_fd_sc_hd__nand2_2
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3974__A1 _4048_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3974__B2 _3410_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4632_ _4716_/A _4513_/A input35/X _5044_/A _4631_/X VGND VGND VPWR VPWR _4632_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_30_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3726__A1 _3716_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4563_ _4563_/A VGND VGND VPWR VPWR _4563_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3726__B2 _3725_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3514_ _3632_/A _3983_/B _3600_/A VGND VGND VPWR VPWR _3653_/C sky130_fd_sc_hd__o21a_1
X_4494_ _5140_/C VGND VGND VPWR VPWR _4494_/X sky130_fd_sc_hd__buf_2
XANTENNA__3517__A _3748_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3445_ _3719_/B _3444_/X _3588_/B VGND VGND VPWR VPWR _3571_/C sky130_fd_sc_hd__o21a_2
XANTENNA__5479__A1 _4803_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5479__B2 _6119_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4151__A1 _3350_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5732__A _5732_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4634__A2_N _4630_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3376_ _3749_/B VGND VGND VPWR VPWR _3376_/X sky130_fd_sc_hd__clkbuf_8
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6164_ _6203_/CLK _6164_/D VGND VGND VPWR VPWR _6164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5115_ _4843_/A _4581_/C _5078_/A _5711_/A _4923_/A VGND VGND VPWR VPWR _5115_/Y
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA__4348__A _4759_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3252__A _3956_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ _6204_/CLK _6095_/D VGND VGND VPWR VPWR _6095_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5100__B1 _4642_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5046_ _5046_/A _5444_/A VGND VGND VPWR VPWR _5046_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4067__B _4067_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3662__B1 _3376_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5939__C1 _5938_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5179__A _5179_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4083__A _4083_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5948_ _6106_/Q _4807_/A _5905_/X _5947_/X VGND VGND VPWR VPWR _5948_/X sky130_fd_sc_hd__o211a_1
XFILLER_25_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4757__A3 _4725_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3965__A1 _3871_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5954__A2 _5944_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5879_ _5877_/X _4931_/X _5878_/Y _5782_/X VGND VGND VPWR VPWR _5879_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_21_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4811__A _4811_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4914__B1 _5822_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3427__A _3586_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4390__A1 _4243_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4127__D1 _4126_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4142__A1 _3406_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4142__B2 _3841_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5890__B2 _4459_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4258__A _4696_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3162__A _3162_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input17_A memory_dmem_request_put[43] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5642__A1 _4629_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4748__A3 _5711_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5945__A2 _4967_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3101__S _3105_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5158__B1 _5220_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4721__A _5263_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4440__B _4942_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5173__A3 _5102_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4905__B1 _4503_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6060__CLK _6207_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3982__D _4088_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3337__A _3621_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4920__A3 _4672_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output85_A _2991_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4133__A1 _4061_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3230_ _3882_/B VGND VGND VPWR VPWR _3230_/X sky130_fd_sc_hd__clkbuf_4
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5881__B2 _4305_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5881__A1 _5025_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3161_ _3161_/A VGND VGND VPWR VPWR _3161_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4168__A _4168_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3892__B1 _3464_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3239__A3 _3230_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3092_ _6188_/Q _6080_/Q _3094_/S VGND VGND VPWR VPWR _3093_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5094__C1 _5093_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3644__B1 _3499_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5802_ _5756_/X _5757_/X _5799_/Y _5801_/Y VGND VGND VPWR VPWR _5802_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3994_ _3614_/A _4149_/D _3525_/A _3711_/B _3648_/A VGND VGND VPWR VPWR _3994_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__5936__A2 _4917_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3947__A1 _4083_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5932__A2_N _5931_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5733_ _5955_/D _5733_/B _5813_/B VGND VGND VPWR VPWR _5733_/Y sky130_fd_sc_hd__nand3_1
X_5664_ _4644_/X _4642_/X _4961_/Y _4584_/X VGND VGND VPWR VPWR _5664_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5149__B1 _4744_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4615_ _4329_/X _4330_/X _4728_/A VGND VGND VPWR VPWR _4937_/B sky130_fd_sc_hd__o21ai_4
X_5595_ _5595_/A VGND VGND VPWR VPWR _6157_/D sky130_fd_sc_hd__clkbuf_1
X_4546_ _4854_/A VGND VGND VPWR VPWR _5118_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__3247__A _3311_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4477_ _4759_/A VGND VGND VPWR VPWR _4788_/B sky130_fd_sc_hd__buf_2
XFILLER_104_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3428_ _3902_/A VGND VGND VPWR VPWR _3428_/X sky130_fd_sc_hd__buf_2
XFILLER_100_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3359_ _3359_/A _3359_/B _3359_/C VGND VGND VPWR VPWR _3806_/B sky130_fd_sc_hd__and3_1
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input9_A memory_dmem_request_put[35] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6147_ _6147_/CLK _6147_/D VGND VGND VPWR VPWR _6147_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__5872__A1 input11/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3883__B1 _3762_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5085__C1 _5084_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6078_ _6176_/CLK _6078_/D VGND VGND VPWR VPWR _6078_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3710__A _3998_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5029_ _5029_/A VGND VGND VPWR VPWR _5029_/X sky130_fd_sc_hd__buf_2
XFILLER_66_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5927__A2 _5973_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4060__B1 _3868_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5637__A _5637_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6083__CLK _6202_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4541__A _4541_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4260__B _4264_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5155__A3 _5152_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4899__C1 _5182_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3157__A _3858_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4902__A3 _4898_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3705__A4 _3910_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5560__B1 _4976_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5372__A _5508_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4115__A1 _3680_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5863__A1 _4726_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3874__B1 _3512_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4418__A2 _5976_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3620__A _3781_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5311__S _5317_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output123_A _3020_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4716__A _4716_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5379__B1 _5378_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3929__A1 _3732_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5918__A2 _5167_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4051__B1 _3717_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5547__A _5988_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4170__B _4170_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4400_ _4442_/A VGND VGND VPWR VPWR _4533_/A sky130_fd_sc_hd__buf_2
XANTENNA__3067__A _3067_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5380_ _5376_/Y _5377_/Y _6098_/Q _5382_/B VGND VGND VPWR VPWR _5383_/A sky130_fd_sc_hd__a2bb2o_1
X_4331_ _4527_/C _4527_/D _4329_/X _4330_/X VGND VGND VPWR VPWR _4414_/A sky130_fd_sc_hd__o2bb2a_2
XFILLER_5_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4106__B2 _3932_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4262_ _4301_/D _4260_/Y _4261_/Y VGND VGND VPWR VPWR _4601_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__4106__A1 _3572_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3213_ _3442_/B _3440_/B VGND VGND VPWR VPWR _3746_/B sky130_fd_sc_hd__nand2b_4
XANTENNA__5854__A1 _4668_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_86_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6001_ _6207_/Q _6203_/Q VGND VGND VPWR VPWR _6009_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__3865__B1 _3522_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4193_ _5392_/C _4225_/A _4193_/C VGND VGND VPWR VPWR _4717_/A sky130_fd_sc_hd__and3b_1
XANTENNA__3006__S _3010_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3144_ _3311_/B VGND VGND VPWR VPWR _3437_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__4409__A2 _4405_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3075_ _6196_/Q _6072_/Q _3083_/S VGND VGND VPWR VPWR _3076_/A sky130_fd_sc_hd__mux2_2
XANTENNA__5082__A2 _5078_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4290__B1 _4259_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3977_ _3631_/X _3574_/X _3626_/X _3967_/X _3567_/X VGND VGND VPWR VPWR _3977_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4593__A1 _5008_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5716_ _5076_/X _4459_/X _5192_/X _4556_/X _4950_/A VGND VGND VPWR VPWR _5716_/X
+ sky130_fd_sc_hd__o41a_2
XFILLER_10_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5790__B1 _5774_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5647_ _5822_/A VGND VGND VPWR VPWR _5811_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5542__B1 _5491_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5578_ _5578_/A VGND VGND VPWR VPWR _6149_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4529_ _4578_/A _4734_/A VGND VGND VPWR VPWR _4661_/A sky130_fd_sc_hd__nand2_1
XFILLER_104_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4648__A2 _5971_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5845__A1 _4570_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3856__B1 _6032_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5058__C1 _5687_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3320__A2 _3814_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4536__A _4536_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3608__A0 _3756_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3440__A _3440_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5209__A2_N _5208_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4805__C1 _4804_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4820__A2 _4929_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6173__D _6173_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4033__B1 _4032_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4271__A _4811_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5230__C1 _5755_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5781__B1 _5780_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5367__A _6147_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5396__A1_N _6178_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5533__B1 _5504_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5306__S _5306_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4149__C _4152_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5049__C1 _4935_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4446__A _4585_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput9 memory_dmem_request_put[35] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_4
XFILLER_91_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5064__A2 _4350_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3350__A _3350_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3075__A1 _6072_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6083__D _6083_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4880_ _4671_/X _5944_/C _4878_/Y _5755_/C VGND VGND VPWR VPWR _4880_/Y sky130_fd_sc_hd__a31oi_4
X_3900_ _3859_/A _3653_/A _3643_/A VGND VGND VPWR VPWR _3900_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_60_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3831_ _3831_/A VGND VGND VPWR VPWR _3831_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4024__B1 _3302_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3762_ _3762_/A VGND VGND VPWR VPWR _3762_/X sky130_fd_sc_hd__buf_2
XANTENNA__5277__A _6063_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4181__A _4219_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3509__B _3589_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5501_ _5501_/A _5501_/B VGND VGND VPWR VPWR _5502_/A sky130_fd_sc_hd__and2_1
X_3693_ _3659_/D _3673_/B _3429_/X _3380_/X VGND VGND VPWR VPWR _3695_/C sky130_fd_sc_hd__o211a_1
XANTENNA__5524__B1 _5491_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5432_ _5432_/A VGND VGND VPWR VPWR _5433_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_114_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5363_ _6051_/Q _6095_/Q _5365_/S VGND VGND VPWR VPWR _5364_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3550__A2 _3592_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3525__A _3525_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4314_ _4405_/A _4341_/B _4518_/A VGND VGND VPWR VPWR _4699_/A sky130_fd_sc_hd__and3_2
XANTENNA__5827__A1 _5152_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5294_ _5294_/A input2/X _6013_/B VGND VGND VPWR VPWR _5294_/X sky130_fd_sc_hd__and3_1
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4245_ _4245_/A VGND VGND VPWR VPWR _4246_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_59_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4176_ _4217_/C _4217_/D VGND VGND VPWR VPWR _4230_/C sky130_fd_sc_hd__nor2_1
XANTENNA__4356__A _4369_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3853__A3 _3680_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3127_ _6052_/Q _6096_/Q _3127_/S VGND VGND VPWR VPWR _3128_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3260__A _3260_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5055__A2 _5720_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3058_ _6189_/Q _6065_/Q _3060_/S VGND VGND VPWR VPWR _3059_/A sky130_fd_sc_hd__mux2_2
XANTENNA__3066__A1 _6068_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6004__A1 _6203_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4015__B1 _3699_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5763__B1 _4948_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4522__C _5715_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4318__A1 _4293_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6121__CLK _6123_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5530__A3 _5529_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5818__A1 _5420_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6168__D _6168_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4266__A _4266_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3170__A _4004_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4006__B1 _3574_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4557__A1 _4457_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5097__A _5899_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4557__B2 _4556_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5754__B1 _4964_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6002__A1_N _3096_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5506__B1 _5388_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3345__A _3345_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5809__A1 _5045_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6078__D _6078_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4030_ _3376_/X _4026_/X _4029_/X _3562_/A VGND VGND VPWR VPWR _4030_/Y sky130_fd_sc_hd__a211oi_4
XFILLER_84_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5037__A2 _5019_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3080__A _3080_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4176__A _4217_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5981_ _5708_/Y _5978_/Y _5237_/X _5980_/Y _4767_/X VGND VGND VPWR VPWR _5982_/B
+ sky130_fd_sc_hd__o221ai_2
XFILLER_52_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3048__A1 _6173_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4796__A1 _4782_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4932_ _4927_/X _5680_/C _4930_/X _4931_/X VGND VGND VPWR VPWR _4932_/Y sky130_fd_sc_hd__o22ai_1
XANTENNA__3599__A2 _3598_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5993__B1 _5410_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4863_ _5745_/A _5034_/C _5240_/B _5079_/B _5721_/C VGND VGND VPWR VPWR _4863_/X
+ sky130_fd_sc_hd__o221a_2
XANTENNA__4548__A1 _5976_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4794_ _4819_/A VGND VGND VPWR VPWR _4794_/X sky130_fd_sc_hd__buf_6
X_3814_ _3814_/A VGND VGND VPWR VPWR _3975_/D sky130_fd_sc_hd__buf_2
XANTENNA__6144__CLK _6146_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5438__C _5438_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3745_ _4089_/A _3499_/X _3271_/A _3594_/X VGND VGND VPWR VPWR _3748_/C sky130_fd_sc_hd__o211a_1
XFILLER_118_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3771__A2 _3770_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3676_ _3139_/X _3671_/X _3672_/X _3675_/X VGND VGND VPWR VPWR _3676_/Y sky130_fd_sc_hd__a31oi_2
Xoutput110 _3065_/X VGND VGND VPWR VPWR memory_dmem_response_get[2] sky130_fd_sc_hd__buf_2
X_5415_ _5415_/A VGND VGND VPWR VPWR _6103_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3255__A _3461_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput121 _3016_/X VGND VGND VPWR VPWR memory_imem_response_get[10] sky130_fd_sc_hd__buf_2
Xoutput143 _2999_/X VGND VGND VPWR VPWR memory_imem_response_get[3] sky130_fd_sc_hd__buf_2
Xoutput132 _3038_/X VGND VGND VPWR VPWR memory_imem_response_get[20] sky130_fd_sc_hd__buf_2
XFILLER_99_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5346_ _6180_/Q _6087_/Q _5350_/S VGND VGND VPWR VPWR _5347_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4720__A1 _4716_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5277_ _6063_/Q _5570_/C VGND VGND VPWR VPWR _5285_/A sky130_fd_sc_hd__nand2_1
XANTENNA__4079__A3 _3223_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4228_ input9/X _4717_/A _4718_/A input17/X _4804_/A VGND VGND VPWR VPWR _4228_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4484__B1 _6136_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3287__A1 _3243_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4159_ _4124_/B _3844_/X _3910_/A _3553_/X _3717_/X VGND VGND VPWR VPWR _4159_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_28_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3039__A1 _6169_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3995__C1 _4073_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4539__A1 _5079_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5736__B1 _5735_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3211__A1 _4135_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3165__A _3165_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3514__A2 _3983_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4711__A1 _4345_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input47_A memory_dmem_request_put[73] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4475__B1 _4860_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4708__B _5152_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3612__B _4083_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6017__CLK _6155_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5019__A2 _5017_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5975__B1 _5735_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6167__CLK _6197_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4443__B _4860_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3450__A1 _4102_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5727__B1 _5403_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput12 memory_dmem_request_put[38] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__buf_2
X_3530_ _3521_/Y _3522_/X _3241_/X _3529_/X VGND VGND VPWR VPWR _3530_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__3753__A2 _3734_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput45 memory_dmem_request_put[71] VGND VGND VPWR VPWR _4405_/B sky130_fd_sc_hd__clkbuf_4
Xinput23 memory_dmem_request_put[49] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput34 memory_dmem_request_put[60] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput56 memory_dmem_request_put[82] VGND VGND VPWR VPWR _4219_/D sky130_fd_sc_hd__clkbuf_1
Xinput78 memory_imem_request_put[4] VGND VGND VPWR VPWR _3387_/B sky130_fd_sc_hd__buf_4
Xinput67 memory_dmem_request_put[93] VGND VGND VPWR VPWR _4171_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_115_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3461_ _3461_/A _3461_/B VGND VGND VPWR VPWR _3480_/A sky130_fd_sc_hd__or2_1
XFILLER_6_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3392_ _3919_/A _4083_/A _3893_/C _3749_/C _3860_/A VGND VGND VPWR VPWR _3392_/Y
+ sky130_fd_sc_hd__a311oi_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3505__A2 _3483_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4163__C1 _4162_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6180_ _6204_/CLK _6180_/D VGND VGND VPWR VPWR _6180_/Q sky130_fd_sc_hd__dfxtp_1
X_5200_ _6057_/Q _5040_/X _5166_/Y _5199_/Y VGND VGND VPWR VPWR _6057_/D sky130_fd_sc_hd__a2bb2oi_1
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5131_ _5131_/A _5444_/A VGND VGND VPWR VPWR _5131_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5721__C _5721_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5062_ _5062_/A VGND VGND VPWR VPWR _5062_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_111_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4013_ _3536_/X _3701_/X _3501_/Y _4036_/C _4012_/X VGND VGND VPWR VPWR _4013_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_65_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5964_ _5176_/X _5179_/X _5025_/Y _5753_/X VGND VGND VPWR VPWR _5964_/X sky130_fd_sc_hd__a31o_1
XFILLER_52_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5966__B1 _5940_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5895_ _4692_/X _4960_/X _5028_/X _4771_/X _5755_/C VGND VGND VPWR VPWR _5895_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4915_ _6051_/Q _4629_/X _4630_/X _4905_/X _4914_/X VGND VGND VPWR VPWR _6051_/D
+ sky130_fd_sc_hd__o32a_1
X_4846_ _4483_/X _4485_/X _5028_/A _5133_/A VGND VGND VPWR VPWR _4846_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5718__B1 _4924_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5194__A1 _4305_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4777_ _4777_/A VGND VGND VPWR VPWR _4777_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__4941__A1 _4422_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4941__B2 _4940_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3728_ _3822_/A VGND VGND VPWR VPWR _3728_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3659_ _4034_/A _3904_/B _3966_/C _3659_/D VGND VGND VPWR VPWR _3659_/X sky130_fd_sc_hd__or4_2
XANTENNA__4154__C1 _4044_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5497__A2 _5405_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5329_ _5329_/A VGND VGND VPWR VPWR _6079_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5654__C1 _4999_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3432__B _3432_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4544__A _5000_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2990__C _6179_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5421__A2 _5412_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5957__B1 _5905_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3213__A_N _3442_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5078__C _5687_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5709__B1 _4387_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6181__D _6181_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5185__A1 _5712_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2999__A _2999_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3196__B1 _3161_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4932__A1 _4927_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4932__B2 _4931_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4145__C1 _3868_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5893__C1 _5892_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4160__A2 _3673_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5822__B _5822_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3623__A _3959_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4448__B1 _5903_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5660__A2 _4574_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3671__A1 _3666_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4454__A _4640_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5948__B1 _5905_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5269__B input3/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4700_ _4700_/A VGND VGND VPWR VPWR _5016_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _5680_/A _5680_/B _5680_/C VGND VGND VPWR VPWR _5680_/X sky130_fd_sc_hd__and3_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3974__A2 _4065_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6091__D _6091_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4631_ input11/X _4717_/A _4718_/A input19/X _4804_/A VGND VGND VPWR VPWR _4631_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_30_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5285__A _5285_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4562_ _5903_/C VGND VGND VPWR VPWR _4563_/A sky130_fd_sc_hd__buf_6
XANTENNA__3726__A2 _3537_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3513_ _3513_/A VGND VGND VPWR VPWR _3600_/A sky130_fd_sc_hd__clkbuf_2
X_4493_ _4623_/A VGND VGND VPWR VPWR _5140_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_116_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3444_ _3802_/B _3437_/B _3895_/A _3591_/A VGND VGND VPWR VPWR _3444_/X sky130_fd_sc_hd__o2bb2a_2
XFILLER_89_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5479__A2 _5090_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5884__C1 _4618_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5732__B _5732_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3375_ _3589_/B VGND VGND VPWR VPWR _3749_/B sky130_fd_sc_hd__buf_2
XANTENNA__3533__A _3911_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4151__A2 _4105_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ _6197_/CLK _6163_/D VGND VGND VPWR VPWR _6163_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4629__A _4629_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5114_ _5101_/Y _5104_/X _4393_/X _5113_/Y VGND VGND VPWR VPWR _5127_/A sky130_fd_sc_hd__o211ai_2
XFILLER_57_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ _6204_/CLK _6094_/D VGND VGND VPWR VPWR _6094_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5100__A1 _5004_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3252__B _3687_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _5045_/A VGND VGND VPWR VPWR _5444_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3662__A1 _3658_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4364__A _4364_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5939__B1 _5937_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4083__B _4083_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5947_ input14/X _5395_/A _5163_/A _5093_/A VGND VGND VPWR VPWR _5947_/X sky130_fd_sc_hd__a211o_1
XFILLER_13_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3965__A2 _3457_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5954__A3 _5148_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5878_ _5878_/A _5878_/B _5878_/C _5971_/B VGND VGND VPWR VPWR _5878_/Y sky130_fd_sc_hd__nand4_4
XFILLER_21_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4829_ _4878_/B _4551_/A _4864_/B VGND VGND VPWR VPWR _4829_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__3708__A _3708_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4914__A1 _4908_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4914__B2 _4913_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4390__A2 _4985_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4127__C1 _3685_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4678__B1 _4643_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4142__A2 _4073_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6176__D _6176_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5642__A2 _4630_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5158__A1 _5141_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3618__A _3643_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5309__S _5317_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6205__CLK _6205_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4440__C _4551_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4905__A1 _4767_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4669__B1 _4668_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4133__A2 _3904_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3353__A _3353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5881__A2 _5880_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3160_ _3673_/A VGND VGND VPWR VPWR _3161_/A sky130_fd_sc_hd__buf_2
XANTENNA__4168__B _4168_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3892__A1 _3829_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3091_ _3091_/A VGND VGND VPWR VPWR _3091_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__6086__D _6086_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5094__B1 _5092_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3644__B2 _3543_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3644__A1 _3633_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4841__B1 _5746_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4184__A _4301_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5801_ _5800_/X _4762_/Y _5145_/X VGND VGND VPWR VPWR _5801_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_35_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3993_ _3748_/A _3988_/Y _3989_/X _3562_/A _3992_/X VGND VGND VPWR VPWR _4002_/B
+ sky130_fd_sc_hd__o311a_1
X_5732_ _5732_/A _5732_/B _5973_/C VGND VGND VPWR VPWR _5813_/B sky130_fd_sc_hd__nand3_1
XANTENNA__3947__A2 _3975_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4912__A _5924_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5149__A1 _5147_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3528__A _3528_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5663_ _5657_/Y _5662_/Y _5175_/A VGND VGND VPWR VPWR _5674_/A sky130_fd_sc_hd__a21o_1
X_4614_ _4614_/A VGND VGND VPWR VPWR _4707_/D sky130_fd_sc_hd__clkbuf_4
X_5594_ _6157_/Q _6025_/Q _5594_/S VGND VGND VPWR VPWR _5595_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4545_ _5073_/A VGND VGND VPWR VPWR _5971_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__3247__B _3461_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5743__A _5743_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4476_ _5170_/A VGND VGND VPWR VPWR _5711_/A sky130_fd_sc_hd__clkbuf_4
X_3427_ _3586_/A VGND VGND VPWR VPWR _3902_/A sky130_fd_sc_hd__buf_2
XANTENNA__4359__A _4878_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3263__A _3468_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6146_ _6146_/CLK _6146_/D VGND VGND VPWR VPWR _6146_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ _3287_/X _3290_/X _3356_/Y _6017_/Q _3357_/X VGND VGND VPWR VPWR _6017_/D
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5872__A2 _5420_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3883__A1 _4149_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3883__B2 _3710_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5085__B1 _5220_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6077_ _6203_/CLK _6077_/D VGND VGND VPWR VPWR _6077_/Q sky130_fd_sc_hd__dfxtp_1
X_3289_ _3786_/A VGND VGND VPWR VPWR _4103_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5028_ _5028_/A VGND VGND VPWR VPWR _5028_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3635__A1 _4124_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3710__B _3719_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4596__C1 _4595_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3399__B1 _3653_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5927__A3 _4839_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4060__A1 _3335_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3438__A _3756_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5155__A4 _4582_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4899__B1 _4815_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3157__B _3278_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5560__A1 _5437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5848__C1 _5769_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4115__A2 _4073_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5863__A2 _5070_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3874__A1 _3410_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3620__B _4034_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3112__S _3116_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output116_A _3073_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5379__A1 _5376_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4732__A _4732_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3929__A2 _3926_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4051__A1 _3536_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5547__B _5547_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4339__C1 _5179_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3348__A _3687_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5563__A _5563_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4330_ _4602_/A VGND VGND VPWR VPWR _4330_/X sky130_fd_sc_hd__buf_2
XFILLER_99_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4261_ _6133_/Q VGND VGND VPWR VPWR _4261_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5839__C1 _5175_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4106__A2 _3797_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4179__A _4218_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5854__A2 _4296_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3212_ _3513_/A VGND VGND VPWR VPWR _4034_/A sky130_fd_sc_hd__buf_2
XFILLER_86_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3314__B1 _3767_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6000_ _6000_/A VGND VGND VPWR VPWR _6201_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3865__A1 _4039_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3865__B2 _3975_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4192_ _5438_/D input7/X VGND VGND VPWR VPWR _4193_/C sky130_fd_sc_hd__nor2_1
X_3143_ _3226_/A VGND VGND VPWR VPWR _3311_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4814__B1 _4780_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3074_ _3096_/A VGND VGND VPWR VPWR _3083_/S sky130_fd_sc_hd__buf_2
XANTENNA__5082__A3 _5079_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4290__A1 _5211_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4642__A _4642_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3976_ _3701_/X _3340_/X _4128_/B _3975_/Y _3838_/X VGND VGND VPWR VPWR _3976_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__4593__A2 _5009_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5715_ _5715_/A _5715_/B _5968_/B VGND VGND VPWR VPWR _5715_/X sky130_fd_sc_hd__and3_1
XFILLER_109_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3258__A _3344_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5646_ _5646_/A VGND VGND VPWR VPWR _5646_/X sky130_fd_sc_hd__buf_2
XANTENNA__5790__B2 _5789_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5542__B2 _6139_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5542__A1 _5523_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5577_ _6149_/Q _6016_/Q _5583_/S VGND VGND VPWR VPWR _5578_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4528_ _5073_/A VGND VGND VPWR VPWR _5687_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_2_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4459_ _4459_/A VGND VGND VPWR VPWR _4459_/X sky130_fd_sc_hd__buf_2
XANTENNA__4089__A _4089_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4648__A3 _4917_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5845__A2 _4571_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3856__B2 _3822_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3856__A1 _3840_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5058__B1 _5079_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6129_ _6145_/CLK _6129_/D VGND VGND VPWR VPWR _6129_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3608__A1 _3779_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3440__B _3440_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6050__CLK _6196_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4805__B1 _4718_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4552__A _4815_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5230__B1 _4487_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4033__A1 _4018_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5781__A1 _4924_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5367__B _6146_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3168__A _3632_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5533__A1 _4801_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5533__B2 _4254_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input77_A memory_imem_request_put[3] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5383__A _5383_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4741__C1 _4604_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3615__B _3680_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4149__D _4149_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4727__A _5188_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5049__B1 _5048_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3631__A _3631_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5322__S _5328_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5064__A3 _4852_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5558__A _5988_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4462__A _4462_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3830_ _3829_/X _3654_/X _3830_/C _3830_/D VGND VGND VPWR VPWR _3830_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__4024__A1 _4021_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5221__B1 _5206_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3761_ _3761_/A VGND VGND VPWR VPWR _3762_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5277__B _5570_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4181__B _4219_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3783__B1 _3537_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3078__A _3078_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5500_ _5495_/X _4229_/X _5498_/X _6125_/Q _5499_/X VGND VGND VPWR VPWR _5501_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3692_ _3692_/A VGND VGND VPWR VPWR _3695_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__4980__C1 _4979_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5524__A1 _5523_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5524__B2 _6133_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5431_ _5431_/A _5431_/B VGND VGND VPWR VPWR _5968_/A sky130_fd_sc_hd__nand2_1
XANTENNA__3535__B1 _3534_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3806__A _3806_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5362_ _5362_/A VGND VGND VPWR VPWR _6094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4313_ _4313_/A VGND VGND VPWR VPWR _4518_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5827__A2 _5971_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3017__S _3021_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5293_ _6206_/Q _6204_/Q input2/X VGND VGND VPWR VPWR _5293_/X sky130_fd_sc_hd__and3b_1
XFILLER_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4244_ _4244_/A VGND VGND VPWR VPWR _4246_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_19_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4637__A _5191_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6073__CLK _6074_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3541__A _3891_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4175_ _4217_/A _4217_/B VGND VGND VPWR VPWR _4230_/B sky130_fd_sc_hd__nor2_1
X_3126_ _3126_/A VGND VGND VPWR VPWR _3126_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5055__A3 _4541_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3057_ _3057_/A VGND VGND VPWR VPWR _3057_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4015__A1 _3968_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4372__A _4415_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6004__A2 _5293_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5468__A _5468_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5212__B1 _5179_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5763__A1 _5190_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3959_ _3955_/X _3959_/B _4146_/A _3959_/D VGND VGND VPWR VPWR _3959_/X sky130_fd_sc_hd__and4b_1
XANTENNA__3774__B1 _3633_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4318__A2 _4246_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5629_ _5629_/A VGND VGND VPWR VPWR _5638_/S sky130_fd_sc_hd__buf_2
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3451__A _3538_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3170__B _3648_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6184__D _6184_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4006__A1 _4135_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4282__A _4282_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4557__A2 _4548_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5754__A1 _5752_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3765__B1 _3749_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5506__A1 _6126_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3626__A _3841_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5317__S _5317_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6096__CLK _6204_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5809__A2 _5470_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4457__A _4890_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5255__A2_N _5040_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5037__A3 _5024_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6094__D _6094_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4176__B _4217_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5980_ _4836_/X _5213_/X _5959_/X _5979_/Y _5961_/X VGND VGND VPWR VPWR _5980_/Y
+ sky130_fd_sc_hd__a32oi_4
XFILLER_18_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4931_ _4931_/A VGND VGND VPWR VPWR _4931_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__4796__A2 _4790_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3599__A3 _3453_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5993__A1 _5998_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4862_ _4862_/A VGND VGND VPWR VPWR _5721_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_32_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4192__A _5438_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5288__A _5508_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5640__A_N _6099_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3813_ _3622_/X _3812_/Y _3242_/X VGND VGND VPWR VPWR _3816_/B sky130_fd_sc_hd__a21oi_2
XFILLER_32_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4548__A2 _5971_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4793_ _5903_/C VGND VGND VPWR VPWR _4793_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_60_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5438__D _5438_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3744_ _3744_/A _3744_/B VGND VGND VPWR VPWR _3744_/X sky130_fd_sc_hd__or2_1
X_3675_ _3673_/Y _3593_/X _3674_/X _3724_/B VGND VGND VPWR VPWR _3675_/X sky130_fd_sc_hd__o31a_1
XANTENNA__3771__A3 _3727_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3536__A _3536_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput100 _3104_/X VGND VGND VPWR VPWR memory_dmem_response_get[20] sky130_fd_sc_hd__buf_2
X_5414_ _5414_/A _5422_/B VGND VGND VPWR VPWR _5415_/A sky130_fd_sc_hd__and2_1
XANTENNA__3255__B _3272_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput122 _3018_/X VGND VGND VPWR VPWR memory_imem_response_get[11] sky130_fd_sc_hd__buf_2
Xoutput133 _3040_/X VGND VGND VPWR VPWR memory_imem_response_get[21] sky130_fd_sc_hd__buf_2
Xoutput111 _3126_/X VGND VGND VPWR VPWR memory_dmem_response_get[30] sky130_fd_sc_hd__buf_2
XFILLER_99_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput144 _3003_/X VGND VGND VPWR VPWR memory_imem_response_get[4] sky130_fd_sc_hd__buf_2
XANTENNA__4720__A2 _4513_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5345_ _5345_/A VGND VGND VPWR VPWR _6086_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5751__A _6185_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5276_ _5276_/A VGND VGND VPWR VPWR _6062_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5380__A1_N _5376_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4367__A _4895_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4227_ _4227_/A VGND VGND VPWR VPWR _4513_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5681__B1 _4661_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4484__A1 _4482_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3271__A _3271_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3287__A2 _3268_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4158_ _3558_/X _3716_/X _3868_/X _3628_/A VGND VGND VPWR VPWR _4158_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4089_ _4089_/A _4089_/B VGND VGND VPWR VPWR _4089_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3109_ _3109_/A VGND VGND VPWR VPWR _3109_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_55_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3995__B1 _3362_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4539__A2 _4534_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5736__A1 _5733_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3747__B1 _3593_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3211__A2 _3205_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3446__A _3603_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_2_3_0_CLK clkbuf_2_3_0_CLK/A VGND VGND VPWR VPWR clkbuf_3_7_0_CLK/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6179__D _6179_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4711__A2 _4691_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5661__A _5661_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4277__A _6134_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4475__A1 _4329_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3181__A _3330_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4708__C _4891_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3612__C _3680_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5672__B1 _5676_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5019__A3 _4870_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5424__B1 _5405_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5975__A1 _5715_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5975__B2 _5974_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3450__A2 _3426_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5727__A1 _5045_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5836__A _5836_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3738__B1 _3815_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput13 memory_dmem_request_put[39] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput24 memory_dmem_request_put[50] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_1
Xinput35 memory_dmem_request_put[61] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_1
Xinput46 memory_dmem_request_put[72] VGND VGND VPWR VPWR _4285_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_115_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput79 memory_imem_request_put[5] VGND VGND VPWR VPWR _3233_/A sky130_fd_sc_hd__clkbuf_4
Xinput57 memory_dmem_request_put[83] VGND VGND VPWR VPWR _4219_/C sky130_fd_sc_hd__clkbuf_1
Xinput68 memory_dmem_request_put[94] VGND VGND VPWR VPWR _4168_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_115_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3460_ _3663_/A _3876_/A _3468_/A VGND VGND VPWR VPWR _3460_/X sky130_fd_sc_hd__a21o_2
XFILLER_97_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3391_ _3647_/A VGND VGND VPWR VPWR _3860_/A sky130_fd_sc_hd__buf_4
XANTENNA__3505__A3 _3490_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4163__B1 _3828_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6089__D _6089_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5130_ input28/X _4978_/X _5042_/X input12/X VGND VGND VPWR VPWR _5131_/A sky130_fd_sc_hd__a22o_1
XANTENNA__5112__C1 _5111_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5061_ _5061_/A VGND VGND VPWR VPWR _5061_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5663__B1 _5175_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4012_ _3525_/X _3170_/X _3654_/X VGND VGND VPWR VPWR _4012_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__3091__A _3091_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5963_ _4431_/X _4937_/Y _4870_/X _4541_/X VGND VGND VPWR VPWR _5963_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5966__A1 _5734_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6111__CLK _6123_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3977__B1 _3967_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4914_ _4908_/X _4721_/X _5822_/A _4913_/X VGND VGND VPWR VPWR _4914_/X sky130_fd_sc_hd__o22a_1
XFILLER_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5894_ _5882_/Y _5886_/Y _5845_/X _5893_/X VGND VGND VPWR VPWR _5894_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__3030__S _3032_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5718__A1 _5761_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4845_ _4614_/A _4738_/B _4772_/A _4696_/A VGND VGND VPWR VPWR _5133_/A sky130_fd_sc_hd__a31o_1
XFILLER_33_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5132__A2_N _4991_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4776_ _4926_/A _4926_/C _4640_/A _4811_/A VGND VGND VPWR VPWR _4928_/A sky130_fd_sc_hd__o211ai_4
XANTENNA__4650__A _4855_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5194__A2 _5192_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5746__A _5746_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3729__B1 _6024_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3727_ _4103_/C VGND VGND VPWR VPWR _3727_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4941__A2 _4423_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3658_ _3621_/D _3773_/B _3583_/A _3657_/X VGND VGND VPWR VPWR _3658_/X sky130_fd_sc_hd__a31o_2
XANTENNA__4154__B1 _3802_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3589_ _3611_/A _3589_/B VGND VGND VPWR VPWR _4128_/A sky130_fd_sc_hd__or2_2
XANTENNA__5497__A3 _5224_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3901__B1 _3900_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5328_ _6187_/Q _6079_/Q _5328_/S VGND VGND VPWR VPWR _5329_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5481__A _5481_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5700__A2_N _5646_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5654__B1 _4621_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5259_ _5256_/X _2986_/C _5388_/A VGND VGND VPWR VPWR _6060_/D sky130_fd_sc_hd__a21oi_1
XFILLER_87_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3665__C1 _3744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5406__B1 _5405_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5957__A1 _6107_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4971__A2_N _4536_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4090__C1 _3218_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5421__A3 _5431_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5078__D _5078_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5709__A1 _4838_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5185__A2 _5181_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4560__A _5228_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3196__A1 _3178_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3176__A _3870_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4932__A2 _5680_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3607__C _3781_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4145__B1 _3910_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3904__A _3904_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5893__B1 _5889_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3623__B _3623_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4448__B2 _5079_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4448__A1 _4437_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output146_A _3007_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5645__B1 _5013_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6134__CLK _6146_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3671__A2 _3668_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5948__A1 _6106_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3974__A3 _3553_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4470__A _4614_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5566__A _5566_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4908__C1 _4907_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4630_ _4630_/A VGND VGND VPWR VPWR _4630_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4384__B1 _4815_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5285__B _5285_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4561_ _4340_/Y _5818_/S _4341_/Y _4432_/A VGND VGND VPWR VPWR _5903_/C sky130_fd_sc_hd__o211a_1
XFILLER_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4492_ _4474_/X _4480_/X _4665_/A _4491_/X VGND VGND VPWR VPWR _4492_/X sky130_fd_sc_hd__o211a_1
X_3512_ _3512_/A VGND VGND VPWR VPWR _3512_/X sky130_fd_sc_hd__buf_2
XFILLER_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3443_ _3461_/B _3443_/B VGND VGND VPWR VPWR _3591_/A sky130_fd_sc_hd__and2b_1
XANTENNA__4136__B1 _3161_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5479__A3 _5445_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5884__B1 _5829_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5732__C _5973_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3814__A _3814_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6162_ _6197_/CLK _6162_/D VGND VGND VPWR VPWR _6162_/Q sky130_fd_sc_hd__dfxtp_1
X_5113_ _4836_/X _5105_/X _5108_/X _4746_/A _5112_/Y VGND VGND VPWR VPWR _5113_/Y
+ sky130_fd_sc_hd__o311ai_2
X_3374_ _3572_/A _4073_/A _4152_/A _3797_/A VGND VGND VPWR VPWR _3374_/X sky130_fd_sc_hd__a31o_2
XFILLER_69_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4151__A3 _4149_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5636__A0 _6176_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6093_ _6204_/CLK _6093_/D VGND VGND VPWR VPWR _6093_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5100__A2 _4675_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5044_/A VGND VGND VPWR VPWR _5045_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3662__A2 _3661_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5939__A1 _4679_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5946_ _5693_/Y _5943_/X _5945_/X VGND VGND VPWR VPWR _5946_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4083__C _4083_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5877_ _5976_/C _5008_/X _5009_/X _4360_/X VGND VGND VPWR VPWR _5877_/X sky130_fd_sc_hd__a31o_1
XFILLER_40_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4380__A _4462_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4828_ _5016_/A VGND VGND VPWR VPWR _4843_/B sky130_fd_sc_hd__buf_2
XANTENNA__5476__A _5476_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5086__A2_N _5040_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4759_ _4759_/A _4860_/A _4759_/C VGND VGND VPWR VPWR _4876_/A sky130_fd_sc_hd__nand3_1
XANTENNA__4914__A2 _4721_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4390__A3 _4986_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4127__B1 _4124_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4678__A1 _4421_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5875__B1 _5874_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3724__A _3724_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6157__CLK _6197_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3443__B _3443_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3886__C1 _3574_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5627__A0 _6172_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4555__A _5061_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6192__D _6192_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5039__A2_N _6053_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3810__C1 _3809_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5158__A2 _5142_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4366__B1 _4601_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4905__A2 _4868_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4440__D _5211_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4118__B1 _3374_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5866__B1 _4924_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4669__A1 _5140_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4669__B2 _4431_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3877__C1 _3350_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4133__A3 _4128_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3892__A2 _3720_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3090_ _6187_/Q _6079_/Q _3094_/S VGND VGND VPWR VPWR _3091_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5094__A1 _5090_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3644__A2 _3711_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4841__A1 _4838_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4841__B2 _4739_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5794__A1_N _4786_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3992_ _3992_/A _3992_/B _3992_/C VGND VGND VPWR VPWR _3992_/X sky130_fd_sc_hd__or3_1
X_5800_ _4317_/A _4363_/A _4488_/X _5240_/D _4255_/Y VGND VGND VPWR VPWR _5800_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5731_ _5731_/A _5731_/B VGND VGND VPWR VPWR _5732_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5296__A _5352_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5149__A2 _5148_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5662_ _5060_/X _5658_/Y _5031_/X _5661_/Y VGND VGND VPWR VPWR _5662_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_30_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4613_ _5746_/D _4610_/X _4612_/X _4345_/A VGND VGND VPWR VPWR _4613_/X sky130_fd_sc_hd__a31o_1
X_5593_ _5593_/A VGND VGND VPWR VPWR _6156_/D sky130_fd_sc_hd__clkbuf_1
X_4544_ _5000_/A VGND VGND VPWR VPWR _5976_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_116_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5743__B _5743_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4109__B1 _4108_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4475_ _4329_/X _4330_/X _4860_/C VGND VGND VPWR VPWR _5170_/A sky130_fd_sc_hd__o21ai_1
XFILLER_104_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3544__A _3780_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5857__B1 _5856_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3426_ _3522_/A _3425_/X _3673_/A VGND VGND VPWR VPWR _3426_/X sky130_fd_sc_hd__o21a_2
XFILLER_97_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6145_ _6145_/CLK _6145_/D VGND VGND VPWR VPWR _6145_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3357_ _3891_/A VGND VGND VPWR VPWR _3357_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3883__A2 _3520_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6176_/CLK _6076_/D VGND VGND VPWR VPWR _6076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5027_ _5971_/D _5025_/Y _4739_/X _5026_/X _5782_/A VGND VGND VPWR VPWR _5027_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_73_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5085__A1 _5057_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3288_ _3918_/A _3918_/C _3918_/B VGND VGND VPWR VPWR _3786_/A sky130_fd_sc_hd__nor3_1
XANTENNA__4375__A _4811_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3635__A2 _3634_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3710__C _3710_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4045__C1 _4044_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4596__B1 _4584_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3399__A1 _3841_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5793__C1 _5118_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3719__A _3998_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4060__A2 _3847_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5929_ _5235_/X _4967_/X _5928_/Y _5145_/X VGND VGND VPWR VPWR _5929_/Y sky130_fd_sc_hd__a22oi_2
XANTENNA__3438__B _3438_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4899__A1 _4878_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3157__C _3157_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5560__A2 _5439_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5848__B1 _5847_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4115__A3 _4111_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5863__A3 _4742_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6187__D _6187_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3874__A2 _3254_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input22_A memory_dmem_request_put[48] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4285__A _4301_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5379__A2 _5377_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output109_A _3124_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3929__A3 _3781_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4732__B _4732_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3629__A _3687_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4051__A2 _3844_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4339__B1 _4328_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3547__D1 _3546_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output90_A _3084_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3364__A _4034_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5839__B1 _5838_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4106__A3 _3911_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4260_ _4268_/A _4264_/C VGND VGND VPWR VPWR _4260_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4179__B _4218_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5854__A3 _4960_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3314__A1 _3867_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3211_ _4135_/B _3205_/X _3208_/X _3692_/A VGND VGND VPWR VPWR _3211_/X sky130_fd_sc_hd__o211a_1
X_4191_ input8/X VGND VGND VPWR VPWR _4225_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__6097__D _6097_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3142_ _3695_/B VGND VGND VPWR VPWR _3142_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3865__A2 _3799_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4814__A1 _4864_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4195__A _4195_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3073_ _3073_/A VGND VGND VPWR VPWR _3073_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4923__A _4923_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4290__A2 _4815_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4027__C1 _3659_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3975_ _3975_/A _3975_/B _3975_/C _3975_/D VGND VGND VPWR VPWR _3975_/Y sky130_fd_sc_hd__nand4_1
X_5714_ _4570_/Y _4571_/X _5705_/Y _5713_/X VGND VGND VPWR VPWR _5725_/A sky130_fd_sc_hd__o22ai_1
X_5645_ _6180_/Q _5166_/A _5013_/X _5644_/X VGND VGND VPWR VPWR _6180_/D sky130_fd_sc_hd__a22o_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3002__A0 _6020_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5542__A2 _5757_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5576_ _5576_/A VGND VGND VPWR VPWR _6148_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4750__B1 _4864_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4527_ _4527_/A _4536_/A _4527_/C _4527_/D VGND VGND VPWR VPWR _5073_/A sky130_fd_sc_hd__nand4_4
XANTENNA__3274__A _4152_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4458_ _4533_/A _5008_/A _5009_/A VGND VGND VPWR VPWR _4459_/A sky130_fd_sc_hd__and3_4
XANTENNA__4089__B _4089_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3409_ _3648_/A VGND VGND VPWR VPWR _3410_/A sky130_fd_sc_hd__buf_2
XANTENNA__4502__B1 _4224_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4389_ _4361_/X _4370_/X _4388_/X VGND VGND VPWR VPWR _4389_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_58_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6128_ _6147_/CLK _6128_/D VGND VGND VPWR VPWR _6128_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3856__A2 _3855_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5058__A1 _5096_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4805__A1 input14/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6059_ _6207_/CLK _6059_/D VGND VGND VPWR VPWR _6059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4805__B2 input22/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6007__B1 _5410_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4018__C1 _3580_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5230__A1 _4353_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4569__B1 _4568_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5766__C1 _5725_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4033__A2 _4024_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5230__B2 _5167_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5781__A2 _5063_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5367__C _6145_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5533__A2 _4482_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5383__B _5383_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3184__A _3443_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4741__B1 _5016_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3615__C _3871_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5603__S _5605_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5049__A1 _4552_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3123__S _3127_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4009__C1 _3577_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5558__B _5558_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4024__A2 _4023_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3359__A _3359_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3760_ _3881_/A VGND VGND VPWR VPWR _3760_/X sky130_fd_sc_hd__buf_2
XFILLER_20_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5221__B2 _5220_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3783__A1 _3157_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4980__B1 _4977_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3691_ _3684_/X _3690_/Y _3624_/X VGND VGND VPWR VPWR _3691_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5574__A _5618_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5430_ _5430_/A VGND VGND VPWR VPWR _6107_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5524__A2 _4287_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3535__A1 _3830_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3535__B2 _3830_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3806__B _3806_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5361_ _6050_/Q _6094_/Q _5361_/S VGND VGND VPWR VPWR _5362_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5293__B _6204_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4312_ _4482_/A _4308_/X _4986_/A _6138_/Q VGND VGND VPWR VPWR _4421_/A sky130_fd_sc_hd__o31a_2
X_5292_ _6204_/Q VGND VGND VPWR VPWR _5292_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4243_ _4243_/A VGND VGND VPWR VPWR _4243_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_101_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4918__A _4918_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3822__A _3822_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4174_ _4174_/A _4174_/B VGND VGND VPWR VPWR _4230_/A sky130_fd_sc_hd__nor2_2
X_3125_ _6051_/Q _6095_/Q _3127_/S VGND VGND VPWR VPWR _3126_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3056_ _6045_/Q _6177_/Q _3056_/S VGND VGND VPWR VPWR _3057_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5996__C1 _5388_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3471__B1 _3470_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5212__A1 _5211_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4015__A2 _4014_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5468__B _5468_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5212__B2 _5106_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3269__A _3904_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3958_ _3679_/X _4124_/B _3205_/X _3543_/Y _3992_/B VGND VGND VPWR VPWR _3959_/B
+ sky130_fd_sc_hd__o41ai_2
XANTENNA__5763__A2 _5761_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3774__A1 _3549_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4971__B1 _4404_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3623__D_N _3622_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5484__A _5484_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3889_ _3881_/Y _3888_/X _3624_/X _3787_/X VGND VGND VPWR VPWR _3889_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4318__A3 _4246_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5628_ _5628_/A VGND VGND VPWR VPWR _6172_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5559_ _5559_/A VGND VGND VPWR VPWR _6144_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4723__B1 _4189_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4828__A _5016_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3732__A _4034_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3170__C _4065_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4563__A _4563_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4006__A2 _3814_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3179__A _3443_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5754__A2 _5753_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3765__A1 _3867_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4962__B1 _4856_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5394__A _5420_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5506__A2 _5504_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4714__B1 _4634_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_CLK CLK VGND VGND VPWR VPWR clkbuf_0_CLK/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__3642__A _3642_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4738__A _4738_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5333__S _5339_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5978__C1 _5977_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5569__A _5569_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4473__A _4926_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4930_ _5098_/A VGND VGND VPWR VPWR _4930_/X sky130_fd_sc_hd__buf_2
XANTENNA__4796__A3 _4795_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5993__A2 _5571_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4861_ _4936_/A VGND VGND VPWR VPWR _5079_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__4192__B input7/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3812_ _3238_/X _3426_/X _3862_/A VGND VGND VPWR VPWR _3812_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3089__A _3089_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4792_ _4792_/A VGND VGND VPWR VPWR _5829_/A sky130_fd_sc_hd__buf_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3743_ _3734_/Y _3738_/Y _3742_/X _3688_/X VGND VGND VPWR VPWR _3744_/B sky130_fd_sc_hd__o2bb2a_1
X_3674_ _3767_/D _3674_/B _3674_/C VGND VGND VPWR VPWR _3674_/X sky130_fd_sc_hd__and3_2
XFILLER_9_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput101 _3106_/X VGND VGND VPWR VPWR memory_dmem_response_get[21] sky130_fd_sc_hd__buf_2
XANTENNA__6040__CLK _6202_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5413_ input11/X _5412_/X _5395_/X _5398_/X _6103_/Q VGND VGND VPWR VPWR _5414_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_99_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput123 _3020_/X VGND VGND VPWR VPWR memory_imem_response_get[12] sky130_fd_sc_hd__buf_2
Xoutput134 _3042_/X VGND VGND VPWR VPWR memory_imem_response_get[23] sky130_fd_sc_hd__buf_2
Xoutput112 _3128_/X VGND VGND VPWR VPWR memory_dmem_response_get[31] sky130_fd_sc_hd__buf_2
XANTENNA__3028__S _3032_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5344_ _6058_/Q _6086_/Q _5350_/S VGND VGND VPWR VPWR _5345_/A sky130_fd_sc_hd__mux2_1
Xoutput145 _3005_/X VGND VGND VPWR VPWR memory_imem_response_get[5] sky130_fd_sc_hd__buf_2
XANTENNA__4720__A3 input37/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5275_ _5275_/A _5275_/B _6014_/B VGND VGND VPWR VPWR _5276_/A sky130_fd_sc_hd__and3_1
XFILLER_101_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4226_ _5438_/C VGND VGND VPWR VPWR _4716_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5130__B1 _5042_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6190__CLK _6205_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5681__A1 _5761_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4484__A2 _4308_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3287__A3 _3284_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4157_ _4148_/X _3477_/X _4088_/C _4156_/Y VGND VGND VPWR VPWR _4157_/X sky130_fd_sc_hd__a211o_1
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3108_ _6180_/Q _6087_/Q _3116_/S VGND VGND VPWR VPWR _3109_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3996__A1_N _3645_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4088_ _3839_/X _4088_/B _4088_/C _4088_/D VGND VGND VPWR VPWR _4088_/X sky130_fd_sc_hd__and4b_1
XANTENNA__4383__A _4734_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3444__B1 _3895_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3039_ _6037_/Q _6169_/Q _3043_/S VGND VGND VPWR VPWR _3040_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3995__A1 _3406_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5197__B1 _4685_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3747__A1 _3299_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5736__A2 _5734_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4944__B1 _4618_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3727__A _4103_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3446__B _3446_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4711__A3 _4694_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3462__A _3480_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5661__B _5661_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5121__B1 _5120_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4475__A2 _4330_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4708__D _4708_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6195__D _6195_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5672__A1 _4633_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3683__B1 _3649_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3612__D _3612_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5424__A1 input14/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3435__B1 _3345_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4293__A _4293_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5975__A2 _4390_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4632__C1 _4631_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3450__A3 _3431_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5727__A2 _5455_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5836__B _5836_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3738__A1 _3736_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6063__CLK _6201_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5328__S _5328_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput14 memory_dmem_request_put[40] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_4
Xinput25 memory_dmem_request_put[51] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_1
Xinput36 memory_dmem_request_put[62] VGND VGND VPWR VPWR input36/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__6013__A _6207_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput47 memory_dmem_request_put[73] VGND VGND VPWR VPWR _4317_/A sky130_fd_sc_hd__buf_4
Xinput58 memory_dmem_request_put[84] VGND VGND VPWR VPWR _4217_/B sky130_fd_sc_hd__clkbuf_1
Xinput69 memory_dmem_request_put[95] VGND VGND VPWR VPWR _4168_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_115_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4163__A1 _3300_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3390_ _3522_/A VGND VGND VPWR VPWR _3749_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_111_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5112__B1 _4541_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3372__A _3956_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5060_ _4668_/A _5000_/A _5118_/B _4675_/A VGND VGND VPWR VPWR _5060_/X sky130_fd_sc_hd__o31a_2
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5663__A1 _5657_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4011_ _4002_/X _4010_/Y _3821_/X _6038_/Q _3822_/X VGND VGND VPWR VPWR _6038_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4871__C1 _5078_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3426__B1 _3673_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5962_ _5959_/X _5661_/A _5960_/X _5961_/X VGND VGND VPWR VPWR _5962_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5299__A _5299_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3977__A1 _3631_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5966__A2 _5962_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4913_ _6131_/Q _4975_/A _4224_/A VGND VGND VPWR VPWR _4913_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3977__B2 _3567_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5893_ _5756_/X _5757_/X _5889_/X _5892_/X VGND VGND VPWR VPWR _5893_/X sky130_fd_sc_hd__a211o_1
X_4844_ _4878_/C _4878_/D _4649_/A VGND VGND VPWR VPWR _5028_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__5718__A2 _4996_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4931__A _4931_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4650__B _5899_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4775_ _4692_/A _4864_/C _4937_/A _4259_/A _4673_/B VGND VGND VPWR VPWR _4967_/A
+ sky130_fd_sc_hd__o2111ai_4
XANTENNA__5746__B _5746_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3729__A1 _3715_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3729__B2 _3728_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3726_ _3716_/X _3537_/X _3142_/X _3725_/X _3302_/X VGND VGND VPWR VPWR _3726_/Y
+ sky130_fd_sc_hd__o221ai_4
X_3657_ _3657_/A _3657_/B _3657_/C VGND VGND VPWR VPWR _3657_/X sky130_fd_sc_hd__and3_1
X_3588_ _3594_/A _3588_/B _3588_/C VGND VGND VPWR VPWR _3588_/X sky130_fd_sc_hd__and3_2
XANTENNA__4154__B2 _4153_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4154__A1 _3674_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4378__A _4378_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3901__A1 _3834_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5327_ _5327_/A VGND VGND VPWR VPWR _6078_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5103__B1 _4757_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3282__A _3282_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5654__A1 _4369_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5258_ _5545_/A VGND VGND VPWR VPWR _5388_/A sky130_fd_sc_hd__buf_4
XFILLER_29_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5189_ _4374_/X _4378_/Y _5706_/B _4582_/X VGND VGND VPWR VPWR _5189_/X sky130_fd_sc_hd__a31o_1
XFILLER_68_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4209_ _4209_/A VGND VGND VPWR VPWR _5818_/S sky130_fd_sc_hd__buf_2
XANTENNA__3665__B1 _3664_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5406__A1 input10/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5957__A2 _4241_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4090__B1 _3482_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6086__CLK _6203_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5709__A2 _5029_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5185__A3 _5183_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3457__A _3457_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3196__A2 _3183_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5590__A0 _6155_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3607__D _3781_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4145__A1 _3460_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4145__B2 _3875_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5342__A0 _6057_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4288__A _4527_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3904__B _3904_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5893__A1 _5756_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input52_A memory_dmem_request_put[78] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3623__C _3623_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3192__A _3343_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4448__A2 _4440_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5645__A1 _6180_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5645__B2 _5644_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4853__C1 _4585_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output139_A _3053_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3671__A3 _3910_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4605__C1 _4604_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3408__B1 _3401_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5948__A2 _4807_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4081__B1 _6041_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4103__B_N _4096_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4908__B1 _5805_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4384__A1 _4878_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4560_ _5228_/A VGND VGND VPWR VPWR _4746_/A sky130_fd_sc_hd__buf_4
XANTENNA__3367__A _3582_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5030__C1 _5029_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5581__A0 _6151_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4491_ _4487_/Y _4488_/X _4843_/C _5240_/C VGND VGND VPWR VPWR _4491_/X sky130_fd_sc_hd__a31o_1
X_3511_ _3841_/A _3746_/A VGND VGND VPWR VPWR _3512_/A sky130_fd_sc_hd__nand2_4
XFILLER_6_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5582__A _5582_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3442_ _3272_/A _3442_/B VGND VGND VPWR VPWR _3895_/A sky130_fd_sc_hd__and2b_2
XANTENNA__4136__B2 _4061_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4136__A1 _3536_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5333__A0 _6053_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5884__A1 _5878_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5884__B2 _5878_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3373_ _3966_/B VGND VGND VPWR VPWR _4152_/A sky130_fd_sc_hd__clkbuf_2
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4198__A _4515_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6161_ _6201_/CLK _6161_/D VGND VGND VPWR VPWR _6161_/Q sky130_fd_sc_hd__dfxtp_1
X_5112_ _5109_/Y _5110_/Y _4541_/X _5111_/X VGND VGND VPWR VPWR _5112_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_97_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5636__A1 _6044_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6092_ _6204_/CLK _6092_/D VGND VGND VPWR VPWR _6092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5100__A3 _5080_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_85_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4926__A _4926_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ input26/X _4978_/X _5042_/X input10/X VGND VGND VPWR VPWR _5046_/A sky130_fd_sc_hd__a22o_1
Xclkbuf_2_2_0_CLK clkbuf_2_3_0_CLK/A VGND VGND VPWR VPWR clkbuf_3_5_0_CLK/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5939__A2 _5935_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3041__S _3043_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5945_ _4679_/X _4967_/X _5944_/Y _4657_/A _4964_/A VGND VGND VPWR VPWR _5945_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4072__B1 _3624_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4661__A _4661_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5757__A _5757_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5876_ _6191_/Q _4715_/X _5858_/Y _5875_/Y VGND VGND VPWR VPWR _6191_/D sky130_fd_sc_hd__a2bb2oi_1
X_4827_ _4827_/A VGND VGND VPWR VPWR _5102_/A sky130_fd_sc_hd__buf_4
XANTENNA__3277__A _3500_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4758_ _4955_/A VGND VGND VPWR VPWR _5152_/B sky130_fd_sc_hd__buf_4
XANTENNA__5572__B1 _5570_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4689_ _5191_/A VGND VGND VPWR VPWR _5745_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_107_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3709_ _4074_/B _3157_/C _3911_/B _4065_/B _4105_/B VGND VGND VPWR VPWR _3709_/X
+ sky130_fd_sc_hd__o41a_2
XFILLER_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4127__A1 _3636_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5324__A0 _6185_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4678__A2 _4699_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5875__A1 _5871_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3724__B _3724_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3886__B1 _3885_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5627__A1 _6040_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4836__A _4856_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3638__B1 _3816_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4555__B _4555_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5667__A _5667_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5386__B _5386_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3810__B1 _3763_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3187__A _4004_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4366__B2 _4602_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4118__A1 _3403_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5315__A0 _6181_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6101__CLK _6145_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5866__A1 _5240_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4669__A2 _5140_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3877__B1 _3844_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4746__A _4746_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_67_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3892__A3 _3512_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3650__A _3781_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5094__A2 _5444_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4841__A2 _4839_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3991_ _3588_/B _3593_/D _3703_/A _3643_/A _3990_/X VGND VGND VPWR VPWR _3992_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_74_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4054__B1 _3748_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5251__C1 _5250_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4481__A _4642_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5730_ _4398_/X _4671_/X _5944_/C _4657_/A VGND VGND VPWR VPWR _5733_/B sky130_fd_sc_hd__a31o_1
XANTENNA__3801__B1 _3571_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5661_ _5661_/A _5661_/B VGND VGND VPWR VPWR _5661_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4612_ _4273_/Y _4211_/A _4536_/X _4619_/B VGND VGND VPWR VPWR _4612_/X sky130_fd_sc_hd__o211a_1
X_5592_ _6156_/Q _6024_/Q _5594_/S VGND VGND VPWR VPWR _5593_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4543_ _4543_/A VGND VGND VPWR VPWR _5000_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4109__A1 _3580_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5306__A0 _6193_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4474_ _4852_/A _4865_/A _4472_/X _4865_/D _4742_/A VGND VGND VPWR VPWR _4474_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__5857__A1 _4964_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3425_ _3525_/A _3631_/A _3780_/A VGND VGND VPWR VPWR _3425_/X sky130_fd_sc_hd__and3_1
XFILLER_112_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6144_ _6146_/CLK _6144_/D VGND VGND VPWR VPWR _6144_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3356_ _3293_/X _3300_/X _3302_/X _3355_/X VGND VGND VPWR VPWR _3356_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_100_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4656__A _4656_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _3243_/X _3268_/Y _3284_/X _3286_/X VGND VGND VPWR VPWR _3287_/X sky130_fd_sc_hd__a31o_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6075_ _6176_/CLK _6075_/D VGND VGND VPWR VPWR _6075_/Q sky130_fd_sc_hd__dfxtp_1
X_5026_ _4437_/A _5009_/X _5008_/X _4472_/X VGND VGND VPWR VPWR _5026_/X sky130_fd_sc_hd__a31o_4
XFILLER_85_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4817__C1 _4816_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5085__A2 _5059_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4045__B1 _4043_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5793__B1 _4673_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4596__A1 _4573_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3399__A2 _3847_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5928_ _5076_/X _4604_/X _5098_/X _4967_/X VGND VGND VPWR VPWR _5928_/Y sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__5487__A _5487_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3719__B _3719_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4060__A3 _4059_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5859_ _4777_/X _4778_/X _4581_/C _4890_/B _5944_/B VGND VGND VPWR VPWR _5859_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_70_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3438__C _4152_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6124__CLK _6147_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4899__A2 _4878_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3157__D _3586_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3735__A _3780_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5848__A1 _5843_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4566__A _4566_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3470__A _3611_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4284__B1 _6135_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4285__B _4285_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input15_A memory_dmem_request_put[41] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5397__A _5499_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4732__C _4732_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3629__B _3687_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5784__B1 _5754_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4339__B2 _4332_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4339__A1 _5687_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4121__B1_N _4120_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3547__C1 _4036_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3645__A _3645_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5839__A1 _5018_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3314__A2 _4135_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3210_ _3864_/B VGND VGND VPWR VPWR _3692_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4190_ _5646_/A VGND VGND VPWR VPWR _4190_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4476__A _5170_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_67_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3141_ _3707_/A VGND VGND VPWR VPWR _3695_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_94_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3380__A _3603_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4814__A2 _4643_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3072_ _6195_/Q _6071_/Q _3072_/S VGND VGND VPWR VPWR _3073_/A sky130_fd_sc_hd__mux2_4
XANTENNA__5472__C1 _5471_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4027__B1 _3574_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5775__B1 _5118_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3974_ _4048_/B _4065_/B _3553_/X _3631_/X _3410_/A VGND VGND VPWR VPWR _4128_/B
+ sky130_fd_sc_hd__o32a_2
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6147__CLK _6147_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5713_ _5708_/Y _5709_/Y _5237_/A _5712_/Y VGND VGND VPWR VPWR _5713_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5527__B1 _5504_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5644_ _4975_/X _5444_/A _5490_/X _5643_/X VGND VGND VPWR VPWR _5644_/X sky130_fd_sc_hd__a31o_1
XFILLER_108_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3002__A1 _6152_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3555__A _3687_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5542__A3 _5529_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5575_ _6148_/Q _6017_/Q _5583_/S VGND VGND VPWR VPWR _5576_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4526_ _5188_/C VGND VGND VPWR VPWR _5878_/B sky130_fd_sc_hd__buf_2
XANTENNA__4750__A1 _4777_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4457_ _4890_/C VGND VGND VPWR VPWR _4457_/X sky130_fd_sc_hd__clkbuf_4
X_3408_ _3674_/B _3807_/A _3401_/Y _3407_/X VGND VGND VPWR VPWR _3408_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4502__A1 _4633_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4388_ _4374_/X _4378_/Y _5102_/B _4387_/X VGND VGND VPWR VPWR _4388_/X sky130_fd_sc_hd__a31o_1
XANTENNA_input7_A memory_dmem_request_put[33] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6127_ _6147_/CLK _6127_/D VGND VGND VPWR VPWR _6127_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3856__A3 _3821_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5058__A2 _4777_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_85_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4386__A _4555_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3339_ _3864_/B VGND VGND VPWR VPWR _3546_/A sky130_fd_sc_hd__clkbuf_2
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3290__A _4103_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6058_ _6207_/CLK _6058_/D VGND VGND VPWR VPWR _6058_/Q sky130_fd_sc_hd__dfxtp_1
X_5009_ _5009_/A VGND VGND VPWR VPWR _5009_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_54_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4805__A2 _4717_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6007__A1 _5291_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4569__A1 _4746_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4018__B1 _4015_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5230__A2 _5123_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5766__B1 _5765_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5367__D _6144_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5781__A3 _5064_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5518__B1 _6131_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3529__C1 _3537_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5533__A3 _5092_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4741__A1 _4738_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5383__C _5383_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3615__D _3666_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6198__D _6198_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5151__D1 _4316_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5680__A _5680_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4296__A _5744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5049__A2 _4783_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output121_A _3016_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4009__B1 _4008_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4024__A3 _3508_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3359__B _3359_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3783__A2 _3780_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4980__A1 _4716_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3690_ _4124_/C _3645_/B _3612_/X _3685_/X _3689_/Y VGND VGND VPWR VPWR _3690_/Y
+ sky130_fd_sc_hd__o2111ai_1
XANTENNA__2991__B1 _6060_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3375__A _3589_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5524__A3 _5498_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3535__A2 _3533_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3806__C _3816_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5360_ _5360_/A VGND VGND VPWR VPWR _6093_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5293__C input2/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4311_ _4405_/A _4333_/A _4313_/A VGND VGND VPWR VPWR _4787_/A sky130_fd_sc_hd__and3_1
X_5291_ input2/X _6205_/Q _6179_/Q _6202_/Q VGND VGND VPWR VPWR _5291_/X sky130_fd_sc_hd__and4b_2
XFILLER_114_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4242_ _4224_/X _4237_/X _4239_/X _4241_/X VGND VGND VPWR VPWR _4242_/X sky130_fd_sc_hd__o2bb2a_2
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4173_ _4301_/C VGND VGND VPWR VPWR _4405_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_95_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3124_ _3124_/A VGND VGND VPWR VPWR _3124_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4934__A _4934_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3055_ _3055_/A VGND VGND VPWR VPWR _3055_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5996__B1 _5995_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3471__A1 _3571_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5748__B1 _5740_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3957_ _3612_/D _4035_/C _3700_/A VGND VGND VPWR VPWR _3992_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__5212__A2 _4552_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3269__B _3754_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5763__A3 _5762_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3774__A2 _3881_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4971__B2 _4405_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3888_ _3636_/X _3522_/X _3882_/X _3635_/X _3887_/X VGND VGND VPWR VPWR _3888_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__5484__B _5528_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4318__A4 _4246_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5627_ _6172_/Q _6040_/Q _5627_/S VGND VGND VPWR VPWR _5628_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3285__A _3301_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5920__B1 _4665_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5558_ _5988_/A _5558_/B VGND VGND VPWR VPWR _5559_/A sky130_fd_sc_hd__or2_1
XANTENNA__4723__B2 _4722_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3918__D_N _3538_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4509_ _4975_/A VGND VGND VPWR VPWR _4630_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_105_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5489_ _5201_/X _5202_/Y _5405_/X _6011_/B _5488_/X VGND VGND VPWR VPWR _6122_/D
+ sky130_fd_sc_hd__o311ai_1
XFILLER_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4487__B1 _4864_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3732__B _3904_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5684__C1 _5683_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5005__A _5005_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3986__A_N _3839_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5987__B1 _5570_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5739__B1 _5738_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4962__A1 _4783_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3765__A2 _3767_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input82_A memory_imem_request_put[8] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3195__A _3195_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5911__B1 _5782_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4714__A1 _6048_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4714__B2 _4713_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3922__C1 _3921_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5614__S _5616_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3642__B _3648_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4738__B _4738_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4754__A _4754_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5978__B1 _5228_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3989__C1 _3802_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4860_ _4860_/A _4860_/B _4860_/C VGND VGND VPWR VPWR _4936_/A sky130_fd_sc_hd__nand3_1
XFILLER_33_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3811_ _3806_/X _3810_/Y _3727_/X _6029_/Q _3728_/X VGND VGND VPWR VPWR _6029_/D
+ sky130_fd_sc_hd__a32o_1
X_4791_ _4243_/A _4482_/B _4247_/A _4738_/B _4318_/Y VGND VGND VPWR VPWR _4792_/A
+ sky130_fd_sc_hd__o311a_2
XANTENNA__5585__A _5618_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3742_ _3534_/X _3938_/B _3608_/X _3741_/Y VGND VGND VPWR VPWR _3742_/X sky130_fd_sc_hd__a31o_1
X_3673_ _3673_/A _3673_/B VGND VGND VPWR VPWR _3673_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__5902__B1 _5901_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5412_ _5432_/A VGND VGND VPWR VPWR _5412_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3913__C1 _4149_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput113 _3067_/X VGND VGND VPWR VPWR memory_dmem_response_get[3] sky130_fd_sc_hd__buf_2
Xoutput124 _3022_/X VGND VGND VPWR VPWR memory_imem_response_get[13] sky130_fd_sc_hd__buf_2
Xoutput102 _3109_/X VGND VGND VPWR VPWR memory_dmem_response_get[22] sky130_fd_sc_hd__buf_2
X_5343_ _5343_/A VGND VGND VPWR VPWR _6085_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__4929__A _4929_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput146 _3007_/X VGND VGND VPWR VPWR memory_imem_response_get[6] sky130_fd_sc_hd__buf_2
Xoutput135 _3044_/X VGND VGND VPWR VPWR memory_imem_response_get[24] sky130_fd_sc_hd__buf_2
XANTENNA__5115__D1 _4923_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4469__B1 _4468_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5274_ input5/X VGND VGND VPWR VPWR _6014_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__5130__A1 input28/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4225_ _4225_/A VGND VGND VPWR VPWR _5438_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5130__B2 input12/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5681__A2 _5118_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4484__A3 _4309_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4156_ _4151_/X _4155_/X _3508_/A VGND VGND VPWR VPWR _4156_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_55_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3107_ _5294_/A VGND VGND VPWR VPWR _3116_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_55_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4087_ _3749_/X _4082_/X _4086_/Y _3707_/X VGND VGND VPWR VPWR _4088_/B sky130_fd_sc_hd__a31o_1
XANTENNA__5969__B1 _5905_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4641__B1 _5710_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3444__B2 _3591_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3038_ _3038_/A VGND VGND VPWR VPWR _3038_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3995__A2 _3382_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5197__A1 _4420_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5495__A _5715_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4989_ _5392_/C _5438_/C _4193_/C _4195_/A VGND VGND VPWR VPWR _5042_/A sky130_fd_sc_hd__a31o_2
XFILLER_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4944__A1 _4680_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3747__A2 _3319_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4157__C1 _4156_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5121__A1 _4882_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3462__B _3462_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5672__A2 _4501_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4880__B1 _5755_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3683__A1 _3682_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4574__A _4574_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5424__A2 _5395_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3435__A1 _3315_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4293__B _4293_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4632__B1 _5044_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3918__A _3918_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3738__A2 _3737_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput15 memory_dmem_request_put[41] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__buf_2
Xinput26 memory_dmem_request_put[52] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_1
Xinput37 memory_dmem_request_put[63] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__6013__B _6013_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput48 memory_dmem_request_put[74] VGND VGND VPWR VPWR _4333_/A sky130_fd_sc_hd__clkbuf_4
Xinput59 memory_dmem_request_put[85] VGND VGND VPWR VPWR _4217_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__5896__C1 _5118_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3653__A _3653_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4163__A2 _3807_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5344__S _5350_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5112__A1 _5109_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5663__A2 _5662_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4010_ _3895_/X _3760_/X _3722_/X _3763_/X _4009_/X VGND VGND VPWR VPWR _4010_/Y
+ sky130_fd_sc_hd__o311ai_2
XANTENNA__3123__A0 _6050_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4871__B1 _4956_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3613__D_N _3562_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3426__A1 _3522_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5961_ _5076_/X _4971_/X _4395_/A _4316_/X VGND VGND VPWR VPWR _5961_/X sky130_fd_sc_hd__a31o_1
XFILLER_52_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3977__A2 _3574_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4912_ _5924_/A VGND VGND VPWR VPWR _5822_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5820__C1 _4984_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5892_ _4959_/X _5890_/X _5891_/X _4875_/X VGND VGND VPWR VPWR _5892_/X sky130_fd_sc_hd__o211a_2
X_4843_ _4843_/A _4843_/B _4843_/C VGND VGND VPWR VPWR _4843_/X sky130_fd_sc_hd__and3_1
XANTENNA__5718__A3 _4887_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3828__A _3828_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4774_ _5073_/A VGND VGND VPWR VPWR _4937_/A sky130_fd_sc_hd__buf_4
XANTENNA__4650__C _5710_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5746__C _5746_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3729__A2 _3726_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3725_ _4126_/B _3718_/X _3721_/Y _3724_/Y VGND VGND VPWR VPWR _3725_/X sky130_fd_sc_hd__o31a_1
XANTENNA__3039__S _3043_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3656_ _3649_/Y _3655_/X _4102_/A VGND VGND VPWR VPWR _3656_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__4659__A _4728_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3587_ _3956_/C _3983_/C _3278_/A VGND VGND VPWR VPWR _3594_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__4154__A2 _3881_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3898__D1 _3897_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3563__A _4036_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3362__B1 _3983_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4378__B _4673_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3901__A2 _3895_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5326_ _6186_/Q _6078_/Q _5328_/S VGND VGND VPWR VPWR _5327_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5103__A1 _5048_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5257_ input5/X VGND VGND VPWR VPWR _5545_/A sky130_fd_sc_hd__inv_2
XANTENNA__5654__A2 _5867_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4208_ _4282_/A _4244_/A _4264_/C _4245_/A VGND VGND VPWR VPWR _4209_/A sky130_fd_sc_hd__nor4_4
XANTENNA__3114__A0 _6047_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5188_ _5188_/A _5188_/B _5188_/C _5188_/D VGND VGND VPWR VPWR _5706_/B sky130_fd_sc_hd__nand4_4
XFILLER_68_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3665__B2 _3562_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3665__A1 _3646_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_83_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4394__A _4642_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4139_ _4039_/B _4135_/X _4136_/X _4138_/X VGND VGND VPWR VPWR _4139_/X sky130_fd_sc_hd__a31o_1
XFILLER_43_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5406__A2 _5395_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4090__A1 _3299_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4090__B2 _3510_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5709__A3 _4385_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5590__A1 _6023_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3473__A _3870_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4145__A2 _3762_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5342__A1 _6085_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3904__C _3904_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4288__B _4298_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5893__A2 _5757_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input45_A memory_dmem_request_put[71] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5645__A2 _5166_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3105__A0 _6058_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4853__B1 _4255_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3656__A1 _3649_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3408__A1 _3674_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4605__B1 _4960_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3408__B2 _3407_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6030__CLK _6045_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4081__A1 _4072_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4081__B2 _3891_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5339__S _5339_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3648__A _3648_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4908__A1 _4716_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4384__A2 _4883_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5030__B1 _4927_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6180__CLK _6204_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5581__A1 _6019_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3510_ _3586_/A _3719_/B _3983_/C _4092_/D VGND VGND VPWR VPWR _3510_/X sky130_fd_sc_hd__or4_4
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4490_ _4929_/A VGND VGND VPWR VPWR _4843_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_6_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3383__A _3383_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4479__A _4543_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3441_ _3873_/B VGND VGND VPWR VPWR _3719_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__4136__A2 _3829_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5333__A1 _6081_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5884__A2 _4956_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3372_ _3956_/B VGND VGND VPWR VPWR _4073_/A sky130_fd_sc_hd__clkbuf_2
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6160_ _6201_/CLK _6160_/D VGND VGND VPWR VPWR _6160_/Q sky130_fd_sc_hd__dfxtp_1
X_5111_ _4693_/X _4735_/Y _5050_/Y _4890_/B _4572_/X VGND VGND VPWR VPWR _5111_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _6204_/CLK _6091_/D VGND VGND VPWR VPWR _6091_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4844__B1 _4649_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4926__B _4926_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _5042_/A VGND VGND VPWR VPWR _5042_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4942__A _4942_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5944_ _5944_/A _5944_/B _5944_/C _5944_/D VGND VGND VPWR VPWR _5944_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__4072__A1 _4064_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5757__B _5757_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5875_ _5871_/X _5845_/X _5874_/X VGND VGND VPWR VPWR _5875_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3558__A _3968_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4826_ _4821_/Y _4822_/X _4823_/X _4825_/Y VGND VGND VPWR VPWR _4826_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_61_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4757_ _4369_/C _4619_/B _4725_/A _4882_/A VGND VGND VPWR VPWR _4757_/X sky130_fd_sc_hd__a31o_2
XANTENNA__5572__B2 _5571_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4688_ _4869_/A VGND VGND VPWR VPWR _5829_/C sky130_fd_sc_hd__clkbuf_4
X_3708_ _3708_/A VGND VGND VPWR VPWR _3911_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4127__A2 _4123_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3639_ _3628_/X _3635_/X _3637_/X _3638_/Y VGND VGND VPWR VPWR _3639_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5324__A1 _6077_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4532__C1 _4531_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3293__A _3526_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5875__A2 _5845_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3886__B2 _3549_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3886__A1 _3551_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5309_ _6194_/Q _6070_/Q _5317_/S VGND VGND VPWR VPWR _5310_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3638__A1 _3881_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6053__CLK _6196_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4555__C _4787_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4852__A _4852_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4063__A1 _3926_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5667__B _5667_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4571__B _4859_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3810__A1 _3760_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3468__A _3468_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5386__C _6014_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5012__B1 _5011_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4118__A2 _3815_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5315__A1 _6073_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5866__A2 _5903_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3877__A1 _3343_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3877__B2 _3876_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4746__B _4746_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4826__B1 _4823_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4841__A3 _4840_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5251__B1 _4395_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3990_ _3397_/A _3781_/C _3657_/C _3582_/B _3600_/A VGND VGND VPWR VPWR _3990_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_62_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4054__A1 _4053_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3801__A1 _3614_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5660_ _4369_/D _4574_/A _4440_/Y _4675_/A VGND VGND VPWR VPWR _5661_/B sky130_fd_sc_hd__o211ai_4
XANTENNA__3378__A _3436_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4611_ _4729_/B VGND VGND VPWR VPWR _4619_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_90_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5593__A _5593_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5591_ _5591_/A VGND VGND VPWR VPWR _6155_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4542_ _4532_/Y _4539_/X _4541_/X VGND VGND VPWR VPWR _4542_/X sky130_fd_sc_hd__a21o_1
X_4473_ _4926_/C VGND VGND VPWR VPWR _4865_/D sky130_fd_sc_hd__buf_2
XANTENNA__4109__A2 _3911_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5306__A1 _6069_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3424_ _3802_/A VGND VGND VPWR VPWR _3780_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5857__A2 _5140_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4002__A _4002_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4937__A _4937_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3841__A _3841_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3355_ _3324_/X _3352_/Y _3508_/A VGND VGND VPWR VPWR _3355_/X sky130_fd_sc_hd__a21o_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6143_ _6205_/CLK _6143_/D VGND VGND VPWR VPWR _6143_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6076__CLK _6176_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _6074_/CLK _6074_/D VGND VGND VPWR VPWR _6074_/Q sky130_fd_sc_hd__dfxtp_1
X_3286_ _3828_/A VGND VGND VPWR VPWR _3286_/X sky130_fd_sc_hd__buf_2
X_5025_ _4707_/D _4619_/B _5003_/C VGND VGND VPWR VPWR _5025_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__4817__B1 _4813_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3052__S _3054_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5490__B1 _5042_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4672__A _4672_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5242__B1 _4836_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4045__B2 _3975_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4045__A1 _3764_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4596__A2 _4583_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5793__A1 _4296_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5927_ _5118_/Y _5973_/B _4839_/Y _4563_/X VGND VGND VPWR VPWR _5927_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_53_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3288__A _3918_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5858_ _5734_/X _5856_/Y _5982_/C _5175_/X _5857_/Y VGND VGND VPWR VPWR _5858_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_21_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3438__D _3983_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5789_ _5175_/X _5784_/Y _5673_/A _5788_/Y VGND VGND VPWR VPWR _5789_/Y sky130_fd_sc_hd__o211ai_4
X_4809_ _4801_/X _4802_/X _4806_/Y _4808_/Y _4189_/A VGND VGND VPWR VPWR _4809_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3735__B _4092_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5008__A _5008_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5848__A2 _5844_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4808__B1 _4224_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4284__A1 _4293_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4285__C _4301_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4582__A _4875_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5233__B1 _4954_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5784__A1 _5778_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5784__B2 _5783_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3795__B1 _3539_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3198__A _3822_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4992__C1 _5042_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4339__A2 _5687_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3926__A _4048_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3547__B1 _3476_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3645__B _3645_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6099__CLK _6207_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5839__A2 _4456_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2985__B_N _6060_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_2_1_0_CLK clkbuf_2_1_0_CLK/A VGND VGND VPWR VPWR clkbuf_3_3_0_CLK/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3140_ _3353_/A VGND VGND VPWR VPWR _3707_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3380__B _3781_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3071_ _3071_/A VGND VGND VPWR VPWR _3071_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5472__B1 _5540_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4814__A3 _4864_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3483__C1 _3374_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4027__A1 _3549_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5775__A1 _5761_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5224__B1 _5223_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5712_ _5712_/A _5746_/A _5712_/C _5712_/D VGND VGND VPWR VPWR _5712_/Y sky130_fd_sc_hd__nand4_1
X_3973_ _3961_/Y _3972_/Y _3821_/X _6036_/Q _3822_/X VGND VGND VPWR VPWR _6036_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_50_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5914__A1_N _4657_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5527__A1 _4801_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5527__B2 _4277_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5643_ _5643_/A _5643_/B _6123_/Q VGND VGND VPWR VPWR _5643_/X sky130_fd_sc_hd__and3_1
X_5574_ _5618_/A VGND VGND VPWR VPWR _5583_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_116_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4525_ _4729_/B VGND VGND VPWR VPWR _5188_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__4750__A2 _4778_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4456_ _5667_/B _5029_/A _4780_/A _4623_/A VGND VGND VPWR VPWR _4456_/X sky130_fd_sc_hd__or4_4
XANTENNA__4667__A _4855_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4387_ _4642_/A VGND VGND VPWR VPWR _4387_/X sky130_fd_sc_hd__buf_2
X_3407_ _3403_/X _3767_/D _3882_/B _3374_/X VGND VGND VPWR VPWR _3407_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4502__A2 _4501_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_85_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3338_ _3835_/A _3499_/A VGND VGND VPWR VPWR _3338_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__3571__A _3571_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6126_ _6207_/CLK _6126_/D VGND VGND VPWR VPWR _6126_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5058__A3 _4778_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_85_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3615__A_N _3308_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3269_ _3904_/A _3754_/A VGND VGND VPWR VPWR _4074_/C sky130_fd_sc_hd__nor2_4
XFILLER_46_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6057_ _6203_/CLK _6057_/D VGND VGND VPWR VPWR _6057_/Q sky130_fd_sc_hd__dfxtp_1
X_5008_ _5008_/A VGND VGND VPWR VPWR _5008_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_73_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4018__A1 _3699_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5498__A _5529_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6007__A2 _5294_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5215__B1 _5214_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4018__B2 _4017_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4569__A2 _4563_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5766__A1 _5175_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3777__B1 _3562_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5518__A1 _5495_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5518__B2 _5503_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3746__A _3746_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3529__B1 _3749_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4741__A2 _4729_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5151__C1 _4574_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4577__A _5067_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5680__B _5680_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3481__A _3876_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5049__A3 _4890_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4009__A1 _4003_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output114_A _3069_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4009__B2 _3479_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5201__A input6/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5206__B1 _5204_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4965__C1 _5005_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3359__C _3359_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3768__B1 _3695_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3783__A3 _3782_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4980__A2 _4513_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2991__A1 _3060_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3940__B1 _3939_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4310_ _4482_/A _4308_/X _4309_/X _6137_/Q VGND VGND VPWR VPWR _5061_/A sky130_fd_sc_hd__o31a_1
X_5290_ _5285_/X _5286_/Y _5289_/Y VGND VGND VPWR VPWR _6064_/D sky130_fd_sc_hd__a21oi_1
XFILLER_114_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4241_ _4807_/A VGND VGND VPWR VPWR _4241_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3391__A _3647_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5693__B1 _4563_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4172_ _4205_/A _4205_/B _4205_/C _4205_/D VGND VGND VPWR VPWR _4301_/C sky130_fd_sc_hd__and4_4
X_3123_ _6050_/Q _6094_/Q _3127_/S VGND VGND VPWR VPWR _3124_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4934__B _4934_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3054_ _6044_/Q _6176_/Q _3054_/S VGND VGND VPWR VPWR _3055_/A sky130_fd_sc_hd__mux2_1
XANTENNA__6114__CLK _6123_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5996__A1 _5570_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3471__A2 _3468_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5748__B2 _5747_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5748__A1 _4570_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3956_ _3956_/A _3956_/B _3956_/C VGND VGND VPWR VPWR _4035_/C sky130_fd_sc_hd__or3_1
XANTENNA__5212__A3 _4953_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4950__A _4950_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3566__A _3802_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3887_ _3717_/X _3883_/X _3476_/B _3886_/Y VGND VGND VPWR VPWR _3887_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3774__A3 _3195_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5626_ _5626_/A VGND VGND VPWR VPWR _6171_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5920__A1 _5918_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5557_ _5256_/A _5260_/A _5431_/B _6144_/Q _5482_/X VGND VGND VPWR VPWR _5558_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_117_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3931__B1 _3308_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5488_ _6122_/Q _4239_/X _4801_/X _5092_/X VGND VGND VPWR VPWR _5488_/X sky130_fd_sc_hd__a2bb2o_1
X_4508_ _5805_/A VGND VGND VPWR VPWR _4975_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4397__A _5188_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4439_ _4926_/B VGND VGND VPWR VPWR _4551_/A sky130_fd_sc_hd__buf_4
XANTENNA__4487__A1 _4483_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5684__B1 _5682_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3732__C _3904_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_86_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6109_ _6123_/CLK _6109_/D VGND VGND VPWR VPWR _6109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5987__A1 _5984_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5987__B2 _5998_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5021__A _5021_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5739__B2 _4793_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4860__A _4860_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4962__A2 _4827_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3476__A _3476_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3765__A3 _3882_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3195__B _3195_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5911__A1 _5712_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input75_A memory_imem_request_put[11] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4714__A2 _4629_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3922__B1 _3909_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4738__C _4772_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5675__B1 _5651_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6137__CLK _6146_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5630__S _5638_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5978__A1 _5976_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5427__B1 _5398_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3989__B1 _3319_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4938__C1 _4937_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4790_ _4680_/X _4783_/X _5761_/A _4785_/X _4789_/X VGND VGND VPWR VPWR _4790_/X
+ sky130_fd_sc_hd__a311o_1
X_3810_ _3760_/X _3457_/X _3762_/X _3763_/X _3809_/X VGND VGND VPWR VPWR _3810_/Y
+ sky130_fd_sc_hd__o311ai_2
X_3741_ _3509_/Y _3740_/Y _3282_/A VGND VGND VPWR VPWR _3741_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3386__A _3386_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3672_ _3223_/X _3230_/X _3653_/X _3327_/X VGND VGND VPWR VPWR _3672_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5902__A1 _4858_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5411_ _5406_/Y _5409_/Y _5410_/X VGND VGND VPWR VPWR _6102_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__3913__B1 _4073_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput114 _3069_/X VGND VGND VPWR VPWR memory_dmem_response_get[4] sky130_fd_sc_hd__buf_2
Xoutput125 _3025_/X VGND VGND VPWR VPWR memory_imem_response_get[14] sky130_fd_sc_hd__buf_2
Xoutput103 _3111_/X VGND VGND VPWR VPWR memory_dmem_response_get[23] sky130_fd_sc_hd__buf_2
X_5342_ _6057_/Q _6085_/Q _5350_/S VGND VGND VPWR VPWR _5343_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5115__C1 _5711_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4929__B _4929_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput147 _3009_/X VGND VGND VPWR VPWR memory_imem_response_get[7] sky130_fd_sc_hd__buf_2
Xoutput136 _3047_/X VGND VGND VPWR VPWR memory_imem_response_get[25] sky130_fd_sc_hd__buf_2
XFILLER_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5666__B1 _4730_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4469__A1 _4457_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5273_ _5286_/B input3/X _5272_/Y VGND VGND VPWR VPWR _5275_/B sky130_fd_sc_hd__a21o_1
XFILLER_102_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5130__A2 _4978_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4224_ _4224_/A VGND VGND VPWR VPWR _4224_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4945__A _4945_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4155_ _3666_/X _3308_/X _4152_/X _4154_/X VGND VGND VPWR VPWR _4155_/X sky130_fd_sc_hd__a31o_1
XFILLER_68_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3106_ _3106_/A VGND VGND VPWR VPWR _3106_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4664__B _4664_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4086_ _3975_/A _4083_/X _4085_/Y VGND VGND VPWR VPWR _4086_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5969__A1 _6108_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4641__A1 _4855_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3060__S _3060_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3037_ _6036_/Q _6168_/Q _3043_/S VGND VGND VPWR VPWR _3038_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4680__A _4680_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5197__A2 _4464_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4988_ _4984_/X _5757_/C _5757_/D _6117_/Q _4987_/X VGND VGND VPWR VPWR _4988_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_109_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4944__A2 _4761_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3601__C1 _4073_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3296__A _3799_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3939_ _4105_/B _3271_/A _3904_/D _3938_/X VGND VGND VPWR VPWR _3939_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3747__A3 _3968_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4157__B1 _4088_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5609_ _5609_/A VGND VGND VPWR VPWR _6163_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5016__A _5016_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5657__B1 _5656_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5121__A2 _5118_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4855__A _4855_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4880__A1 _4671_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3683__A2 _3350_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_86_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3435__A2 _3513_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4093__C1 _4092_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4632__A1 _4716_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3918__B _3918_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput16 memory_dmem_request_put[42] VGND VGND VPWR VPWR _5431_/A sky130_fd_sc_hd__clkbuf_2
Xinput27 memory_dmem_request_put[53] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4148__B1 _4146_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput49 memory_dmem_request_put[75] VGND VGND VPWR VPWR _4341_/B sky130_fd_sc_hd__buf_2
Xinput38 memory_dmem_request_put[64] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__6013__C _6013_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5896__B1 _5903_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3934__A _3975_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4012__B1_N _3654_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5625__S _5627_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3653__B _3653_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5648__A0 _6145_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5112__A2 _5110_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4765__A _4765_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3123__A1 _6094_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4871__A1 _4565_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3426__A2 _3425_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5960_ _4750_/Y _5899_/X _4965_/Y _5782_/X VGND VGND VPWR VPWR _5960_/X sky130_fd_sc_hd__a31o_1
XFILLER_52_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5891_ _5211_/X _5745_/B _5903_/D _5213_/X VGND VGND VPWR VPWR _5891_/X sky130_fd_sc_hd__a31o_1
X_4911_ _2986_/B _5640_/D _4984_/A _5162_/A VGND VGND VPWR VPWR _5924_/A sky130_fd_sc_hd__o2bb2a_2
XANTENNA__5820__B1 _5163_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3977__A3 _3626_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5596__A _5618_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4842_ _4950_/A _4841_/Y _4732_/B VGND VGND VPWR VPWR _4842_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4773_ _4945_/A _4852_/A _4353_/A _5188_/A VGND VGND VPWR VPWR _4773_/Y sky130_fd_sc_hd__o211ai_4
XANTENNA__5746__D _5746_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3729__A3 _3727_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4650__D _4879_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3724_ _3724_/A _3724_/B VGND VGND VPWR VPWR _3724_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4139__B1 _4138_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3655_ _3652_/Y _3653_/X _3654_/X VGND VGND VPWR VPWR _3655_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5887__B1 _4923_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3844__A _3893_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3362__A1 _3632_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3586_ _3586_/A _3663_/A _3876_/A VGND VGND VPWR VPWR _4116_/B sky130_fd_sc_hd__and3_2
XANTENNA__3898__C1 _3699_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3901__A3 _3215_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5325_ _5325_/A VGND VGND VPWR VPWR _6077_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5103__A2 _5018_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4378__C _4673_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5256_ _5256_/A VGND VGND VPWR VPWR _5256_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4675__A _4675_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4207_ _4265_/C VGND VGND VPWR VPWR _4245_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3114__A1 _6090_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5187_ _5755_/A _5976_/B _4574_/X _5976_/A _4675_/X VGND VGND VPWR VPWR _5187_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_68_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3665__A2 _3656_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4138_ _3926_/X _4137_/X _3709_/X VGND VGND VPWR VPWR _4138_/X sky130_fd_sc_hd__o21a_1
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4069_ _3626_/X _3254_/X _3830_/C _3938_/B _4068_/X VGND VGND VPWR VPWR _4069_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__4075__C1 _4074_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4090__A2 _4089_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3050__A0 _6042_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4123__A2_N _3571_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3754__A _3754_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3889__C1 _3787_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3904__D _3904_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4288__C _4358_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3105__A1 _6086_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input38_A memory_dmem_request_put[64] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4585__A _4585_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4853__A1 _4317_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3656__A2 _3655_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4066__C1 _3860_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4605__A1 _4777_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5802__B1 _5799_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3408__A2 _3807_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4081__A2 _4080_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5030__A1 _4761_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3648__B _3648_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4908__A2 _4513_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5030__B2 _4726_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3041__A0 _6038_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5869__B1 _5102_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5355__S _5361_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3440_ _3440_/A _3440_/B VGND VGND VPWR VPWR _3873_/B sky130_fd_sc_hd__and2_2
XANTENNA__4136__A3 _3830_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3371_ _3437_/C VGND VGND VPWR VPWR _3956_/B sky130_fd_sc_hd__clkbuf_2
X_5110_ _4761_/X _4328_/X _4882_/X _4829_/Y _4574_/X VGND VGND VPWR VPWR _5110_/Y
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_88_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6090_ _6176_/CLK _6090_/D VGND VGND VPWR VPWR _6090_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4278__A1_N _4266_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5041_ _4984_/X _5757_/C _5757_/D _6118_/Q _4987_/X VGND VGND VPWR VPWR _5041_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__4844__A1 _4878_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4926__C _4926_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3830__C _3830_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3804__C1 _3282_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5943_ _5093_/A _4362_/X _5529_/A _4364_/X _5942_/Y VGND VGND VPWR VPWR _5943_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__4072__A2 _4071_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5757__C _5757_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5874_ _5924_/A _5874_/B VGND VGND VPWR VPWR _5874_/X sky130_fd_sc_hd__or2_1
X_4825_ _4750_/Y _4917_/A _4824_/X VGND VGND VPWR VPWR _4825_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3558__B _4149_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3032__A0 _6034_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4756_ _4273_/Y _4211_/A _4536_/X _4707_/C VGND VGND VPWR VPWR _5829_/B sky130_fd_sc_hd__o211a_4
X_4687_ _4937_/B VGND VGND VPWR VPWR _5755_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__3574__A _3574_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3707_ _3707_/A VGND VGND VPWR VPWR _3707_/X sky130_fd_sc_hd__buf_2
X_3638_ _3881_/A _3535_/X _3816_/A VGND VGND VPWR VPWR _3638_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5483__A2_N _6120_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4532__B1 _4374_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3569_ _3564_/X _3815_/C _3208_/X _3568_/X VGND VGND VPWR VPWR _3569_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3886__A2 _3553_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5308_ _5365_/S VGND VGND VPWR VPWR _5317_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_0_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6100__D _6100_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5239_ _5102_/D _5008_/X _5009_/X _4547_/Y VGND VGND VPWR VPWR _5239_/X sky130_fd_sc_hd__a31o_1
XFILLER_102_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3638__A2 _3535_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3099__A0 _6055_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4852__B _5048_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4063__A2 _4062_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3749__A _4044_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5667__C _5899_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4571__C _4859_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3468__B _3468_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3810__A2 _3457_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5012__A1 _5002_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3484__A _3871_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5866__A3 _4875_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4523__B1 _4512_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3877__A2 _3875_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4000__A2_N _3998_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_67_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output144_A _3003_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4826__B2 _4825_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5251__A1 _5755_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3659__A _4034_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4054__A2 _3926_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3801__A2 _3447_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4610_ _5188_/A VGND VGND VPWR VPWR _4610_/X sky130_fd_sc_hd__buf_4
XANTENNA__5874__A _5924_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5590_ _6155_/Q _6023_/Q _5594_/S VGND VGND VPWR VPWR _5591_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4762__B1 _4761_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4541_ _4541_/A VGND VGND VPWR VPWR _4541_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3394__A _3815_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4472_ _4566_/A VGND VGND VPWR VPWR _4472_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__4109__A3 _3533_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3423_ _3447_/C _3870_/B VGND VGND VPWR VPWR _3525_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5857__A3 _4604_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4002__B _4002_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6142_ _6145_/CLK _6142_/D VGND VGND VPWR VPWR _6142_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4937__B _4937_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3354_ _3838_/A VGND VGND VPWR VPWR _3508_/A sky130_fd_sc_hd__buf_4
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3841__B _3841_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4817__A1 _4657_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _6074_/CLK _6073_/D VGND VGND VPWR VPWR _6073_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ _3301_/A VGND VGND VPWR VPWR _3828_/A sky130_fd_sc_hd__clkbuf_1
X_5024_ _5140_/A _5020_/X _5021_/X _5023_/X VGND VGND VPWR VPWR _5024_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_57_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5490__B2 _4906_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5490__A1 input31/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4953__A _5182_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5242__A1 _5239_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5778__C1 _5777_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4045__A2 _4042_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5793__A2 _5078_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5926_ _5028_/X _5880_/X _4930_/X _5148_/A _5179_/X VGND VGND VPWR VPWR _5926_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_53_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4450__C1 _4449_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3288__B _3918_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5857_ _4964_/X _5140_/D _4604_/X _5856_/Y VGND VGND VPWR VPWR _5857_/Y sky130_fd_sc_hd__o31ai_1
X_5788_ _5716_/X _5787_/Y _4498_/X VGND VGND VPWR VPWR _5788_/Y sky130_fd_sc_hd__o21ai_1
X_4808_ _6130_/Q _4807_/X _4224_/X VGND VGND VPWR VPWR _4808_/Y sky130_fd_sc_hd__o21ai_1
X_4739_ _4739_/A VGND VGND VPWR VPWR _4739_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3735__C _3904_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5848__A3 _5845_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4505__B1 _4242_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6020__CLK _6155_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4723__A1_N _4720_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6170__CLK _6203_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4808__A1 _6130_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4284__A2 _4246_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4285__D _4405_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5233__A1 _5076_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3479__A _4036_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5784__A2 _5781_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3795__A1 _3580_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4992__B1 input9/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3547__A1 _3327_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3635__B1_N _3838_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3380__C _4034_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3070_ _6194_/Q _6070_/Q _3072_/S VGND VGND VPWR VPWR _3071_/A sky130_fd_sc_hd__mux2_4
XFILLER_0_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5472__A1 _5444_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2992__S _2998_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3483__B1 _3482_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4027__A2 _3871_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5224__A1 input32/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5711_ _5711_/A _5711_/B _5745_/A VGND VGND VPWR VPWR _5712_/D sky130_fd_sc_hd__and3_2
XANTENNA__5775__A2 _5878_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3972_ _3142_/X _3971_/Y _3762_/X _3300_/X _3302_/X VGND VGND VPWR VPWR _3972_/Y
+ sky130_fd_sc_hd__o221ai_1
XANTENNA__4983__B1 _6052_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5527__A2 _4268_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5642_ _4629_/X _4630_/X _5410_/X VGND VGND VPWR VPWR _6179_/D sky130_fd_sc_hd__o21a_1
XANTENNA__4735__B1 _5182_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5573_ _5629_/A VGND VGND VPWR VPWR _5618_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__6043__CLK _6045_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4524_ _5667_/A VGND VGND VPWR VPWR _4524_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_116_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4948__A _4948_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4455_ _4654_/A _4363_/A _5756_/A VGND VGND VPWR VPWR _4623_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__4499__C1 _4498_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4386_ _4555_/B VGND VGND VPWR VPWR _4642_/A sky130_fd_sc_hd__clkbuf_2
X_3406_ _3406_/A VGND VGND VPWR VPWR _3767_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__6193__CLK _6196_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3337_ _3621_/A VGND VGND VPWR VPWR _3499_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3571__B _3571_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6125_ _6147_/CLK _6125_/D VGND VGND VPWR VPWR _6125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3268_ _3268_/A _3359_/A VGND VGND VPWR VPWR _3268_/Y sky130_fd_sc_hd__nand2_1
X_6056_ _6196_/CLK _6056_/D VGND VGND VPWR VPWR _6056_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ _4878_/Y _5118_/D _4644_/X _5006_/X VGND VGND VPWR VPWR _5007_/X sky130_fd_sc_hd__a211o_1
XFILLER_39_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3199_ _3891_/A VGND VGND VPWR VPWR _5388_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6007__A3 _6013_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5215__A1 _5836_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3299__A _3299_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4018__A2 _4013_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4569__A3 _5755_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5766__A2 _5760_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3777__A1 _3775_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5909_ _6192_/Q _4715_/X _5894_/Y _5908_/Y VGND VGND VPWR VPWR _6192_/D sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__5518__A2 _4908_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3746__B _3746_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3529__A1 _3403_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5923__C1 _5922_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3762__A _3762_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5151__B1 _4829_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5680__C _5680_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3481__B _3588_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input20_A memory_dmem_request_put[46] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4662__C1 _4661_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3465__B1 _3463_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4009__A2 _4005_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5206__A1 _4629_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5206__B2 _5205_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3768__A1 _3674_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output107_A _3120_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4965__B1 _5000_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6066__CLK _6203_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4980__A3 input40/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2991__A2 _6013_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3940__A1 _3936_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5363__S _5365_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5142__B1 _4568_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4240_ _5648_/S VGND VGND VPWR VPWR _4807_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5693__A1 _5720_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4171_ _4171_/A _4171_/B VGND VGND VPWR VPWR _4205_/D sky130_fd_sc_hd__nor2_1
XFILLER_67_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3122_ _3122_/A VGND VGND VPWR VPWR _3122_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_82_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3053_ _3053_/A VGND VGND VPWR VPWR _3053_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5996__A2 _5994_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5748__A2 _4571_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6209__151 VGND VGND VPWR VPWR _6209__151/HI memory_imem_response_get[27] sky130_fd_sc_hd__conb_1
X_3955_ _3910_/B _3975_/B _3359_/C _3954_/X _3299_/B VGND VGND VPWR VPWR _3955_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_51_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3847__A _3847_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3566__B _3870_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3886_ _3551_/A _3553_/A _3885_/X _3549_/X _3574_/X VGND VGND VPWR VPWR _3886_/Y
+ sky130_fd_sc_hd__a221oi_2
X_5625_ _6171_/Q _6039_/Q _5627_/S VGND VGND VPWR VPWR _5626_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3058__S _3060_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5920__A2 _5919_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5556_ _5405_/X _5555_/X _5388_/A VGND VGND VPWR VPWR _6143_/D sky130_fd_sc_hd__a21oi_1
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3392__C1 _3860_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3931__A1 _3867_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5487_ _5487_/A VGND VGND VPWR VPWR _6121_/D sky130_fd_sc_hd__clkbuf_1
X_4507_ _5648_/S VGND VGND VPWR VPWR _5805_/A sky130_fd_sc_hd__buf_2
XFILLER_117_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4438_ _4769_/A VGND VGND VPWR VPWR _4754_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3582__A _3686_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4487__A2 _4485_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5684__A1 _4556_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4369_ _4369_/A _5188_/A _4369_/C _4369_/D VGND VGND VPWR VPWR _4369_/Y sky130_fd_sc_hd__nand4_4
XANTENNA__3732__D _3732_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6108_ _6145_/CLK _6108_/D VGND VGND VPWR VPWR _6108_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6039_ _6074_/CLK _6039_/D VGND VGND VPWR VPWR _6039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5987__A2 _5985_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6089__CLK _6176_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_0_0_CLK clkbuf_2_1_0_CLK/A VGND VGND VPWR VPWR clkbuf_3_1_0_CLK/A sky130_fd_sc_hd__clkbuf_2
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4860__B _4860_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4947__B1 _4538_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4962__A3 _4552_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3476__B _3476_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5911__A2 _5102_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4714__A3 _4630_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input68_A memory_dmem_request_put[94] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3922__A1 _6034_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3492__A _3959_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5675__B2 _5674_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5427__A1 input15/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5427__B2 _6107_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4635__C1 _4472_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3989__A1 _3932_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5978__A2 _4556_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5928__A1_N _5076_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4938__B1 _5712_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3667__A _3870_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3740_ _3761_/A _4149_/A _3704_/X VGND VGND VPWR VPWR _3740_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_20_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3610__B1 _3608_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3671_ _3666_/X _3668_/X _3910_/A _3670_/Y VGND VGND VPWR VPWR _3671_/X sky130_fd_sc_hd__a31o_1
XFILLER_9_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5902__A2 _4859_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5363__A0 _6051_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5410_ _5422_/B VGND VGND VPWR VPWR _5410_/X sky130_fd_sc_hd__buf_6
XFILLER_114_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3913__A1 _3593_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3913__B2 _3525_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4498__A _5125_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput115 _3071_/X VGND VGND VPWR VPWR memory_dmem_response_get[5] sky130_fd_sc_hd__buf_2
Xoutput104 _3113_/X VGND VGND VPWR VPWR memory_dmem_response_get[24] sky130_fd_sc_hd__buf_2
X_5341_ _5352_/A VGND VGND VPWR VPWR _5350_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_114_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4929__C _4929_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5115__B1 _5078_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput148 _3011_/X VGND VGND VPWR VPWR memory_imem_response_get[8] sky130_fd_sc_hd__buf_2
Xoutput126 _3027_/X VGND VGND VPWR VPWR memory_imem_response_get[15] sky130_fd_sc_hd__buf_2
Xoutput137 _3049_/X VGND VGND VPWR VPWR memory_imem_response_get[26] sky130_fd_sc_hd__buf_2
XANTENNA__5666__B2 _5731_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5666__A1 _5782_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4469__A2 _4306_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5272_ _5570_/C input3/X _6062_/Q VGND VGND VPWR VPWR _5272_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3677__B1 _3539_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4223_ _4199_/X _5044_/A _5648_/S _4222_/X VGND VGND VPWR VPWR _4224_/A sky130_fd_sc_hd__a31o_2
X_4154_ _3674_/B _3881_/B _3802_/X _4153_/Y _4044_/B VGND VGND VPWR VPWR _4154_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_83_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4085_ _4084_/X _3208_/X _3649_/Y VGND VGND VPWR VPWR _4085_/Y sky130_fd_sc_hd__a21oi_1
X_3105_ _6058_/Q _6086_/Q _3105_/S VGND VGND VPWR VPWR _3106_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4664__C _4664_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3036_ _3036_/A VGND VGND VPWR VPWR _3036_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5969__A2 _4807_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4641__A2 _5745_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_83_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5197__A3 _4793_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3577__A _3838_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4987_ _6146_/Q VGND VGND VPWR VPWR _4987_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4944__A3 _4878_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3601__B1 _3746_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3938_ _4042_/C _3938_/B _3938_/C VGND VGND VPWR VPWR _3938_/X sky130_fd_sc_hd__and3_1
XFILLER_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3869_ _3867_/X _3910_/C _3773_/C _3603_/X _3868_/X VGND VGND VPWR VPWR _3869_/Y
+ sky130_fd_sc_hd__a311oi_1
XANTENNA__5159__A2_N _6056_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4157__A1 _4148_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5608_ _6163_/Q _6031_/Q _5616_/S VGND VGND VPWR VPWR _5609_/A sky130_fd_sc_hd__mux2_1
XANTENNA__6103__D _6103_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5539_ _5093_/X _4341_/B _4802_/X _6138_/Q _5482_/X VGND VGND VPWR VPWR _5540_/B
+ sky130_fd_sc_hd__o32a_1
XFILLER_11_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5106__B1 _4873_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4201__A _4201_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5657__A1 _4732_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3716__A1_N _3832_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4855__B _4996_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_86_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4880__A2 _5944_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4617__C1 _4946_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4093__B1 _3992_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4983__A2_N _4982_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4632__A2 _4513_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3840__B1 _3839_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3487__A _4073_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3918__C _3918_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput28 memory_dmem_request_put[54] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_1
Xinput17 memory_dmem_request_put[43] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4148__B2 _4147_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4148__A1 _3695_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6104__CLK _6146_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput39 memory_dmem_request_put[65] VGND VGND VPWR VPWR input39/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5896__A1 _4754_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3934__B _3934_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3356__C1 _3355_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3653__C _3653_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5648__A1 _5560_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4871__A2 _5711_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5555__B1_N _6143_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4084__B1 _3983_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5890_ _4824_/X _4878_/Y _5107_/A _4459_/A VGND VGND VPWR VPWR _5890_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_93_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4910_ _4910_/A VGND VGND VPWR VPWR _5162_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5820__A1 input9/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4841_ _4838_/X _4839_/Y _4840_/X _5746_/D _4739_/X VGND VGND VPWR VPWR _4841_/Y
+ sky130_fd_sc_hd__a32oi_2
XANTENNA__3397__A _3397_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4772_ _4772_/A VGND VGND VPWR VPWR _4945_/A sky130_fd_sc_hd__buf_4
X_3723_ _3701_/A _3512_/X _3722_/X _3673_/Y _3524_/X VGND VGND VPWR VPWR _3724_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4139__A1 _4039_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3654_ _4083_/B VGND VGND VPWR VPWR _3654_/X sky130_fd_sc_hd__buf_2
XFILLER_106_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5887__A1 _4890_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5887__B2 _4534_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3898__B1 _3896_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3585_ _3749_/B VGND VGND VPWR VPWR _3862_/A sky130_fd_sc_hd__buf_2
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3362__A2 _3858_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5324_ _6185_/Q _6077_/Q _5328_/S VGND VGND VPWR VPWR _5325_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4956__A _4956_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_102_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5103__A3 _5944_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5255_ _6059_/Q _5040_/X _5227_/X _5254_/Y VGND VGND VPWR VPWR _6059_/D sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__4847__C1 _4420_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4206_ _4283_/A VGND VGND VPWR VPWR _4264_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__3860__A _3860_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5186_ _5177_/Y _5180_/Y _4950_/X _5185_/X VGND VGND VPWR VPWR _5186_/Y sky130_fd_sc_hd__a211oi_4
XFILLER_95_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4137_ _3835_/X _3305_/A _4152_/B _4061_/X VGND VGND VPWR VPWR _4137_/X sky130_fd_sc_hd__o22a_1
XFILLER_113_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4068_ _3893_/C _3653_/B _3668_/A _3902_/A VGND VGND VPWR VPWR _4068_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4075__B1 _3938_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3019_ _6028_/Q _6160_/Q _3021_/S VGND VGND VPWR VPWR _3020_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5575__A0 _6148_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3100__A _3100_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6127__CLK _6147_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3050__A1 _6174_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3754__B _3754_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3889__B1 _3624_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4288__D _4354_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4853__A2 _4234_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4066__B1 _3438_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4605__A2 _4778_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5802__B2 _5801_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5802__A1 _5756_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3813__B1 _3242_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4081__A3 _3821_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4908__A3 input39/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5030__A2 _5028_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3041__A1 _6170_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5636__S _5638_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5869__A1 _4487_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output99_A _3061_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3370_ _3904_/A VGND VGND VPWR VPWR _3572_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3537__C_N _3491_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3680__A _3680_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5646_/A VGND VGND VPWR VPWR _5040_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4844__A2 _4878_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3830__D _3830_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4057__B1 _6040_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5942_ _5167_/X _5880_/X _4773_/Y VGND VGND VPWR VPWR _5942_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5254__C1 _5253_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3804__B1 _3803_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5400__A input5/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5757__D _5757_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5873_ _6103_/Q _5805_/A _5905_/A _5872_/X VGND VGND VPWR VPWR _5874_/B sky130_fd_sc_hd__o211a_1
XFILLER_21_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4824_ _4483_/X _4485_/X _4649_/A _5188_/D VGND VGND VPWR VPWR _4824_/X sky130_fd_sc_hd__o22a_4
XANTENNA__3558__C _3660_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5557__B1 _6144_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4755_ _5761_/D _4437_/Y _4754_/X _5034_/B VGND VGND VPWR VPWR _4755_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3032__A1 _6166_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3706_ _3701_/X _3705_/X _3661_/Y VGND VGND VPWR VPWR _3706_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5309__A0 _6194_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4686_ _4942_/A VGND VGND VPWR VPWR _4686_/X sky130_fd_sc_hd__buf_4
X_3637_ _3524_/X _3342_/X _4124_/D _3636_/X _3749_/D VGND VGND VPWR VPWR _3637_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__3066__S _3072_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4532__A1 _4431_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3568_ _3968_/A _3932_/B _3567_/X _3710_/C _4092_/C VGND VGND VPWR VPWR _3568_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_115_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4686__A _4942_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5307_ _5307_/A VGND VGND VPWR VPWR _6069_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3499_ _3499_/A VGND VGND VPWR VPWR _3499_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_69_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5238_ _5232_/Y _5236_/Y _5237_/X VGND VGND VPWR VPWR _5238_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__3099__A1 _6083_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5169_ _4740_/X _5102_/B _4457_/X _4652_/X VGND VGND VPWR VPWR _5169_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_29_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4852__C _4852_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5796__B1 _5704_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5310__A _5310_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4571__D _4800_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3749__B _3749_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3468__C _3621_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3810__A3 _3762_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5012__A2 _5004_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5866__A4 _4792_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4523__B2 _4522_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4523__A1 _4629_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input50_A memory_dmem_request_put[76] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output137_A _3049_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3005__A _3005_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5251__A2 _4369_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5787__B1 _5228_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5220__A _5220_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3659__B _3904_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5539__B1 _6138_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5874__B _5874_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4762__A1 _5152_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4540_ _4835_/A VGND VGND VPWR VPWR _4541_/A sky130_fd_sc_hd__buf_2
X_4471_ _4926_/B VGND VGND VPWR VPWR _4865_/A sky130_fd_sc_hd__buf_2
XANTENNA__4109__A4 _3962_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3422_ _3491_/A VGND VGND VPWR VPWR _4102_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__6201__D _6201_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6141_ _6145_/CLK _6141_/D VGND VGND VPWR VPWR _6141_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4937__C _4999_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3353_ _3353_/A VGND VGND VPWR VPWR _3838_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4278__B1 _4277_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3284_ _3359_/B _3815_/C _3674_/B _3359_/C _3283_/Y VGND VGND VPWR VPWR _3284_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _6074_/CLK _6072_/D VGND VGND VPWR VPWR _6072_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4817__A2 _4812_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5023_ _4931_/A _4740_/X _5782_/A _4948_/A VGND VGND VPWR VPWR _5023_/X sky130_fd_sc_hd__a31o_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5490__A2 _4978_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5242__A2 _5240_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5778__B1 _5006_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4450__B1 _4420_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5925_ _5915_/Y _5921_/Y _5845_/X _5924_/X VGND VGND VPWR VPWR _5925_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_34_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5856_ _5850_/X _5851_/X _4732_/B _5855_/X VGND VGND VPWR VPWR _5856_/Y sky130_fd_sc_hd__o22ai_4
XANTENNA__3288__C _3918_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4807_ _4807_/A VGND VGND VPWR VPWR _4807_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3585__A _3749_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5787_ _5722_/Y _5785_/X _5786_/X _5228_/X VGND VGND VPWR VPWR _5787_/Y sky130_fd_sc_hd__a31oi_1
X_2999_ _2999_/A VGND VGND VPWR VPWR _2999_/X sky130_fd_sc_hd__clkbuf_1
X_4738_ _4738_/A _4738_/B _4772_/A VGND VGND VPWR VPWR _4739_/A sky130_fd_sc_hd__and3_1
XANTENNA__5950__B1 _5941_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4669_ _5140_/A _5140_/B _4668_/X _4431_/X VGND VGND VPWR VPWR _4669_/Y sky130_fd_sc_hd__o22ai_2
XANTENNA__4505__B2 _4504_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5702__B1 _5701_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6111__D _6111_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5305__A _5305_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4269__B1 _4234_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4808__A2 _4807_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4284__A3 _4308_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5218__C1 _5217_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5040__A _5646_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5233__A2 _4971_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3795__A2 _3794_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4992__A1 _5438_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3495__A _3621_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3547__A2 _3543_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5941__B1 _5940_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3952__C1 _3701_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6021__D _6021_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3704__C1 _3468_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3380__D _3904_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5457__C1 _5456_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5472__A2 _5433_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3483__A1 _3621_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4027__A3 _3482_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3971_ _3962_/X _3963_/X _3964_/X _3970_/X VGND VGND VPWR VPWR _3971_/Y sky130_fd_sc_hd__a211oi_2
XANTENNA__5224__A2 _4978_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5710_ _5710_/A VGND VGND VPWR VPWR _5712_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_90_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4983__B2 _4190_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2994__A0 _6016_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5527__A3 _5092_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5641_ _5445_/X _5640_/X _5410_/X VGND VGND VPWR VPWR _6178_/D sky130_fd_sc_hd__o21a_1
XANTENNA__4735__A1 _5211_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5932__B1 _4190_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5572_ _6199_/Q _5985_/A _5570_/X _5571_/X VGND VGND VPWR VPWR _5629_/A sky130_fd_sc_hd__o2bb2a_1
X_4523_ _4629_/A _4630_/A _4512_/Y _4522_/X VGND VGND VPWR VPWR _4523_/X sky130_fd_sc_hd__o22a_1
XFILLER_116_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4454_ _4640_/A VGND VGND VPWR VPWR _5667_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__5696__C1 _5148_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4499__B1 _4495_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3405_ _3781_/D VGND VGND VPWR VPWR _3406_/A sky130_fd_sc_hd__clkbuf_4
X_4385_ _4385_/A VGND VGND VPWR VPWR _5102_/B sky130_fd_sc_hd__buf_2
XFILLER_105_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3336_ _3582_/C _3437_/C VGND VGND VPWR VPWR _3835_/A sky130_fd_sc_hd__or2_2
XANTENNA__3571__C _3571_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5125__A _5125_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6124_ _6147_/CLK _6124_/D VGND VGND VPWR VPWR _6124_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4964__A _4964_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6074_/CLK _6055_/D VGND VGND VPWR VPWR _6055_/Q sky130_fd_sc_hd__dfxtp_1
X_5006_ _5006_/A VGND VGND VPWR VPWR _5006_/X sky130_fd_sc_hd__clkbuf_2
X_3267_ _3246_/X _3249_/X _3612_/D _3998_/C _3266_/X VGND VGND VPWR VPWR _3268_/A
+ sky130_fd_sc_hd__a41o_1
XANTENNA__4120__C1 _3806_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3757__B1_N _3282_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3198_ _3822_/A VGND VGND VPWR VPWR _3891_/A sky130_fd_sc_hd__buf_2
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5215__A2 _5213_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3299__B _3299_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4569__A4 _4956_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6106__D _6106_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5908_ _5902_/Y _5955_/A _5907_/X _5769_/X VGND VGND VPWR VPWR _5908_/Y sky130_fd_sc_hd__a211oi_2
XANTENNA__3777__A2 _3776_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5839_ _5018_/D _4456_/X _5838_/Y _5175_/A VGND VGND VPWR VPWR _5839_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__5518__A3 _5498_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3529__A2 _3524_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4204__A _4265_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5923__B1 _5905_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5151__A1 _5755_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4662__B1 _5680_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3465__B2 _3464_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input13_A memory_dmem_request_put[39] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5206__A2 _4630_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6016__D _6016_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4965__A1 _4865_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3768__A2 _3748_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5914__B1 _5004_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3940__A2 _3699_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5142__A1 _5136_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5693__A2 _5720_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4170_ _4170_/A _4170_/B VGND VGND VPWR VPWR _4205_/C sky130_fd_sc_hd__nor2_1
XFILLER_95_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3121_ _6049_/Q _6093_/Q _3127_/S VGND VGND VPWR VPWR _3122_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4653__B1 _4652_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3052_ _6043_/Q _6175_/Q _3054_/S VGND VGND VPWR VPWR _3053_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3954_ _3932_/B _3847_/B _4004_/A VGND VGND VPWR VPWR _3954_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3847__B _3847_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3885_ _3773_/A _3756_/C _3841_/B _4042_/C VGND VGND VPWR VPWR _3885_/X sky130_fd_sc_hd__a31o_1
X_5624_ _5624_/A VGND VGND VPWR VPWR _6170_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3916__C1 _3546_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6160__CLK _6201_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4959__A _5020_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5555_ _2986_/B _5640_/D _6143_/Q VGND VGND VPWR VPWR _5555_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__3392__B1 _3749_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3931__A2 _3881_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5486_ _5486_/A _5501_/B VGND VGND VPWR VPWR _5487_/A sky130_fd_sc_hd__and2_1
X_4506_ _5643_/B VGND VGND VPWR VPWR _4629_/A sky130_fd_sc_hd__clkbuf_2
X_4437_ _4437_/A _5048_/A VGND VGND VPWR VPWR _4437_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3582__B _3582_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5669__C1 _5668_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5684__A2 _5680_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4368_ _4832_/A VGND VGND VPWR VPWR _4369_/C sky130_fd_sc_hd__buf_4
XFILLER_98_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4892__B1 _4541_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input5_A RST_N VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6107_ _6147_/CLK _6107_/D VGND VGND VPWR VPWR _6107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3319_ _3509_/A VGND VGND VPWR VPWR _3319_/X sky130_fd_sc_hd__clkbuf_4
X_4299_ _4268_/A _4244_/A _4308_/A _4245_/A _6134_/Q VGND VGND VPWR VPWR _4354_/A
+ sky130_fd_sc_hd__o41ai_4
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6038_ _6202_/CLK _6038_/D VGND VGND VPWR VPWR _6038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5987__A3 _5986_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4860__C _4860_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4947__A1 _4552_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4633__S _4633_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3476__C _3476_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3907__C1 _4036_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3773__A _3773_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4869__A _4869_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5911__A3 _4610_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3922__A2 _3891_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5427__A2 _5412_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4635__B1 _4955_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3989__A2 _3720_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6033__CLK _6202_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4938__A1 _4398_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5060__B1 _4675_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6183__CLK _6204_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3667__B _3667_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3610__A1 _4105_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3610__B2 _3938_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3670_ _3659_/D _3673_/B _3488_/X VGND VGND VPWR VPWR _3670_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5363__A1 _6095_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2998__S _2998_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3913__A2 _3653_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3374__B1 _3797_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput116 _3073_/X VGND VGND VPWR VPWR memory_dmem_response_get[6] sky130_fd_sc_hd__buf_2
Xoutput105 _3115_/X VGND VGND VPWR VPWR memory_dmem_response_get[25] sky130_fd_sc_hd__buf_2
X_5340_ _5340_/A VGND VGND VPWR VPWR _6084_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5115__A1 _4843_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput149 _3014_/X VGND VGND VPWR VPWR memory_imem_response_get[9] sky130_fd_sc_hd__buf_2
Xoutput127 _3029_/X VGND VGND VPWR VPWR memory_imem_response_get[16] sky130_fd_sc_hd__buf_2
Xoutput138 _3051_/X VGND VGND VPWR VPWR memory_imem_response_get[28] sky130_fd_sc_hd__buf_2
X_5271_ _5269_/Y _5270_/X _6062_/Q VGND VGND VPWR VPWR _5275_/A sky130_fd_sc_hd__a21o_1
XFILLER_114_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5666__A2 _4773_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4222_ _5757_/A _4985_/A _4986_/A _6147_/Q VGND VGND VPWR VPWR _4222_/X sky130_fd_sc_hd__o31a_1
XANTENNA__4874__B1 _4686_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3677__A1 _3508_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4153_ _3761_/A _3572_/A _3515_/B _3643_/A VGND VGND VPWR VPWR _4153_/Y sky130_fd_sc_hd__a31oi_1
X_4084_ _4004_/C _3581_/A _3703_/A _3983_/X VGND VGND VPWR VPWR _4084_/X sky130_fd_sc_hd__a31o_1
XFILLER_56_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5403__A _5757_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3104_ _3104_/A VGND VGND VPWR VPWR _3104_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4626__B1 _4596_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3035_ _6035_/Q _6167_/Q _3043_/S VGND VGND VPWR VPWR _3036_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4641__A3 _4843_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3858__A _3858_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4986_ _4986_/A VGND VGND VPWR VPWR _5757_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_24_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5051__B1 _5050_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3937_ _3910_/B _3626_/X _3573_/X _3923_/Y VGND VGND VPWR VPWR _3937_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5197__A4 _5176_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3601__A1 _3406_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3868_ _3868_/A VGND VGND VPWR VPWR _3868_/X sky130_fd_sc_hd__buf_2
XANTENNA__4689__A _5191_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3799_ _3799_/A _3847_/B _4149_/B VGND VGND VPWR VPWR _3799_/X sky130_fd_sc_hd__and3_2
XANTENNA__4157__A2 _3477_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5607_ _5618_/A VGND VGND VPWR VPWR _5616_/S sky130_fd_sc_hd__clkbuf_2
X_5538_ _5538_/A VGND VGND VPWR VPWR _6137_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5106__A1 _5008_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5106__B2 _4692_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5657__A2 _4822_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5469_ _5469_/A VGND VGND VPWR VPWR _6115_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__6056__CLK _6196_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4855__C _5761_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4880__A3 _4878_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4617__B1 _5034_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4093__A1 _3567_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5290__B1 _5289_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4632__A3 input35/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3840__A1 _3828_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput18 memory_dmem_request_put[44] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input80_A memory_imem_request_put[6] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4599__A _5067_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4148__A2 _4143_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput29 memory_dmem_request_put[55] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5896__A2 _5903_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3934__C _3934_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3356__B1 _3302_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3108__A0 _6180_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4084__A1 _4004_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5820__A2 _5395_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4840_ _4882_/A VGND VGND VPWR VPWR _4840_/X sky130_fd_sc_hd__buf_4
XFILLER_33_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5033__B1 _5721_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4771_ _5721_/B VGND VGND VPWR VPWR _4771_/X sky130_fd_sc_hd__buf_2
XANTENNA__6204__D _6204_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3722_ _3633_/A _4073_/A _3457_/A VGND VGND VPWR VPWR _3722_/X sky130_fd_sc_hd__a21o_2
XANTENNA__3595__B1 _3748_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3653_ _3653_/A _3653_/B _3653_/C VGND VGND VPWR VPWR _3653_/X sky130_fd_sc_hd__and3_2
XANTENNA__4139__A2 _4135_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5887__A2 _5761_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4302__A _4354_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3898__A1 _3998_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3584_ _4124_/D _3525_/X _3548_/X _3583_/X VGND VGND VPWR VPWR _3584_/Y sky130_fd_sc_hd__a211oi_1
X_5323_ _5323_/A VGND VGND VPWR VPWR _6076_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__6079__CLK _6203_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4847__B1 _5102_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4956__B _5971_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5254_ _5229_/X _5238_/Y _5015_/A _5253_/Y VGND VGND VPWR VPWR _5254_/Y sky130_fd_sc_hd__o211ai_4
X_5185_ _5712_/C _5181_/X _5183_/X _5184_/Y _4652_/X VGND VGND VPWR VPWR _5185_/X
+ sky130_fd_sc_hd__o311a_2
X_4205_ _4205_/A _4205_/B _4205_/C _4205_/D VGND VGND VPWR VPWR _4283_/A sky130_fd_sc_hd__nand4_4
XANTENNA__5133__A _5133_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4136_ _3536_/A _3829_/X _3830_/C _3161_/A _4061_/X VGND VGND VPWR VPWR _4136_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_3_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4067_ _4067_/A _4067_/B VGND VGND VPWR VPWR _4067_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4075__A1 _3834_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5272__B1 _6062_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_83_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3018_ _3018_/A VGND VGND VPWR VPWR _3018_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3588__A _3594_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5024__B1 _5023_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4969_ _4957_/X _4966_/Y _4968_/Y _4836_/X VGND VGND VPWR VPWR _4969_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_51_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6114__D _6114_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5575__A1 _6017_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4212__A _4282_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5308__A _5365_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3889__A1 _3881_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4838__B1 _4937_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4882__A _4882_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4066__A1 _3499_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4605__A3 _4864_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3813__A1 _3622_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5802__A2 _5757_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3498__A _3904_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6024__D _6024_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5869__A2 _4891_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4829__B1 _4864_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3501__B1 _3475_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4792__A _4792_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4057__A1 _4047_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5254__B1 _5015_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5941_ _5934_/Y _5939_/Y _5940_/X VGND VGND VPWR VPWR _5941_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4057__B2 _3822_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3804__A1 _4044_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5872_ input11/X _5420_/A _5162_/A _4984_/A VGND VGND VPWR VPWR _5872_/X sky130_fd_sc_hd__a211o_1
X_4823_ _5034_/B VGND VGND VPWR VPWR _4823_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5557__B2 _5482_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5557__A1 _5256_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4754_ _4754_/A VGND VGND VPWR VPWR _4754_/X sky130_fd_sc_hd__buf_4
XANTENNA__3568__B1 _3710_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3705_ _3343_/X _3893_/C _3534_/X _3910_/C _3704_/X VGND VGND VPWR VPWR _3705_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__5309__A1 _6070_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4685_ _4685_/A VGND VGND VPWR VPWR _4685_/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__5726__A2_N _5646_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4517__C1 _4516_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3636_ _4128_/A VGND VGND VPWR VPWR _3636_/X sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_4_8_0_CLK_A clkbuf_4_9_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4532__A2 _4524_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4967__A _4967_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3567_ _3998_/A VGND VGND VPWR VPWR _3567_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_115_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3740__B1 _3704_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3871__A _3871_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5306_ _6193_/Q _6069_/Q _5306_/S VGND VGND VPWR VPWR _5307_/A sky130_fd_sc_hd__mux2_1
X_3498_ _3904_/B VGND VGND VPWR VPWR _4083_/C sky130_fd_sc_hd__buf_4
X_5237_ _5237_/A VGND VGND VPWR VPWR _5237_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5168_ _5167_/X _4290_/Y _4927_/X _4838_/X _5020_/X VGND VGND VPWR VPWR _5168_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_75_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5099_ _5102_/D _5097_/X _5102_/C _5098_/X VGND VGND VPWR VPWR _5099_/X sky130_fd_sc_hd__a31o_1
X_4119_ _3314_/Y _3654_/X _3680_/X _4118_/Y VGND VGND VPWR VPWR _4119_/X sky130_fd_sc_hd__a211o_1
XANTENNA__6109__D _6109_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5245__B1 _5244_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4852__D _4878_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5796__B2 _5795_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4207__A _4265_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3749__C _3749_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3111__A _3111_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5221__A1_N _6058_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5012__A3 _5007_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4756__C1 _4707_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3559__B1 _3308_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5236__A1_N _4957_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5181__C1 _4686_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4877__A _5152_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4523__A2 _4630_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3781__A _3781_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input43_A memory_dmem_request_put[69] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6019__D _6019_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5236__B1 _5234_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5501__A _5501_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5787__A1 _5722_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5220__B _5220_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5251__A3 _5010_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3659__C _3966_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5539__B2 _5482_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5539__A1 _5093_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3956__A _3956_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4762__A2 _4956_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4470_ _4614_/A VGND VGND VPWR VPWR _4852_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3970__B1 _3969_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4787__A _4787_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3421_ _3327_/X _3934_/D _3414_/X _3420_/Y VGND VGND VPWR VPWR _3421_/X sky130_fd_sc_hd__o31a_1
XFILLER_112_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3722__B1 _3457_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3352_ _3327_/X _3335_/X _3338_/Y _3340_/X _3351_/Y VGND VGND VPWR VPWR _3352_/Y
+ sky130_fd_sc_hd__o311ai_1
X_6140_ _6146_/CLK _6140_/D VGND VGND VPWR VPWR _6140_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4937__D _4937_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4278__B2 _4209_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6071_ _6074_/CLK _6071_/D VGND VGND VPWR VPWR _6071_/Q sky130_fd_sc_hd__dfxtp_1
X_3283_ _3934_/C _3815_/A VGND VGND VPWR VPWR _3283_/Y sky130_fd_sc_hd__nand2_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _5022_/A VGND VGND VPWR VPWR _5782_/A sky130_fd_sc_hd__buf_2
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6117__CLK _6145_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5227__B1 _5225_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5778__A1 _5776_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5242__A3 _5241_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4450__A1 _4732_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5924_ _5924_/A _5924_/B VGND VGND VPWR VPWR _5924_/X sky130_fd_sc_hd__or2_1
XANTENNA__3789__B1 _3788_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5855_ _5852_/Y _5721_/B _5853_/X _5854_/X VGND VGND VPWR VPWR _5855_/X sky130_fd_sc_hd__a22o_1
XFILLER_21_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4806_ _4716_/X _4513_/X input38/X _4803_/X _4805_/X VGND VGND VPWR VPWR _4806_/Y
+ sky130_fd_sc_hd__o311ai_4
XANTENNA__3866__A _3918_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5786_ _5944_/B _4960_/X _4693_/X _4541_/A _5029_/X VGND VGND VPWR VPWR _5786_/X
+ sky130_fd_sc_hd__a311o_1
X_2998_ _6019_/Q _6151_/Q _2998_/S VGND VGND VPWR VPWR _2999_/A sky130_fd_sc_hd__mux2_1
X_4737_ _4735_/Y _4610_/X _4736_/Y _5152_/A VGND VGND VPWR VPWR _4737_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__5950__B2 _5949_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5950__A1 _6194_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3077__S _3083_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4668_ _4668_/A _4668_/B _4852_/C VGND VGND VPWR VPWR _4668_/X sky130_fd_sc_hd__and3_4
XANTENNA__3961__B1 _3960_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4697__A _4697_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3619_ _3749_/C _3616_/X _3868_/A _3281_/A VGND VGND VPWR VPWR _3623_/C sky130_fd_sc_hd__o211a_1
XANTENNA__5702__A1 _6111_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4599_ _5067_/A VGND VGND VPWR VPWR _5022_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3713__B1 _3712_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4269__B2 _6134_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4269__A1 _4313_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3106__A _3106_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5466__B1 _5439_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4284__A4 _4246_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5218__B1 _4584_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5321__A _5321_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5233__A3 _4459_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5790__A1_N _6186_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4992__A2 _4227_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5941__A1 _5934_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3952__B1 _3762_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5154__C1 _5153_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4103__C _4103_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3704__B1 _3876_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4400__A _4442_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3016__A _3016_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5457__B1 _5447_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5472__A3 _5470_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5209__B1 _4859_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3483__A2 _3230_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3970_ _3764_/X _3965_/Y _4105_/C _3969_/Y _3975_/C VGND VGND VPWR VPWR _3970_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4968__C1 _4730_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5128__A1_N _6055_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3686__A _3686_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2994__A1 _6149_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5640_ _6099_/Q _6098_/Q _6097_/Q _5640_/D VGND VGND VPWR VPWR _5640_/X sky130_fd_sc_hd__and4b_1
XANTENNA__4735__A2 _4873_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5932__B2 _6193_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5571_ _6199_/Q _5985_/A _6100_/Q _6197_/Q VGND VGND VPWR VPWR _5571_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3943__B1 _3941_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4522_ _4522_/A _5968_/B _5715_/A VGND VGND VPWR VPWR _4522_/X sky130_fd_sc_hd__and3_1
X_4453_ _4878_/B _4551_/A _4878_/A _4854_/A VGND VGND VPWR VPWR _5079_/A sky130_fd_sc_hd__o211ai_4
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3404_ _3437_/C VGND VGND VPWR VPWR _3781_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__5696__B1 _5148_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4499__A1 _5079_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3695__D_N _3694_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4384_ _4878_/B _4883_/A _4815_/D VGND VGND VPWR VPWR _4385_/A sky130_fd_sc_hd__o21ai_4
XFILLER_98_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3335_ _4083_/A _4074_/A _4074_/B VGND VGND VPWR VPWR _3335_/X sky130_fd_sc_hd__and3_1
X_6123_ _6123_/CLK _6123_/D VGND VGND VPWR VPWR _6123_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3266_ _3254_/X _3831_/A _4048_/B _3882_/C _3299_/B VGND VGND VPWR VPWR _3266_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_58_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5448__B1 _5256_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6205_/CLK _6054_/D VGND VGND VPWR VPWR _6054_/Q sky130_fd_sc_hd__dfxtp_1
X_5005_ _5005_/A VGND VGND VPWR VPWR _5118_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__4120__B1 _4117_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3197_ _3139_/X _3142_/X _3157_/X _3173_/Y _3196_/X VGND VGND VPWR VPWR _3197_/X
+ sky130_fd_sc_hd__o32a_2
XFILLER_38_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3299__C _3537_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5907_ _6104_/Q _4975_/A _5905_/X _5906_/X VGND VGND VPWR VPWR _5907_/X sky130_fd_sc_hd__o211a_1
XFILLER_22_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5838_ _4998_/X _5833_/X _5031_/X _5837_/Y VGND VGND VPWR VPWR _5838_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_14_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3529__A3 _3525_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5769_ _5924_/A VGND VGND VPWR VPWR _5769_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__4187__B1 _4238_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5923__A1 _6105_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6122__D _6122_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5316__A _5316_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_3_5_0_CLK_A clkbuf_3_5_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5151__A2 _4524_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4220__A _4230_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4111__B1 _4110_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4662__A1 _5167_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4890__A _4890_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5986__A _6201_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4965__A2 _4480_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3768__A3 _3767_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5914__B2 _5913_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5375__C1 _5374_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3925__B1 _3924_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6032__D _6032_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3940__A3 _3937_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5678__B1 _5677_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5142__A2 _5138_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5693__A3 _4856_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3120_ _3120_/A VGND VGND VPWR VPWR _3120_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_121_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4653__A1 _4648_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3051_ _3051_/A VGND VGND VPWR VPWR _3051_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5850__B1 _4541_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3861__C1 _3934_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6207__D _6207_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3953_ _3867_/X _3975_/A _3567_/X _3338_/Y _3934_/B VGND VGND VPWR VPWR _3953_/X
+ sky130_fd_sc_hd__a311o_1
X_3884_ _3956_/C VGND VGND VPWR VPWR _4042_/C sky130_fd_sc_hd__buf_2
XANTENNA__3847__C _3847_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5623_ _6170_/Q _6038_/Q _5627_/S VGND VGND VPWR VPWR _5624_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3916__B1 _3915_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3392__A1 _3919_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5554_ _5554_/A VGND VGND VPWR VPWR _6142_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5669__B1 _4642_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3931__A3 _3195_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4505_ _6046_/Q _4190_/X _4242_/X _4504_/Y VGND VGND VPWR VPWR _6046_/D sky130_fd_sc_hd__a2bb2oi_1
X_5485_ _4803_/X _5161_/X _5445_/A _5451_/X _6121_/Q VGND VGND VPWR VPWR _5486_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3582__C _3582_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4436_ _4696_/A VGND VGND VPWR VPWR _5048_/A sky130_fd_sc_hd__clkbuf_4
X_4367_ _4895_/A VGND VGND VPWR VPWR _5188_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__4975__A _4975_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3318_ _3586_/A VGND VGND VPWR VPWR _3814_/A sky130_fd_sc_hd__buf_4
XANTENNA__4892__A1 _5976_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6106_ _6146_/CLK _6106_/D VGND VGND VPWR VPWR _6106_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4298_ _4298_/A VGND VGND VPWR VPWR _4536_/A sky130_fd_sc_hd__buf_2
XFILLER_74_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3249_ _3603_/A VGND VGND VPWR VPWR _3249_/X sky130_fd_sc_hd__buf_4
XFILLER_46_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3090__S _3094_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6037_ _6045_/CLK _6037_/D VGND VGND VPWR VPWR _6037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3710__D_N _3611_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5841__B1 _5822_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6117__D _6117_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4947__A2 _4945_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4215__A _4264_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3476__D _3476_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3907__B1 _3906_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3773__B _3773_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5046__A _5046_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4885__A _5878_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5496__A2_N _4239_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4635__A1 _4864_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4096__C1 _4095_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5427__A3 _5431_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5832__B1 _5819_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3843__C1 _3842_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6027__D _6027_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output112_A _3128_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4938__A2 _4935_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5060__A1 _4668_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4399__B1 _4233_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3667__C _3966_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3610__A2 _3607_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5434__A2_N _5425_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4020__C1 _3934_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3374__A1 _3572_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput106 _3117_/X VGND VGND VPWR VPWR memory_dmem_response_get[26] sky130_fd_sc_hd__buf_2
XANTENNA__5115__A2 _4581_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput117 _3076_/X VGND VGND VPWR VPWR memory_dmem_response_get[7] sky130_fd_sc_hd__buf_2
Xoutput128 _3031_/X VGND VGND VPWR VPWR memory_imem_response_get[17] sky130_fd_sc_hd__buf_2
Xoutput139 _3053_/X VGND VGND VPWR VPWR memory_imem_response_get[29] sky130_fd_sc_hd__buf_2
X_5270_ _5286_/B input3/X VGND VGND VPWR VPWR _5270_/X sky130_fd_sc_hd__or2_1
XFILLER_114_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5666__A3 _4965_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4221_ _4309_/A VGND VGND VPWR VPWR _4986_/A sky130_fd_sc_hd__buf_2
XFILLER_101_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4874__A1 _5240_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3677__A2 _3676_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4152_ _4152_/A _4152_/B _4152_/C VGND VGND VPWR VPWR _4152_/X sky130_fd_sc_hd__or3_1
XFILLER_110_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4083_ _4083_/A _4083_/B _4083_/C VGND VGND VPWR VPWR _4083_/X sky130_fd_sc_hd__or3_1
X_3103_ _6057_/Q _6085_/Q _3105_/S VGND VGND VPWR VPWR _3104_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5823__B1 _5687_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3204__A _3956_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4626__B2 _4625_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3034_ _3056_/S VGND VGND VPWR VPWR _3043_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__3858__B _3876_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5051__A1 _5123_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4985_ _4985_/A VGND VGND VPWR VPWR _5757_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__5051__B2 _4736_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3936_ _3418_/X _4074_/A _3519_/X _3543_/Y _3350_/A VGND VGND VPWR VPWR _3936_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_51_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3601__A2 _3779_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3867_ _3867_/A VGND VGND VPWR VPWR _3867_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4658__A2_N _4536_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3798_ _3363_/X _3652_/Y _4105_/A VGND VGND VPWR VPWR _3798_/Y sky130_fd_sc_hd__o21bai_1
X_5606_ _5606_/A VGND VGND VPWR VPWR _6162_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3593__B _3659_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5537_ _5537_/A _5568_/B VGND VGND VPWR VPWR _5538_/A sky130_fd_sc_hd__and2_1
XFILLER_11_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5106__A2 _5009_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5468_ _5468_/A _5468_/B VGND VGND VPWR VPWR _5469_/A sky130_fd_sc_hd__and2_1
X_4419_ _4584_/A VGND VGND VPWR VPWR _4420_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5657__A3 _5652_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5399_ input9/X _5445_/A _5395_/X _5398_/X _6101_/Q VGND VGND VPWR VPWR _5401_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_101_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4855__D _4855_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4078__C1 _3488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_86_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4617__A1 _4707_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5814__B1 _5735_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4093__A2 _3932_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5290__A1 _5285_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3840__A2 _3837_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput19 memory_dmem_request_put[45] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4148__A3 _4144_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3934__D _3934_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3356__A1 _3293_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input73_A memory_dmem_request_put[99] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4798__A1_N _4715_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4305__B1 _4378_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3108__A1 _6087_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_2_2_0_CLK_A clkbuf_2_3_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5504__A _5504_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4069__C1 _4068_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6150__CLK _6197_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4084__A2 _3581_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5033__B2 _5032_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4770_ _4788_/B _4883_/A _5188_/B _5005_/A VGND VGND VPWR VPWR _5721_/B sky130_fd_sc_hd__o211ai_4
XANTENNA__3595__A1 _3271_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3721_ _4124_/D _3720_/X _3749_/D _3327_/X VGND VGND VPWR VPWR _3721_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_9_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3652_ _3512_/A _4135_/C _3832_/A VGND VGND VPWR VPWR _3652_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4139__A3 _4136_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5887__A3 _5170_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3583_ _3583_/A _3773_/A _3583_/C VGND VGND VPWR VPWR _3583_/X sky130_fd_sc_hd__and3_2
XANTENNA__3898__A2 _3731_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5322_ _6184_/Q _6076_/Q _5328_/S VGND VGND VPWR VPWR _5323_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4956__C _5944_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5253_ _5242_/Y _5245_/X _4393_/X _5252_/Y VGND VGND VPWR VPWR _5253_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_102_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4847__A1 _4843_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4847__B2 _4846_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5184_ _5048_/X _5021_/X _5680_/B _4742_/X _5140_/A VGND VGND VPWR VPWR _5184_/Y
+ sky130_fd_sc_hd__o2111ai_1
X_4204_ _4265_/A VGND VGND VPWR VPWR _4244_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5414__A _5414_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4135_ _4135_/A _4135_/B _4135_/C _3299_/B VGND VGND VPWR VPWR _4135_/X sky130_fd_sc_hd__or4b_1
XFILLER_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4066_ _3499_/X _4135_/C _3305_/A _3438_/B _3860_/A VGND VGND VPWR VPWR _4067_/B
+ sky130_fd_sc_hd__a311o_1
XANTENNA__4075__A2 _3428_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5272__A1 _5570_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_4_4_0_CLK_A clkbuf_4_5_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3017_ _6027_/Q _6159_/Q _3021_/S VGND VGND VPWR VPWR _3018_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3588__B _3588_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5024__A1 _5140_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3035__A0 _6035_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4968_ _4930_/X _4967_/X _4959_/X _4730_/Y VGND VGND VPWR VPWR _4968_/Y sky130_fd_sc_hd__o211ai_1
X_4899_ _4878_/C _4878_/D _4815_/C _5182_/A VGND VGND VPWR VPWR _4899_/X sky130_fd_sc_hd__a211o_1
X_3919_ _3919_/A VGND VGND VPWR VPWR _3919_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_20_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6023__CLK _6155_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3889__A2 _3888_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3109__A _3109_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6130__D _6130_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4838__A1 _4480_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5909__A2_N _4715_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6173__CLK _6176_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4066__A2 _4135_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3779__A _3983_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3813__A2 _3812_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3026__A0 _6031_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4403__A _5240_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5869__A3 _4931_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6040__D _6040_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4829__A1 _4878_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3501__A1 _3499_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5254__A1 _5229_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4057__A2 _3787_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5940_ _5643_/A _4501_/X _5905_/X _5125_/A VGND VGND VPWR VPWR _5940_/X sky130_fd_sc_hd__a211o_1
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3804__A2 _4044_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3201__B _3442_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5871_ _5862_/Y _5865_/Y _5870_/Y _4494_/X VGND VGND VPWR VPWR _5871_/X sky130_fd_sc_hd__a22o_1
XFILLER_61_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3017__A0 _6027_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4822_ _4362_/X _4363_/A _4937_/D _5118_/B _4364_/X VGND VGND VPWR VPWR _4822_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5557__A2 _5260_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4753_ _5211_/A VGND VGND VPWR VPWR _5761_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__3568__B2 _4092_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3568__A1 _3968_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6046__CLK _6205_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3704_ _3462_/B _3592_/A _3876_/B _3468_/B VGND VGND VPWR VPWR _3704_/X sky130_fd_sc_hd__o211a_2
XANTENNA__4313__A _4313_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5409__A _6102_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4684_ _4685_/A VGND VGND VPWR VPWR _4952_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__4517__B1 _5805_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3635_ _4124_/C _3634_/X _3838_/A VGND VGND VPWR VPWR _3635_/X sky130_fd_sc_hd__o21ba_1
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3566_ _3802_/B _3870_/A VGND VGND VPWR VPWR _3998_/A sky130_fd_sc_hd__nor2_2
XANTENNA__5190__B1 _5022_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6196__CLK _6196_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4628__A1_N _6047_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3740__A1 _3761_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3497_ _3299_/A _3362_/Y _3305_/A _3571_/A VGND VGND VPWR VPWR _3497_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3871__B _3871_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5305_ _5305_/A VGND VGND VPWR VPWR _6068_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5236_ _4957_/X _5233_/Y _5234_/X _5235_/X VGND VGND VPWR VPWR _5236_/Y sky130_fd_sc_hd__o2bb2ai_1
X_5167_ _5167_/A VGND VGND VPWR VPWR _5167_/X sky130_fd_sc_hd__buf_4
XFILLER_84_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5245__A1 _4541_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5098_ _5098_/A VGND VGND VPWR VPWR _5098_/X sky130_fd_sc_hd__buf_2
X_4118_ _3403_/X _3815_/C _3374_/X VGND VGND VPWR VPWR _4118_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_83_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4049_ _3347_/X _3553_/X _4048_/X VGND VGND VPWR VPWR _4049_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4453__C1 _4854_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3749__D _3749_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6125__D _6125_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3008__A0 _6023_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4756__B1 _4536_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3559__A1 _3438_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5319__A _5365_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5181__B1 _5687_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3781__B _3781_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5989__A _5989_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4893__A _5228_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input36_A memory_dmem_request_put[62] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5236__B2 _5235_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5501__B _5501_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3798__A1 _3363_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5787__A2 _5785_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5220__C _5220_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3302__A _3806_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3659__D _3659_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6069__CLK _6074_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6035__D _6035_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4995__B1 _4241_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5539__A2 _4341_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3956__B _3956_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4762__A3 _4923_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4427__A2_N _4293_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3970__A1 _3764_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3970__B2 _3975_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5172__B1 _4420_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3420_ _4036_/A _3838_/A _3420_/C VGND VGND VPWR VPWR _3420_/Y sky130_fd_sc_hd__nor3_1
XFILLER_98_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3722__A1 _3633_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3351_ _3342_/X _3343_/X _3410_/B _3347_/X _3350_/X VGND VGND VPWR VPWR _3351_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_97_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5899__A _5899_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6070_ _6074_/CLK _6070_/D VGND VGND VPWR VPWR _6070_/Q sky130_fd_sc_hd__dfxtp_1
X_3282_ _3282_/A VGND VGND VPWR VPWR _3815_/A sky130_fd_sc_hd__buf_2
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _5021_/A VGND VGND VPWR VPWR _5021_/X sky130_fd_sc_hd__clkbuf_4
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5227__A1 _5222_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5227__B2 _5226_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3212__A _3513_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5778__A2 _4457_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4308__A _4308_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3789__A1 _5388_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4450__A2 _4410_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5923_ _6105_/Q _5772_/A _5905_/A _5922_/X VGND VGND VPWR VPWR _5924_/B sky130_fd_sc_hd__o211a_1
X_5854_ _4668_/A _4296_/X _4960_/A _4879_/A _4928_/A VGND VGND VPWR VPWR _5854_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4805_ input14/X _4717_/X _4718_/X input22/X _4804_/X VGND VGND VPWR VPWR _4805_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3866__B _3918_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5785_ _5102_/C _4935_/X _5097_/X _4924_/X VGND VGND VPWR VPWR _5785_/X sky130_fd_sc_hd__a31o_2
X_2997_ _2997_/A VGND VGND VPWR VPWR _2997_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4736_ _4369_/A _4296_/X _5867_/C _4621_/A VGND VGND VPWR VPWR _4736_/Y sky130_fd_sc_hd__a31oi_4
XANTENNA__5950__A2 _4799_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4667_ _4855_/D VGND VGND VPWR VPWR _5140_/A sky130_fd_sc_hd__buf_4
XANTENNA__3882__A _4083_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3961__A1 _3508_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4978__A _4978_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3618_ _3643_/A VGND VGND VPWR VPWR _3868_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5702__A2 _4721_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4598_ _4832_/A VGND VGND VPWR VPWR _4946_/A sky130_fd_sc_hd__buf_4
XANTENNA__3713__A1 _3621_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3549_ _3549_/A VGND VGND VPWR VPWR _3549_/X sky130_fd_sc_hd__buf_2
XFILLER_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5293__A_N _6206_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4269__A2 _4268_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5466__A1 input23/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5219_ _5216_/X _5218_/X _4767_/X VGND VGND VPWR VPWR _5220_/B sky130_fd_sc_hd__o21ai_2
X_6199_ _6201_/CLK _6199_/D VGND VGND VPWR VPWR _6199_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5466__B2 input15/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5602__A _5602_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5218__A1 _5170_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4505__A1_N _6046_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3122__A _3122_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4218__A _4218_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_3_1_0_CLK_A clkbuf_3_1_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5926__C1 _5179_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3401__B1 _3350_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5941__A2 _5939_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3952__A1 _3215_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3952__B2 _3876_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5154__B1 _5152_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3792__A _3816_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4103__D _4103_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4901__B1 _4563_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3704__A1 _3462_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_12_0_CLK_A clkbuf_3_6_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5457__A1 _5444_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output142_A _3057_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5209__B2 _4858_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4128__A _4128_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4968__B1 _4959_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3967__A _3967_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3686__B _3746_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3640__B1 _6021_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4366__A2_N _4527_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5393__B1 _4201_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5570_ _6200_/Q _6199_/Q _5570_/C VGND VGND VPWR VPWR _5570_/X sky130_fd_sc_hd__and3b_1
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4521_ _4800_/A VGND VGND VPWR VPWR _5715_/A sky130_fd_sc_hd__buf_2
XANTENNA__3943__B2 _3942_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3943__A1 _3286_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4452_ _4533_/A VGND VGND VPWR VPWR _4878_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3403_ _3968_/A VGND VGND VPWR VPWR _3403_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5696__A1 _4422_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5696__B2 _5695_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4499__A2 _4456_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4383_ _4734_/A VGND VGND VPWR VPWR _4815_/D sky130_fd_sc_hd__buf_4
XANTENNA__3207__A _3754_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3334_ _3876_/A VGND VGND VPWR VPWR _4074_/B sky130_fd_sc_hd__buf_2
XFILLER_58_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5448__A1 _6110_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ _6147_/CLK _6122_/D VGND VGND VPWR VPWR _6122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3265_ _3574_/A VGND VGND VPWR VPWR _3299_/B sky130_fd_sc_hd__buf_2
X_6053_ _6196_/CLK _6053_/D VGND VGND VPWR VPWR _6053_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5448__B2 _5260_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5004_ _5004_/A _5731_/B _5973_/B _5004_/D VGND VGND VPWR VPWR _5004_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__4120__A1 _3707_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4120__B2 _4119_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5422__A _5422_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3196_ _3178_/X _3183_/X _3161_/X _3195_/X VGND VGND VPWR VPWR _3196_/X sky130_fd_sc_hd__o211a_1
XFILLER_26_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5081__C1 _4957_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5906_ input12/X _5395_/A _5529_/A _5403_/X VGND VGND VPWR VPWR _5906_/X sky130_fd_sc_hd__a211o_1
X_5837_ _5834_/X _5836_/Y _4345_/X VGND VGND VPWR VPWR _5837_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__5908__C1 _5769_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3088__S _3094_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4187__A1 _4520_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5768_ _6113_/Q _5643_/A _5767_/X VGND VGND VPWR VPWR _5768_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5384__B1 _5376_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5923__A2 _5772_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4719_ input13/X _4717_/X _4718_/X input21/X _4978_/A VGND VGND VPWR VPWR _4719_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5136__B1 _5135_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5699_ _5691_/Y _5698_/Y _5725_/C VGND VGND VPWR VPWR _5699_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4501__A _4501_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3117__A _3117_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4220__B _4220_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4111__A1 _3967_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5332__A _5332_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4662__A2 _4672_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4890__B _4890_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5986__B _6198_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3787__A _4088_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3622__B1 _3281_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6107__CLK _6147_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5375__B1 _6011_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3925__A1 _3195_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4411__A _4442_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5678__A1 _6110_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4886__C1 _4885_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5142__A3 _4494_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3689__B1 _3688_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3027__A _3027_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3050_ _6042_/Q _6174_/Q _3054_/S VGND VGND VPWR VPWR _3051_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4653__A2 _4581_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5850__A1 _4726_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3861__B1 _3720_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5063__C1 _5005_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3952_ _3215_/X _3359_/C _3762_/X _3876_/X _3701_/X VGND VGND VPWR VPWR _3952_/Y
+ sky130_fd_sc_hd__o221ai_1
X_3883_ _4149_/B _3520_/X _3762_/A _3710_/C VGND VGND VPWR VPWR _3883_/X sky130_fd_sc_hd__o22a_1
X_5622_ _5622_/A VGND VGND VPWR VPWR _6169_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3916__A1 _3645_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3377__C1 _3376_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5553_ _5988_/A _5553_/B VGND VGND VPWR VPWR _5554_/A sky130_fd_sc_hd__or2_1
X_4504_ _4504_/A _4504_/B _4974_/C VGND VGND VPWR VPWR _4504_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__5417__A _6104_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4321__A _4942_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5669__A1 _5190_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3392__A2 _4083_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5484_ _5484_/A _5528_/B VGND VGND VPWR VPWR _6120_/D sky130_fd_sc_hd__nand2_1
X_4435_ _4926_/B VGND VGND VPWR VPWR _4437_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_6_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4366_ _4527_/C _4527_/D _4601_/A _4602_/A VGND VGND VPWR VPWR _4895_/A sky130_fd_sc_hd__o2bb2ai_2
XFILLER_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4892__A2 _4840_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3317_ _3779_/C VGND VGND VPWR VPWR _4089_/B sky130_fd_sc_hd__clkbuf_4
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6105_ _6145_/CLK _6105_/D VGND VGND VPWR VPWR _6105_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5152__A _5152_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4297_ _4527_/A VGND VGND VPWR VPWR _4297_/X sky130_fd_sc_hd__buf_2
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3248_ _3315_/A _3436_/B VGND VGND VPWR VPWR _3603_/A sky130_fd_sc_hd__nand2_2
XFILLER_74_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ _6202_/CLK _6036_/D VGND VGND VPWR VPWR _6036_/Q sky130_fd_sc_hd__dfxtp_1
X_3179_ _3443_/B VGND VGND VPWR VPWR _3330_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__3852__B1 _3301_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5841__B2 _5840_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5841__A1 _6189_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5054__C1 _4937_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5298__S _5306_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4947__A3 _5018_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3604__B1 _3603_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3400__A _4074_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6133__D _6133_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5357__A0 _6061_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3907__A1 _3904_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5742__A1_N _4999_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5109__B1 _5050_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4826__A2_N _4822_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5327__A _5327_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3773__C _3773_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4231__A _4231_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5046__B _5444_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4885__B _5118_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5062__A _5062_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4096__B1 _3707_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4635__A2 _5188_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5832__A1 _5263_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3843__B1 _3699_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4399__A1 _4266_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4406__A _4860_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5060__A2 _5000_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4399__B2 _6135_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3310__A _3614_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output105_A _3115_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5348__A0 _6059_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6043__D _6043_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5237__A _5237_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4020__B1 _3489_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3374__A2 _4073_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput107 _3120_/X VGND VGND VPWR VPWR memory_dmem_response_get[27] sky130_fd_sc_hd__buf_2
Xoutput118 _3078_/X VGND VGND VPWR VPWR memory_dmem_response_get[8] sky130_fd_sc_hd__buf_2
Xoutput129 _3033_/X VGND VGND VPWR VPWR memory_imem_response_get[18] sky130_fd_sc_hd__buf_2
X_4220_ _4230_/A _4220_/B _4220_/C _4220_/D VGND VGND VPWR VPWR _4309_/A sky130_fd_sc_hd__nand4_4
XANTENNA__4874__A2 _4581_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3531__C1 _3530_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4151_ _3350_/X _4105_/C _4149_/X _4150_/Y _3862_/A VGND VGND VPWR VPWR _4151_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4082_ _3831_/A _4124_/D _3249_/X _4124_/C _3756_/X VGND VGND VPWR VPWR _4082_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__4087__B1 _3707_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3102_ _3102_/A VGND VGND VPWR VPWR _3102_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_110_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5823__A1 _4754_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3204__B _3632_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3033_ _3033_/A VGND VGND VPWR VPWR _3033_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5036__C1 _5035_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3220__A _3461_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4316__A _5235_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4984_ _4984_/A VGND VGND VPWR VPWR _4984_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4035__B _4061_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5051__A2 _4735_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3935_ _3695_/A _3931_/Y _3933_/X _3934_/Y _3577_/X VGND VGND VPWR VPWR _3935_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_32_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5339__A0 _6056_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5605_ _6162_/Q _6030_/Q _5605_/S VGND VGND VPWR VPWR _5606_/A sky130_fd_sc_hd__mux2_1
X_3866_ _3918_/A _3918_/C _3918_/B VGND VGND VPWR VPWR _3866_/X sky130_fd_sc_hd__or3_2
XANTENNA__4547__D1 _4673_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3797_ _3797_/A VGND VGND VPWR VPWR _4105_/A sky130_fd_sc_hd__buf_2
XANTENNA__4011__B1 _6038_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3593__C _3614_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_4_0_0_CLK_A clkbuf_4_1_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5536_ input5/X VGND VGND VPWR VPWR _5568_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__4986__A _4986_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5467_ _4977_/X _5433_/A _5805_/C _5451_/X _6115_/Q VGND VGND VPWR VPWR _5468_/A
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3770__C1 _3769_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4418_ _5148_/D _5976_/A _4957_/A _4369_/Y VGND VGND VPWR VPWR _4418_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5581__S _5583_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5511__B1 _5425_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5398_ _5503_/A VGND VGND VPWR VPWR _5398_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4349_ _4769_/A VGND VGND VPWR VPWR _4350_/A sky130_fd_sc_hd__buf_2
XFILLER_99_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4078__B1 _3919_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4617__A2 _4619_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5814__A1 _5813_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6019_ _6155_/CLK _6019_/D VGND VGND VPWR VPWR _6019_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6128__D _6128_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3825__B1 _3562_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5290__A2 _5286_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5027__C1 _5782_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4226__A _5438_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3130__A _3301_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4250__B1 _5756_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3356__A2 _3300_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5750__B1 _5729_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4896__A _4926_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input66_A memory_dmem_request_put[92] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4305__A1 _4347_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3305__A _3305_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4069__B1 _3938_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6038__D _6038_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4084__A3 _3703_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5520__A _5520_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3959__B _3959_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3040__A _3040_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3720_ _3720_/A VGND VGND VPWR VPWR _3720_/X sky130_fd_sc_hd__buf_2
XANTENNA__3975__A _3975_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3595__A2 _3594_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3651_ _3711_/A VGND VGND VPWR VPWR _3832_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5741__B1 _4883_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3582_ _3686_/A _3582_/B _3582_/C VGND VGND VPWR VPWR _3583_/A sky130_fd_sc_hd__and3_2
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5321_ _5321_/A VGND VGND VPWR VPWR _6075_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5252_ _4765_/X _5249_/X _5251_/X _4950_/X VGND VGND VPWR VPWR _5252_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__4847__A2 _4833_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_87_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4956__D _4956_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5183_ _5745_/A _4777_/X _4778_/X _5903_/D _5170_/X VGND VGND VPWR VPWR _5183_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__3504__C1 _3724_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4203_ input1/X VGND VGND VPWR VPWR _4282_/A sky130_fd_sc_hd__inv_2
XANTENNA__5414__B _5422_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3215__A _3710_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4134_ _4127_/Y _4133_/X _3286_/X VGND VGND VPWR VPWR _4134_/X sky130_fd_sc_hd__a21o_1
XFILLER_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4065_ _4065_/A _4065_/B _4092_/C _3495_/X VGND VGND VPWR VPWR _4067_/A sky130_fd_sc_hd__or4b_1
XANTENNA__5272__A2 input3/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5430__A _5430_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3016_ _3016_/A VGND VGND VPWR VPWR _3016_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3588__C _3588_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5024__A2 _5020_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3035__A1 _6167_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4967_ _4967_/A VGND VGND VPWR VPWR _4967_/X sky130_fd_sc_hd__clkbuf_4
X_4898_ _5240_/A _5240_/D _5878_/B _4897_/Y VGND VGND VPWR VPWR _4898_/Y sky130_fd_sc_hd__a31oi_4
XANTENNA__5980__B1 _5979_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3918_ _3918_/A _3918_/B _3918_/C _3538_/A VGND VGND VPWR VPWR _3918_/X sky130_fd_sc_hd__or4b_2
XANTENNA__3991__C1 _3990_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3849_ _4092_/A _3711_/A _3719_/B _3647_/A VGND VGND VPWR VPWR _3849_/X sky130_fd_sc_hd__a31o_1
XFILLER_20_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5519_ _5519_/A _5531_/B VGND VGND VPWR VPWR _5520_/A sky130_fd_sc_hd__and2_1
XFILLER_105_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4299__B1 _6134_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4838__A2 _4437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4066__A3 _3305_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5799__B1 _5798_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5340__A _5340_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3779__B _3983_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3026__A1 _6163_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4223__B1 _4222_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5184__D1 _5140_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5723__B1 _4950_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5515__A _5515_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4829__A2 _4551_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3501__A2 _3911_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5254__A2 _5238_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4057__A3 _4056_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5870_ _5794_/Y _5866_/X _5868_/Y _5869_/Y VGND VGND VPWR VPWR _5870_/Y sky130_fd_sc_hd__o22ai_4
XANTENNA__3804__A3 _3801_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4821_ _4369_/A _4480_/C _4820_/Y VGND VGND VPWR VPWR _4821_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__5557__A3 _5431_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3017__A1 _6159_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4752_ _4750_/Y _4652_/A _4751_/Y _4316_/X VGND VGND VPWR VPWR _4752_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3568__A2 _3932_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5962__B1 _5960_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3703_ _3703_/A VGND VGND VPWR VPWR _3910_/C sky130_fd_sc_hd__clkbuf_2
X_4683_ _4665_/X _4677_/Y _4682_/X VGND VGND VPWR VPWR _4683_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5409__B _5425_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3634_ _3343_/A _3631_/X _3756_/A _3633_/Y VGND VGND VPWR VPWR _3634_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5714__B1 _5705_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4517__A1 _4716_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5190__A1 _4347_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3565_ _3858_/A VGND VGND VPWR VPWR _3932_/B sky130_fd_sc_hd__buf_2
XANTENNA__5425__A _6106_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3496_ _3968_/A _3494_/X _3495_/X VGND VGND VPWR VPWR _3496_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__3740__A2 _4149_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3871__C _3904_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5304_ _6192_/Q _6068_/Q _5306_/S VGND VGND VPWR VPWR _5305_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5235_ _5235_/A VGND VGND VPWR VPWR _5235_/X sky130_fd_sc_hd__buf_4
XANTENNA__5478__C1 _5477_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4150__C1 _3574_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5166_ _5166_/A _5166_/B VGND VGND VPWR VPWR _5166_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5097_ _5899_/C VGND VGND VPWR VPWR _5097_/X sky130_fd_sc_hd__clkbuf_4
X_4117_ _4116_/X _3699_/A _3849_/X _4102_/A VGND VGND VPWR VPWR _4117_/Y sky130_fd_sc_hd__a31oi_2
XANTENNA__5160__A _5822_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5245__A2 _4464_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4048_ _4048_/A _4048_/B _4065_/B VGND VGND VPWR VPWR _4048_/X sky130_fd_sc_hd__or3_1
XFILLER_44_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4453__B1 _4878_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5650__C1 _5649_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5999_ _5999_/A _5999_/B _6014_/B VGND VGND VPWR VPWR _6000_/A sky130_fd_sc_hd__and3_1
XANTENNA__3008__A1 _6155_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4756__A1 _4273_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5953__B1 _5952_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4504__A _4504_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3559__A2 _3558_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3964__C1 _3512_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6141__D _6141_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5705__B1 _4950_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6140__CLK _6146_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5181__A1 _4777_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3781__C _3781_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input29_A memory_dmem_request_put[55] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5787__A3 _5786_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3798__A2 _3652_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4995__B2 _4994_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5539__A3 _4802_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4414__A _4414_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3956__C _3956_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3955__C1 _3299_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6051__D _6051_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3944__A1_N _3866_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3970__A2 _3965_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5172__A1 _5973_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output97_A _3100_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3722__A2 _4073_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3350_ _3350_/A VGND VGND VPWR VPWR _3350_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_112_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5020_ _5020_/A VGND VGND VPWR VPWR _5020_/X sky130_fd_sc_hd__buf_4
X_3281_ _3281_/A VGND VGND VPWR VPWR _3934_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__4132__C1 _3707_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5899__B _5899_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4683__B1 _4682_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5227__A2 _4630_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3789__A2 _6027_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5922_ input13/X _5420_/A _5163_/A _4984_/A VGND VGND VPWR VPWR _5922_/X sky130_fd_sc_hd__a211o_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5853_ _5745_/C _5899_/B _5240_/D _4918_/A VGND VGND VPWR VPWR _5853_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4450__A3 _4418_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5935__B1 _5102_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5784_ _5778_/X _5781_/X _5754_/Y _5783_/Y VGND VGND VPWR VPWR _5784_/Y sky130_fd_sc_hd__a22oi_4
X_4804_ _4804_/A VGND VGND VPWR VPWR _4804_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3866__C _3918_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4735_ _5211_/A _4873_/A _5182_/A VGND VGND VPWR VPWR _4735_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__6163__CLK _6197_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2996_ _6018_/Q _6150_/Q _2998_/S VGND VGND VPWR VPWR _2997_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4666_ _4666_/A VGND VGND VPWR VPWR _5004_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3961__A2 _3951_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4597_ _4926_/C VGND VGND VPWR VPWR _5867_/C sky130_fd_sc_hd__buf_2
X_3617_ _3754_/A VGND VGND VPWR VPWR _3643_/A sky130_fd_sc_hd__buf_2
XANTENNA__3882__B _3882_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5438__A_N _5392_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3713__A2 _3709_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3548_ _3571_/A VGND VGND VPWR VPWR _3548_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_115_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3299__D_N _3491_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3479_ _4036_/A VGND VGND VPWR VPWR _3479_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4994__A input6/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5466__A2 _5437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5218_ _5170_/X _5680_/B _4679_/X _4584_/X _5217_/X VGND VGND VPWR VPWR _5218_/X
+ sky130_fd_sc_hd__o311a_1
X_6198_ _6201_/CLK _6198_/D VGND VGND VPWR VPWR _6198_/Q sky130_fd_sc_hd__dfxtp_1
X_5149_ _5147_/Y _5148_/Y _4744_/X VGND VGND VPWR VPWR _5150_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__3403__A _3968_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5218__A2 _5680_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6136__D _6136_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4218__B _4218_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3743__A2_N _3738_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4234__A _4234_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5926__B1 _4930_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3401__A1 _3830_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3952__A2 _3359_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5154__A1 _5018_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3792__B _3806_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4901__A1 _4899_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3704__A2 _3592_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5457__A2 _5445_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_85_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output135_A _3044_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6036__CLK _6202_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3313__A _3382_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4128__B _4128_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6046__D _6046_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4968__A1 _4930_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5090__B1 _5042_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6186__CLK _6204_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3640__A1 _3625_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2979__B1 _2998_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5917__B1 _5916_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3686__C _3773_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3640__B2 _3541_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3928__C1 _3701_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3983__A _3983_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5393__A1 _5436_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4520_ _4520_/A VGND VGND VPWR VPWR _4800_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3943__A2 _3930_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4451_ _4252_/X _4346_/X _4389_/Y _4393_/X _4450_/Y VGND VGND VPWR VPWR _4504_/A
+ sky130_fd_sc_hd__o311ai_4
X_3402_ _3876_/B VGND VGND VPWR VPWR _3968_/A sky130_fd_sc_hd__buf_2
XANTENNA__5696__A2 _4699_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4382_ _4700_/A VGND VGND VPWR VPWR _4734_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6121_ _6123_/CLK _6121_/D VGND VGND VPWR VPWR _6121_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3333_ _3437_/B VGND VGND VPWR VPWR _3876_/A sky130_fd_sc_hd__clkbuf_2
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3264_ _3754_/A VGND VGND VPWR VPWR _3574_/A sky130_fd_sc_hd__buf_2
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6052_ _6196_/CLK _6052_/D VGND VGND VPWR VPWR _6052_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5448__A2 _5222_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5667_/B _5003_/B _5003_/C _5152_/C VGND VGND VPWR VPWR _5731_/B sky130_fd_sc_hd__nand4_2
XANTENNA__4120__A2 _4115_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5422__B _5422_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3223__A _4065_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3195_ _3195_/A _3195_/B _3194_/X VGND VGND VPWR VPWR _3195_/X sky130_fd_sc_hd__or3b_1
XFILLER_39_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5081__B1 _5080_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5905_ _5905_/A VGND VGND VPWR VPWR _5905_/X sky130_fd_sc_hd__buf_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5836_ _5836_/A _5836_/B VGND VGND VPWR VPWR _5836_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5908__B1 _5907_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3893__A _4149_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4187__A2 _4405_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2979_ _5998_/C _5998_/B _2998_/S VGND VGND VPWR VPWR _2979_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5767_ _5805_/A _5805_/B _5767_/C VGND VGND VPWR VPWR _5767_/X sky130_fd_sc_hd__and3_1
XANTENNA__5384__A1 _5373_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5698_ _5694_/X _5697_/X _5664_/X _4685_/X VGND VGND VPWR VPWR _5698_/Y sky130_fd_sc_hd__a211oi_1
XANTENNA__3395__B1 _3580_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4718_ _4718_/A VGND VGND VPWR VPWR _4718_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4649_ _4649_/A VGND VGND VPWR VPWR _5899_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__5136__A1 _5102_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4220__C _4220_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6059__CLK _6207_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5613__A _5613_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4111__A2 _3495_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3133__A _3918_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4890__C _4890_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5072__B1 _4494_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3622__A1 _3157_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5375__A1 _5368_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4583__C1 _4582_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3925__A2 _3831_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3308__A _3308_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5678__A2 _4721_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4886__B1 _4882_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3689__A1 _3658_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5523__A _5715_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_67_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4653__A3 _4650_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5850__A2 _5706_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3861__A1 _3911_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3861__B2 _4124_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5063__B1 _4697_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3951_ _3139_/X _3946_/X _3947_/Y _3950_/X VGND VGND VPWR VPWR _3951_/X sky130_fd_sc_hd__o31a_1
XFILLER_51_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3882_ _4083_/A _3882_/B _3882_/C VGND VGND VPWR VPWR _3882_/X sky130_fd_sc_hd__and3_1
X_5621_ _6169_/Q _6037_/Q _5627_/S VGND VGND VPWR VPWR _5622_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4602__A _4602_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3916__A2 _4143_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3377__B1 _3369_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5552_ _5256_/A _4218_/C _5260_/A _6142_/Q _5482_/X VGND VGND VPWR VPWR _5553_/B
+ sky130_fd_sc_hd__o32a_1
X_4503_ _4503_/A VGND VGND VPWR VPWR _4974_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__5417__B _5425_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5669__A2 _5667_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3218__A _3700_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3392__A3 _3893_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5483_ _5482_/X _6120_/Q _5445_/A _5131_/Y VGND VGND VPWR VPWR _5484_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__6201__CLK _6201_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4434_ _4890_/C VGND VGND VPWR VPWR _5712_/C sky130_fd_sc_hd__buf_4
XFILLER_113_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4365_ _4769_/C VGND VGND VPWR VPWR _4369_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_98_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3316_ _3956_/C VGND VGND VPWR VPWR _3779_/C sky130_fd_sc_hd__buf_2
XFILLER_86_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4892__A3 _4891_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6104_ _6146_/CLK _6104_/D VGND VGND VPWR VPWR _6104_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5433__A _5433_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5152__B _5152_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5826__C1 _4879_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4296_ _5744_/A VGND VGND VPWR VPWR _4296_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_86_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _6197_/CLK _6035_/D VGND VGND VPWR VPWR _6035_/Q sky130_fd_sc_hd__dfxtp_1
X_3247_ _3311_/B _3461_/B VGND VGND VPWR VPWR _3436_/B sky130_fd_sc_hd__nor2_2
XFILLER_73_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3178_ _3780_/C _3468_/A VGND VGND VPWR VPWR _3178_/X sky130_fd_sc_hd__or2_4
XANTENNA__3852__A1 _4128_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5841__A2 _4629_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5579__S _5583_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5054__B1 _4937_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3604__A1 _3549_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3099__S _3105_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6003__C1 _6002_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5819_ _5819_/A VGND VGND VPWR VPWR _5905_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5357__A1 _6092_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3907__A2 _3464_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5109__A1 _5140_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5762__D1 _5152_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5109__B2 _5048_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3128__A _3128_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4231__B _4231_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4868__B1 _4698_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4885__C _5079_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5739__A2_N _5737_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3540__B1 _3539_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5343__A _5343_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4096__A1 _3340_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4995__A2_N _4991_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3843__A1 _3594_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5832__A2 _4501_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input11_A memory_dmem_request_put[37] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4399__A2 _4272_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5060__A3 _5118_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5348__A1 _6088_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4422__A _4422_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4020__A1 _3195_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3374__A3 _4152_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3038__A _3038_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput119 _3080_/X VGND VGND VPWR VPWR memory_dmem_response_get[9] sky130_fd_sc_hd__buf_2
Xoutput108 _3122_/X VGND VGND VPWR VPWR memory_dmem_response_get[28] sky130_fd_sc_hd__buf_2
XANTENNA__4874__A3 _5903_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4150_ _3668_/X _3549_/X _3831_/A _3603_/X _3574_/X VGND VGND VPWR VPWR _4150_/Y
+ sky130_fd_sc_hd__a311oi_1
XANTENNA__3531__B1 _3516_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5249__A1_N _4547_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput90 _3084_/X VGND VGND VPWR VPWR memory_dmem_response_get[11] sky130_fd_sc_hd__buf_2
X_3101_ _6056_/Q _6084_/Q _3105_/S VGND VGND VPWR VPWR _3102_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4087__A1 _3749_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4081_ _4072_/X _4080_/Y _3821_/X _6041_/Q _3891_/X VGND VGND VPWR VPWR _6041_/D
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5823__A2 _5745_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3032_ _6034_/Q _6166_/Q _3032_/S VGND VGND VPWR VPWR _3033_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5036__B1 _5031_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4983_ _4974_/Y _4982_/X _6052_/Q _4190_/X VGND VGND VPWR VPWR _6052_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4035__C _4035_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3934_ _3975_/A _3934_/B _3934_/C _3934_/D VGND VGND VPWR VPWR _3934_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__3598__B1 _3539_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3865_ _4039_/B _3799_/X _3522_/X _3975_/C _3508_/A VGND VGND VPWR VPWR _3865_/Y
+ sky130_fd_sc_hd__a221oi_1
XANTENNA__5339__A1 _6084_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4332__A _4414_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4547__C1 _5118_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5817__A1_N _6188_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5604_ _5604_/A VGND VGND VPWR VPWR _6161_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__5428__A _5508_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3796_ _3792_/X _3795_/Y _3727_/X _6028_/Q _3728_/X VGND VGND VPWR VPWR _6028_/D
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4011__A1 _4002_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4011__B2 _3822_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3593__D _3593_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4135__D_N _3299_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5535_ _5523_/X _4333_/A _5529_/X _5491_/X _6137_/Q VGND VGND VPWR VPWR _5537_/A
+ sky130_fd_sc_hd__a32o_1
X_5466_ input23/X _5437_/A _5439_/A input15/X VGND VGND VPWR VPWR _5805_/C sky130_fd_sc_hd__a22o_1
XANTENNA__3770__B1 _3763_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4417_ _5029_/A VGND VGND VPWR VPWR _4957_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5511__A1 _5093_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5397_ _5499_/A VGND VGND VPWR VPWR _5503_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5163__A _5163_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4348_ _4759_/A VGND VGND VPWR VPWR _4769_/A sky130_fd_sc_hd__buf_2
XANTENNA_input3_A EN_memory_imem_request_put VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4279_ _4379_/A VGND VGND VPWR VPWR _4860_/B sky130_fd_sc_hd__buf_2
XFILLER_100_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4078__B2 _3428_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4078__A1 _3679_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5814__A2 _4964_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6018_ _6155_/CLK _6018_/D VGND VGND VPWR VPWR _6018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3825__A1 _3775_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5027__B1 _4739_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3411__A _3870_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4507__A _5648_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4250__A1 _4243_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6144__D _6144_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5033__A2_N _5062_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5338__A _5338_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5750__B2 _5749_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4305__A2 _4296_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input59_A memory_dmem_request_put[85] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5073__A _5073_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4710__C1 _4709_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3305__B _3343_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4069__A1 _3626_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5266__B1 _4224_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4417__A _5029_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3321__A _3754_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3959__C _4146_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4242__A2_N _4237_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6054__D _6054_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3975__B _3975_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3595__A3 _3249_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3650_ _3781_/C VGND VGND VPWR VPWR _3711_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__4152__A _4152_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5741__A1 _4649_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3581_ _3581_/A VGND VGND VPWR VPWR _4124_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5320_ _6183_/Q _6075_/Q _5328_/S VGND VGND VPWR VPWR _5321_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3752__B1 _6025_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5251_ _5755_/C _4369_/Y _5010_/X _4395_/A _5250_/X VGND VGND VPWR VPWR _5251_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__3504__B1 _3497_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4202_ _4976_/A VGND VGND VPWR VPWR _5044_/A sky130_fd_sc_hd__clkbuf_2
X_5182_ _5182_/A VGND VGND VPWR VPWR _5903_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_96_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4133_ _4061_/X _3904_/X _4128_/Y _4132_/X VGND VGND VPWR VPWR _4133_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5711__A _5711_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4064_ _4058_/Y _4060_/X _3699_/X _4063_/X _3508_/A VGND VGND VPWR VPWR _4064_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_56_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3015_ _6026_/Q _6158_/Q _3021_/S VGND VGND VPWR VPWR _3016_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4327__A _4527_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4768__C1 _4767_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5024__A3 _5021_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4966_ _4524_/X _4431_/X _4965_/Y VGND VGND VPWR VPWR _4966_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_51_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4897_ _4483_/X _4485_/X _4945_/A _5096_/A VGND VGND VPWR VPWR _4897_/Y sky130_fd_sc_hd__o22ai_4
XANTENNA__5980__A1 _4836_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5980__B2 _5961_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3917_ _3815_/B _3910_/X _4036_/C _3628_/A _3916_/X VGND VGND VPWR VPWR _3917_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3991__B1 _3643_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3848_ _3343_/X _3881_/B _3195_/A _3847_/X VGND VGND VPWR VPWR _3848_/X sky130_fd_sc_hd__a31o_1
XFILLER_22_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3443__A_N _3461_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3779_ _3983_/A _3983_/B _3779_/C VGND VGND VPWR VPWR _4116_/A sky130_fd_sc_hd__and3_2
XANTENNA__3743__B1 _3742_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5518_ _5495_/X _4908_/X _5498_/X _6131_/Q _5503_/A VGND VGND VPWR VPWR _5519_/A
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5592__S _5594_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4299__A1 _4268_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3406__A _3406_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5449_ _5444_/X _5445_/X _5677_/C _5447_/X _5448_/X VGND VGND VPWR VPWR _6110_/D
+ sky130_fd_sc_hd__a311o_1
XANTENNA__5496__B1 _5495_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3593__A_N _4073_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4838__A3 _4865_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6139__D _6139_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5248__B1 _5152_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5799__A1 _5732_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3779__C _3779_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3141__A _3707_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2980__A _6178_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4223__A1 _4199_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5068__A _5152_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3431__C1 _3653_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5184__C1 _4742_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5723__A1 _5719_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4700__A _4700_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3734__B1 _3680_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3316__A _3956_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6049__D _6049_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5239__B1 _4547_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5531__A _5531_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3051__A _3051_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4820_ _4929_/B _4929_/A _4942_/A VGND VGND VPWR VPWR _4820_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__5411__B1 _5410_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _4488_/X _5021_/A _4956_/A VGND VGND VPWR VPWR _4751_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3568__A3 _3567_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5962__B2 _5961_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5962__A1 _5959_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3702_ _3773_/B VGND VGND VPWR VPWR _3703_/A sky130_fd_sc_hd__clkbuf_4
X_4682_ _4679_/X _4619_/X _4657_/X _4681_/Y _5734_/A VGND VGND VPWR VPWR _4682_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3973__B1 _6036_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3633_ _3633_/A _3710_/C VGND VGND VPWR VPWR _3633_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__5714__A1 _4570_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4517__A2 _4513_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5706__A _5706_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5714__B2 _5713_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3725__B1 _3724_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4610__A _5188_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5190__A2 _4673_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3564_ _3499_/A _4065_/A _3799_/A _3528_/A VGND VGND VPWR VPWR _3564_/X sky130_fd_sc_hd__a31o_1
X_3495_ _3621_/D VGND VGND VPWR VPWR _3495_/X sky130_fd_sc_hd__buf_4
XANTENNA__5425__B _5425_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5478__B1 _5540_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5303_ _5303_/A VGND VGND VPWR VPWR _6067_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3226__A _3226_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5234_ _5018_/B _5755_/D _4945_/X _5829_/A _4652_/A VGND VGND VPWR VPWR _5234_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_69_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4150__B1 _3603_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6092__CLK _6204_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5165_ _6121_/Q _4511_/X _5013_/X _5164_/X VGND VGND VPWR VPWR _5166_/B sky130_fd_sc_hd__o211a_1
XFILLER_96_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4116_ _4116_/A _4116_/B _3911_/A VGND VGND VPWR VPWR _4116_/X sky130_fd_sc_hd__or3b_1
X_5096_ _5096_/A VGND VGND VPWR VPWR _5102_/D sky130_fd_sc_hd__buf_2
XFILLER_96_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4453__A1 _4878_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5245__A3 _5243_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4047_ _3477_/X _4036_/X _4039_/Y _4046_/Y _3744_/A VGND VGND VPWR VPWR _4047_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5650__B1 _5676_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5998_ _5998_/A _5998_/B _5998_/C _6201_/Q VGND VGND VPWR VPWR _5999_/B sky130_fd_sc_hd__nand4_1
X_4949_ _4943_/Y _4944_/X _4947_/X _5973_/B VGND VGND VPWR VPWR _4949_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__4756__A2 _4211_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5953__A1 _5951_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4504__B _4504_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3964__B1 _3687_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3959__A_N _3955_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5705__A1 _5683_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3716__B1 _3418_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5181__A2 _4778_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4520__A _4520_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3781__D _3781_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3136__A _3609_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4141__B1 _6044_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5351__A _5351_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2975__A _6197_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4274__A1_N _4266_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5641__B1 _5410_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3955__B1 _3954_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3970__A3 _4105_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5526__A _5526_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4904__C1 _4903_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5172__A2 _5171_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3280_ _3864_/B VGND VGND VPWR VPWR _3281_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4132__B1 _4131_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5899__C _5899_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4683__A1 _4665_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5921_ _4665_/X _4956_/A _5917_/Y _4964_/X _5920_/Y VGND VGND VPWR VPWR _5921_/Y
+ sky130_fd_sc_hd__o311ai_2
XANTENNA__5632__A0 _6174_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5852_ _5079_/A _4534_/X _4572_/X VGND VGND VPWR VPWR _5852_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5935__A1 _5829_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5935__B2 _5167_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5783_ _5712_/D _5176_/X _5782_/X _4874_/X _5752_/Y VGND VGND VPWR VPWR _5783_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_4803_ _5044_/A VGND VGND VPWR VPWR _4803_/X sky130_fd_sc_hd__buf_2
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4734_ _4734_/A VGND VGND VPWR VPWR _5182_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3946__B1 _3945_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2995_ _2995_/A VGND VGND VPWR VPWR _2995_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4665_ _4665_/A VGND VGND VPWR VPWR _4665_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5699__B1 _5725_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5436__A _5436_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4596_ _4573_/X _4583_/Y _4584_/X _4595_/Y VGND VGND VPWR VPWR _4596_/Y sky130_fd_sc_hd__o211ai_4
X_3616_ _3406_/A _4152_/A _3756_/C _3549_/A VGND VGND VPWR VPWR _3616_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4340__A _6138_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3882__C _3882_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4371__B1 _4364_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3547_ _3327_/X _3543_/Y _3476_/A _4036_/B _3546_/X VGND VGND VPWR VPWR _3547_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_115_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4123__B1 _3954_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3478_ _3466_/Y _3476_/X _3477_/X VGND VGND VPWR VPWR _3478_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4994__B _4994_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5217_ _5050_/Y _5944_/D _5074_/X _4556_/A VGND VGND VPWR VPWR _5217_/X sky130_fd_sc_hd__a211o_1
X_6197_ _6197_/CLK _6197_/D VGND VGND VPWR VPWR _6197_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5871__B1 _5870_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5148_ _5148_/A _5148_/B _5148_/C _5148_/D VGND VGND VPWR VPWR _5148_/Y sky130_fd_sc_hd__nand4_1
XFILLER_56_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5079_ _5079_/A _5079_/B _5079_/C VGND VGND VPWR VPWR _5079_/X sky130_fd_sc_hd__and3_1
XANTENNA__5218__A3 _4679_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4218__C _4218_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5623__A0 _6170_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4515__A _4515_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5926__A1 _5028_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3937__B1 _3923_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5926__B2 _5148_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6152__D _6152_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3401__A2 _3410_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5139__C1 _5118_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5154__A2 _4840_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3792__C _3792_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5572__A1_N _6199_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4901__A2 _4900_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4114__B1 _4113_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input41_A memory_dmem_request_put[67] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5457__A3 _5455_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_85_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5862__B1 _5861_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_85_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output128_A _3031_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5614__A0 _6166_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4968__A2 _4967_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5090__A1 input27/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4425__A _4566_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5090__B2 input11/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2979__A1 _5998_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5917__A1 _5123_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3686__D _3802_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3640__A2 _3639_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3928__B1 _3847_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6062__D _6062_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3983__B _3983_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5393__A2 _5392_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3943__A3 _3935_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5256__A _5256_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4450_ _4732_/B _4410_/Y _4418_/X _4420_/X _4449_/Y VGND VGND VPWR VPWR _4450_/Y
+ sky130_fd_sc_hd__o311ai_4
XFILLER_7_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4381_ _4578_/A VGND VGND VPWR VPWR _4883_/A sky130_fd_sc_hd__clkbuf_4
X_3401_ _3830_/D _3410_/B _3350_/X VGND VGND VPWR VPWR _3401_/Y sky130_fd_sc_hd__o21ai_1
X_3332_ _3663_/A VGND VGND VPWR VPWR _4074_/A sky130_fd_sc_hd__clkbuf_2
X_6120_ _6145_/CLK _6120_/D VGND VGND VPWR VPWR _6120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3263_ _3468_/B VGND VGND VPWR VPWR _3882_/C sky130_fd_sc_hd__buf_2
XFILLER_39_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6051_ _6205_/CLK _6051_/D VGND VGND VPWR VPWR _6051_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5853__B1 _4918_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5002_ _4997_/Y _4789_/X _4461_/X _4998_/X _5001_/X VGND VGND VPWR VPWR _5002_/Y
+ sky130_fd_sc_hd__o2111ai_4
X_3194_ _4089_/A VGND VGND VPWR VPWR _3194_/X sky130_fd_sc_hd__buf_2
XFILLER_39_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5605__A0 _6162_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6130__CLK _6207_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5081__A1 _4661_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3616__C1 _3549_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5081__B2 _5021_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5904_ _4794_/X _5903_/X _5982_/C _5125_/A VGND VGND VPWR VPWR _5955_/A sky130_fd_sc_hd__o211a_2
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3092__A0 _6188_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5835_ _5867_/C _4945_/A _4353_/A _4882_/A VGND VGND VPWR VPWR _5836_/B sky130_fd_sc_hd__a31o_1
XANTENNA__5908__A1 _5902_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5369__C1 _6143_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3893__B _3932_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5766_ _5175_/X _5760_/Y _5765_/Y _5725_/C VGND VGND VPWR VPWR _5766_/Y sky130_fd_sc_hd__o211ai_4
XANTENNA__4187__A3 _4859_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2978_ _5985_/B VGND VGND VPWR VPWR _2998_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__5384__A2 _5371_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5697_ _4870_/X _4440_/Y _4967_/X _5696_/Y _4679_/X VGND VGND VPWR VPWR _5697_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3395__A1 _3377_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4717_ _4717_/A VGND VGND VPWR VPWR _4717_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4648_ _4378_/A _5971_/A _4917_/A _5148_/C VGND VGND VPWR VPWR _4648_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5136__A2 _4708_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5166__A _5166_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4579_ _4878_/B VGND VGND VPWR VPWR _4581_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_1_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4220__D _4220_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4111__A3 _3674_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3414__A _4004_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5844__B1 _4420_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6147__D _6147_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5072__A1 _5069_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4890__D _5028_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4245__A _4245_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3083__A0 _6184_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3622__A2 _3621_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5375__A2 _5371_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4583__B1 _4581_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5780__C1 _5779_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3925__A3 _3342_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5076__A _5710_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4335__B1 _4364_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4886__A1 _4672_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3689__A2 _3680_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4099__C1 _3673_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5835__B1 _4882_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6153__CLK _6155_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3846__C1 _3845_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6057__D _6057_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5850__A3 _5148_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3861__A2 _3230_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5063__A1 _4350_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3950_ _3948_/Y _3868_/X _4146_/A _3949_/Y VGND VGND VPWR VPWR _3950_/X sky130_fd_sc_hd__a211o_1
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3881_ _3881_/A _3881_/B VGND VGND VPWR VPWR _3881_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6012__B1 _6207_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5620_ _5620_/A VGND VGND VPWR VPWR _6168_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__3916__A3 _3913_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3377__B2 _3374_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3377__A1 _3361_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5551_ _5551_/A VGND VGND VPWR VPWR _6141_/D sky130_fd_sc_hd__clkbuf_1
X_4502_ _4633_/S _4501_/X _4224_/A VGND VGND VPWR VPWR _4503_/A sky130_fd_sc_hd__a21oi_2
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5482_ _5482_/A VGND VGND VPWR VPWR _5482_/X sky130_fd_sc_hd__clkbuf_2
X_4433_ _4862_/A VGND VGND VPWR VPWR _4890_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4364_ _4364_/A VGND VGND VPWR VPWR _4364_/X sky130_fd_sc_hd__buf_2
XFILLER_113_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4295_ _4860_/A VGND VGND VPWR VPWR _5744_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_98_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3315_ _3315_/A _3606_/A VGND VGND VPWR VPWR _3956_/C sky130_fd_sc_hd__nor2_2
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6103_ _6145_/CLK _6103_/D VGND VGND VPWR VPWR _6103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5826__B1 _4565_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5152__C _5152_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3234__A _3582_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3246_ _3468_/A _3780_/C _3746_/A VGND VGND VPWR VPWR _3246_/X sky130_fd_sc_hd__or3b_2
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ _6202_/CLK _6034_/D VGND VGND VPWR VPWR _6034_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3177_ _3603_/D VGND VGND VPWR VPWR _3468_/A sky130_fd_sc_hd__buf_2
XFILLER_66_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3852__A2 _3722_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5841__A3 _4630_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4065__A _4065_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5054__A1 _4865_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3604__A2 _4004_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6003__B1 _5540_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5818_ _6144_/Q _5420_/A _5818_/S VGND VGND VPWR VPWR _5819_/A sky130_fd_sc_hd__mux2_2
XFILLER_10_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5762__C1 _5107_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3907__A3 _3711_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5749_ _4952_/B _5736_/Y _5673_/A _5748_/Y VGND VGND VPWR VPWR _5749_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_10_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6026__CLK _6045_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5109__A2 _4735_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3409__A _3648_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4231__C _4231_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4868__A1 _4857_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5624__A _5624_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6176__CLK _6176_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4885__D _5240_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4626__A1_N _4570_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3540__A1 _3508_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3144__A _3311_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5817__B1 _5811_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4096__A2 _4090_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2983__A input2/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3843__A2 _3320_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3056__A0 _6045_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4703__A _5003_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3319__A _3509_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4020__A2 _3829_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput109 _3124_/X VGND VGND VPWR VPWR memory_dmem_response_get[29] sky130_fd_sc_hd__buf_2
XFILLER_107_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5534__A _5534_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3531__A1 _3509_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3531__B2 _3517_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput91 _3087_/X VGND VGND VPWR VPWR memory_dmem_response_get[12] sky130_fd_sc_hd__buf_2
X_3100_ _3100_/A VGND VGND VPWR VPWR _3100_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5808__B1 _5804_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4087__A2 _4082_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4080_ _3300_/X _3919_/X _4076_/X _4079_/X _3828_/X VGND VGND VPWR VPWR _4080_/Y
+ sky130_fd_sc_hd__o221ai_2
XANTENNA__5823__A3 _5761_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3031_ _3031_/A VGND VGND VPWR VPWR _3031_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4492__C1 _4491_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5036__A1 _4998_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3598__A1 _3580_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4982_ _4975_/X _4980_/Y _4981_/Y _4189_/A VGND VGND VPWR VPWR _4982_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4795__B1 _4794_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3933_ _4083_/C _3932_/Y _3429_/X _3893_/X VGND VGND VPWR VPWR _3933_/X sky130_fd_sc_hd__o211a_1
XANTENNA__6049__CLK _6205_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3864_ _4083_/B _3864_/B VGND VGND VPWR VPWR _3975_/C sky130_fd_sc_hd__and2_4
XANTENNA__4547__B1 _4259_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5603_ _6161_/Q _6029_/Q _5605_/S VGND VGND VPWR VPWR _5604_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3229__A _4092_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3795_ _3580_/X _3794_/Y _3539_/X VGND VGND VPWR VPWR _3795_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4011__A2 _4010_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5534_ _5534_/A _6011_/B VGND VGND VPWR VPWR _6136_/D sky130_fd_sc_hd__nand2_1
XANTENNA__6199__CLK _6201_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3770__A1 _3760_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5465_ _5444_/X _5445_/X _5772_/C _5540_/A _5464_/X VGND VGND VPWR VPWR _6114_/D
+ sky130_fd_sc_hd__a311o_1
X_4416_ _4585_/A VGND VGND VPWR VPWR _5029_/A sky130_fd_sc_hd__buf_2
XANTENNA__5444__A _5444_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5511__A2 _4802_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5396_ _6178_/Q _2986_/B _4243_/X _4518_/A VGND VGND VPWR VPWR _5499_/A sky130_fd_sc_hd__o2bb2a_2
XFILLER_113_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4347_ _4347_/A VGND VGND VPWR VPWR _5976_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4278_ _4266_/A _4268_/Y _4277_/Y _4209_/A VGND VGND VPWR VPWR _4379_/A sky130_fd_sc_hd__o2bb2ai_4
XANTENNA__4078__A2 _4089_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3229_ _4092_/C VGND VGND VPWR VPWR _3882_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_74_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6017_ _6155_/CLK _6017_/D VGND VGND VPWR VPWR _6017_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3825__A2 _3824_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5027__B2 _5026_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5027__A1 _5971_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4250__A2 _4654_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4538__B1 _4882_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3139__A _3748_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6160__D _6160_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2978__A _5985_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5354__A _5354_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4710__B1 _4708_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4069__A2 _3254_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5266__A1 _6061_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5266__B2 _5265_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3959__D _3959_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output110_A _3065_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4433__A _4862_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3985__D1 _3242_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3975__C _3975_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5529__A _5529_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4152__B _4152_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6070__D _6070_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3049__A _3049_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5741__A2 _4929_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3580_ _3580_/A VGND VGND VPWR VPWR _3580_/X sky130_fd_sc_hd__buf_2
XANTENNA__3752__A1 _3744_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3752__B2 _3728_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5250_ _5096_/A _4414_/A _5078_/B _5152_/D _4461_/A VGND VGND VPWR VPWR _5250_/X
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__5264__A _5643_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3504__A1 _3363_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4201_ _4201_/A VGND VGND VPWR VPWR _4976_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5181_ _4777_/X _4778_/X _5687_/C _5687_/B _4686_/X VGND VGND VPWR VPWR _5181_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__3504__B2 _3502_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4132_ _3692_/A _4129_/Y _4130_/X _4131_/Y _3707_/A VGND VGND VPWR VPWR _4132_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__5711__B _5711_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4608__A _4832_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4063_ _3926_/X _4062_/Y _4036_/B VGND VGND VPWR VPWR _4063_/X sky130_fd_sc_hd__o21ba_1
XFILLER_3_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3512__A _3512_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3014_ _3014_/A VGND VGND VPWR VPWR _3014_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3231__B _3443_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4327__B _4527_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4768__B1 _4252_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4965_ _4865_/C _4480_/C _5000_/A _5005_/A VGND VGND VPWR VPWR _4965_/Y sky130_fd_sc_hd__o211ai_4
X_3916_ _3645_/A _4143_/A _3913_/X _3915_/X _3546_/A VGND VGND VPWR VPWR _3916_/X
+ sky130_fd_sc_hd__o311a_2
XANTENNA__4343__A _4555_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5439__A _5439_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4896_ _4926_/A VGND VGND VPWR VPWR _5096_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5980__A2 _5213_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3847_ _3847_/A _3847_/B _3847_/C VGND VGND VPWR VPWR _3847_/X sky130_fd_sc_hd__and3_2
XANTENNA__3991__A1 _3588_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5193__B1 _4869_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3778_ _3828_/A _3792_/C VGND VGND VPWR VPWR _3778_/X sky130_fd_sc_hd__or2_1
XANTENNA__4940__B1 _4618_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3743__B2 _3688_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5517_ _6130_/Q _5504_/X _5447_/X _5516_/Y VGND VGND VPWR VPWR _6130_/D sky130_fd_sc_hd__a211o_1
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4299__A2 _4244_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5448_ _6110_/Q _5222_/X _5256_/X _5260_/X VGND VGND VPWR VPWR _5448_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5496__B2 _5092_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5379_ _5376_/Y _5377_/Y _5378_/Y VGND VGND VPWR VPWR _6098_/D sky130_fd_sc_hd__a21oi_1
XFILLER_101_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5248__A1 _5118_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_86_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5799__A2 _4765_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4518__A _4518_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3422__A _3491_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6155__D _6155_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5956__C1 _4984_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4253__A _4282_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5349__A _5349_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4223__A2 _5044_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3431__B1 _3429_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5184__B1 _5680_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5723__A2 _5722_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3734__A1 _3238_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input71_A memory_dmem_request_put[97] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5239__A1 _5102_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5531__B _5531_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4428__A _4705_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3332__A _3663_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3670__B1 _3488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6065__D _6065_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3986__B _3986_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5947__C1 _5093_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5411__A1 _5406_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _4777_/A _4778_/A _4864_/B VGND VGND VPWR VPWR _4750_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__5962__A2 _5661_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4681_ _4680_/X _4551_/Y _5079_/A _4605_/X VGND VGND VPWR VPWR _4681_/Y sky130_fd_sc_hd__a31oi_4
X_3701_ _3701_/A VGND VGND VPWR VPWR _3701_/X sky130_fd_sc_hd__buf_2
XANTENNA__4193__A_N _5392_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3973__A1 _3961_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3973__B2 _3822_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3632_ _3632_/A VGND VGND VPWR VPWR _3633_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5714__A2 _4571_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4517__A3 input34/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4922__B1 _5148_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5706__B _5706_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3725__A1 _4126_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5190__A3 _4960_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3563_ _4036_/A VGND VGND VPWR VPWR _4126_/B sky130_fd_sc_hd__clkbuf_2
X_5302_ _6191_/Q _6067_/Q _5306_/S VGND VGND VPWR VPWR _5303_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3494_ _3592_/A _3462_/B _3468_/B _3588_/C VGND VGND VPWR VPWR _3494_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5478__A1 _5444_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5233_ _5076_/X _4971_/X _4459_/X _4954_/X VGND VGND VPWR VPWR _5233_/Y sky130_fd_sc_hd__o31ai_1
XANTENNA__4150__A1 _3668_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5164_ _5161_/X _5772_/B _5163_/X _4984_/X VGND VGND VPWR VPWR _5164_/X sky130_fd_sc_hd__a211o_1
X_4115_ _3680_/X _4073_/X _4111_/X _4114_/Y VGND VGND VPWR VPWR _4115_/X sky130_fd_sc_hd__a31o_1
XFILLER_29_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4338__A _4742_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3242__A _3707_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5095_ _5089_/X _4991_/X _5094_/X VGND VGND VPWR VPWR _5095_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_56_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4046_ _3962_/X _4041_/X _3838_/X _4045_/X VGND VGND VPWR VPWR _4046_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_37_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4989__B1 _4195_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4453__A2 _4551_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5650__A1 _6109_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3661__B1 _3429_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5047__A2_N _4991_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5938__C1 _5757_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5997_ _5998_/A _5998_/B _5998_/C _6201_/Q VGND VGND VPWR VPWR _5999_/A sky130_fd_sc_hd__a31o_1
XANTENNA__4073__A _4073_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4948_ _4948_/A VGND VGND VPWR VPWR _5973_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__5953__A2 _4957_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4504__C _4974_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4879_ _4879_/A VGND VGND VPWR VPWR _5755_/C sky130_fd_sc_hd__buf_2
XANTENNA__3964__A1 _3195_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4801__A _5968_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5705__A2 _5704_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3716__B2 _3674_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5181__A3 _5687_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3417__A _3781_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4913__B1 _4224_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4141__B2 _3891_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4141__A1 _4134_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3152__A _3275_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4248__A _4405_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5641__A1 _5445_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3652__B1 _3832_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5079__A _5079_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3955__A1 _3910_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5157__B1 _4767_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4904__B1 _4685_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3327__A _3571_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4132__A1 _3692_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4683__A2 _4677_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3465__A2_N _3674_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3062__A _5294_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5920_ _5918_/X _5919_/X _4665_/X VGND VGND VPWR VPWR _5920_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5632__A1 _6042_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5851_ _4360_/X _4960_/X _5880_/A _5025_/Y _4957_/A VGND VGND VPWR VPWR _5851_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5782_ _5782_/A VGND VGND VPWR VPWR _5782_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5935__A2 _4930_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4802_ _5203_/A VGND VGND VPWR VPWR _4802_/X sky130_fd_sc_hd__buf_2
XANTENNA__5396__B1 _4243_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2994_ _6016_/Q _6149_/Q _2998_/S VGND VGND VPWR VPWR _2995_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4733_ _4769_/B VGND VGND VPWR VPWR _4873_/A sky130_fd_sc_hd__buf_2
XANTENNA__3946__A1 _3428_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4621__A _4621_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4664_ _4645_/X _4664_/B _4664_/C VGND VGND VPWR VPWR _4664_/Y sky130_fd_sc_hd__nand3b_1
XANTENNA__5699__A1 _5691_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4595_ _4666_/A _4590_/X _4591_/Y _4594_/X VGND VGND VPWR VPWR _4595_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__3237__A _3983_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5708__A1_N _5145_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3615_ _3308_/A _3680_/A _3871_/B _3666_/A VGND VGND VPWR VPWR _3623_/B sky130_fd_sc_hd__and4b_1
X_3546_ _3546_/A VGND VGND VPWR VPWR _3546_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__4371__A1 _4307_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5216_ _5006_/X _4855_/A _5212_/X _4964_/A _5215_/Y VGND VGND VPWR VPWR _5216_/X
+ sky130_fd_sc_hd__o311a_1
X_3477_ _4102_/A VGND VGND VPWR VPWR _3477_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5320__A0 _6183_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5871__A1 _5862_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4123__B2 _3501_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6196_ _6196_/CLK _6196_/D VGND VGND VPWR VPWR _6196_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5871__B2 _4494_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5147_ _5061_/X _5062_/X _5102_/B _5032_/Y VGND VGND VPWR VPWR _5147_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5078_ _5078_/A _5078_/B _5687_/B _5078_/D VGND VGND VPWR VPWR _5078_/X sky130_fd_sc_hd__and4_1
XFILLER_56_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4029_ _4027_/X _4028_/Y _3476_/B VGND VGND VPWR VPWR _4029_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5084__C1 _5083_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4218__D _4218_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5623__A1 _6038_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4831__C1 _5880_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3700__A _3700_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3634__B1 _3633_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5926__A2 _5880_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3937__A1 _3910_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5139__B1 _4786_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3792__D _3792_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3147__A _3272_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4901__A3 _4856_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4114__A1 _3319_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5311__A0 _6195_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5362__A _5362_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5862__A1 _5179_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input34_A memory_dmem_request_put[60] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5614__A1 _6034_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4706__A _4772_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4822__C1 _4364_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3625__B1 _3624_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5090__A2 _4804_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2979__A2 _5998_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5917__A2 _5123_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3640__A3 _3453_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5378__B1 _5288_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3928__A1 _4124_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3389__C1 _3581_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4050__B1 _3520_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5537__A _5537_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6082__CLK _6202_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4441__A _4769_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3983__C _3983_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4380_ _4462_/A VGND VGND VPWR VPWR _4878_/B sky130_fd_sc_hd__buf_4
X_3400_ _4074_/A VGND VGND VPWR VPWR _3830_/D sky130_fd_sc_hd__buf_2
XFILLER_50_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3057__A _3057_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3331_ _3802_/B VGND VGND VPWR VPWR _3663_/A sky130_fd_sc_hd__clkbuf_4
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5302__A0 _6191_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3262_ _3657_/B VGND VGND VPWR VPWR _3468_/B sky130_fd_sc_hd__clkbuf_2
X_6050_ _6196_/CLK _6050_/D VGND VGND VPWR VPWR _6050_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5853__A1 _5745_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5001_ _5944_/A _5971_/C _5944_/D _4742_/X VGND VGND VPWR VPWR _5001_/X sky130_fd_sc_hd__a31o_1
X_3193_ _3780_/C VGND VGND VPWR VPWR _4089_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5605__A1 _6030_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4616__A _4937_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5081__A2 _4464_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3520__A _3732_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3616__B1 _3756_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5903_ _5903_/A _5903_/B _5903_/C _5903_/D VGND VGND VPWR VPWR _5903_/X sky130_fd_sc_hd__and4_1
XANTENNA__3092__A1 _6080_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5834_ _5899_/A _5745_/B _5710_/A _4827_/A _4440_/Y VGND VGND VPWR VPWR _5834_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__5369__B1 _5367_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5908__A2 _5955_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4041__B1 _4040_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5765_ _5735_/X _5764_/Y _5175_/A VGND VGND VPWR VPWR _5765_/Y sky130_fd_sc_hd__o21ai_1
X_2977_ _6199_/Q VGND VGND VPWR VPWR _5985_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5447__A _5545_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4351__A _4566_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5696_ _4422_/A _4699_/X _5148_/B _5695_/X _5148_/A VGND VGND VPWR VPWR _5696_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__3893__C _3893_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3395__A2 _3393_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4716_ _4716_/A VGND VGND VPWR VPWR _4716_/X sky130_fd_sc_hd__buf_2
X_4647_ _5022_/A VGND VGND VPWR VPWR _5148_/C sky130_fd_sc_hd__buf_2
XANTENNA__5136__A3 _5148_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5166__B _5166_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4578_ _4578_/A VGND VGND VPWR VPWR _5711_/B sky130_fd_sc_hd__buf_2
XFILLER_115_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5182__A _5182_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3529_ _3403_/X _3524_/X _3525_/X _3749_/D _3537_/A VGND VGND VPWR VPWR _3529_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__3414__B _3527_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5844__A1 _5235_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6179_ _6205_/CLK _6179_/D VGND VGND VPWR VPWR _6179_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3855__B1 _3142_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4526__A _5188_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3430__A _3746_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5072__A2 _5071_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3083__A1 _6076_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6163__D _6163_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4032__B1 _6039_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4583__A1 _4574_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4261__A _6133_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5780__B1 _5145_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3925__A4 _3653_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4335__A1 _4307_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4886__A2 _4332_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5092__A _5529_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4099__B1 _3418_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5835__A1 _5867_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output140_A _2997_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3846__B1 _3843_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4436__A _4696_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3340__A _3546_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5599__A0 _6159_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5063__A2 _4725_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6073__D _6073_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3880_ _3863_/X _3865_/Y _3624_/X _3866_/X _3879_/X VGND VGND VPWR VPWR _3880_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_16_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6012__A1 _6202_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4023__B1 _4022_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5267__A input4/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3377__A2 _3363_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5550_ _5550_/A _5568_/B VGND VGND VPWR VPWR _5551_/A sky130_fd_sc_hd__and2_1
XANTENNA__4171__A _4171_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5771__B1 _5766_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4501_ _4501_/A VGND VGND VPWR VPWR _4501_/X sky130_fd_sc_hd__buf_4
X_5481_ _5481_/A VGND VGND VPWR VPWR _6119_/D sky130_fd_sc_hd__clkbuf_1
X_4432_ _4432_/A VGND VGND VPWR VPWR _4862_/A sky130_fd_sc_hd__buf_2
XFILLER_6_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3515__A _4004_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4363_ _4363_/A VGND VGND VPWR VPWR _5263_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4294_ _4313_/A _4293_/Y _4234_/A _6133_/Q VGND VGND VPWR VPWR _4860_/A sky130_fd_sc_hd__a22oi_4
X_3314_ _3867_/A _4135_/B _3767_/B VGND VGND VPWR VPWR _3314_/Y sky130_fd_sc_hd__o21ai_4
X_6102_ _6146_/CLK _6102_/D VGND VGND VPWR VPWR _6102_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5826__A1 _4843_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3245_ _3781_/B VGND VGND VPWR VPWR _3746_/A sky130_fd_sc_hd__clkbuf_2
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ _6202_/CLK _6033_/D VGND VGND VPWR VPWR _6033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5152__D _5152_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3837__B1 _4124_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ _3870_/A VGND VGND VPWR VPWR _3780_/C sky130_fd_sc_hd__buf_2
XANTENNA__3250__A _3440_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3852__A3 _3731_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5054__A2 _4865_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4065__B _4065_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4262__B1 _4261_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3604__A3 _3686_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6003__A1 _3060_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4014__B1 _3350_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5817_ _6188_/Q _4715_/X _5811_/Y _5816_/Y VGND VGND VPWR VPWR _6188_/D sky130_fd_sc_hd__a2bb2oi_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5762__B1 _4364_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5748_ _4570_/Y _4571_/X _5740_/Y _5747_/X VGND VGND VPWR VPWR _5748_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5905__A _5905_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4231__D _4231_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5679_ _5676_/X _5678_/X _5811_/A VGND VGND VPWR VPWR _5679_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__4868__A2 _4867_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3425__A _3525_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3540__A2 _3531_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5817__B2 _5816_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6158__D _6158_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4096__A3 _4091_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3160__A _3673_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3056__A1 _6177_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_9_0_CLK clkbuf_4_9_0_CLK/A VGND VGND VPWR VPWR _6207_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4005__B1 _3476_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5753__B1 _4345_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5087__A _5757_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4020__A3 _3720_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6120__CLK _6145_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5505__B1 _5504_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5534__B _6011_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3335__A _4083_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3531__A2 _3510_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput92 _3089_/X VGND VGND VPWR VPWR memory_dmem_response_get[13] sky130_fd_sc_hd__buf_2
XANTENNA__5808__A1 _5791_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5808__B2 _5807_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6068__D _6068_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4087__A3 _4086_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5550__A _5550_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3819__B1 _3492_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4492__B1 _4665_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3030_ _6033_/Q _6165_/Q _3032_/S VGND VGND VPWR VPWR _3031_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4166__A _4301_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5036__A2 _5027_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4981_ _6132_/Q _4807_/X _4224_/X VGND VGND VPWR VPWR _4981_/Y sky130_fd_sc_hd__o21ai_1
X_3932_ _3967_/A _3932_/B VGND VGND VPWR VPWR _3932_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4795__A1 _4668_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3452__D1 _3744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3598__A2 _3597_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3863_ _3161_/X _3857_/Y _3861_/Y _4039_/B VGND VGND VPWR VPWR _3863_/X sky130_fd_sc_hd__a211o_1
XFILLER_32_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4547__A1 _4878_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5602_ _5602_/A VGND VGND VPWR VPWR _6160_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5533_ _4801_/X _4482_/B _5092_/X _5504_/A _4254_/Y VGND VGND VPWR VPWR _5534_/A
+ sky130_fd_sc_hd__a32o_1
X_3794_ _3699_/X _3793_/X _3766_/Y VGND VGND VPWR VPWR _3794_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__4011__A3 _3821_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5725__A _5725_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3770__A2 _3457_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5464_ _6114_/Q _5222_/X _5256_/X _5260_/X VGND VGND VPWR VPWR _5464_/X sky130_fd_sc_hd__o22a_1
X_4415_ _4415_/A VGND VGND VPWR VPWR _4585_/A sky130_fd_sc_hd__buf_2
X_5395_ _5395_/A VGND VGND VPWR VPWR _5395_/X sky130_fd_sc_hd__clkbuf_2
X_4346_ _4306_/Y _4316_/X _4339_/X _4345_/X VGND VGND VPWR VPWR _4346_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3245__A _3781_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5511__A3 _5262_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4277_ _6134_/Q VGND VGND VPWR VPWR _4277_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5460__A _5460_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3228_ _3621_/A _3500_/A VGND VGND VPWR VPWR _4092_/C sky130_fd_sc_hd__nand2_2
XFILLER_86_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6016_ _6197_/CLK _6016_/D VGND VGND VPWR VPWR _6016_/Q sky130_fd_sc_hd__dfxtp_1
X_3159_ _3647_/A VGND VGND VPWR VPWR _3673_/A sky130_fd_sc_hd__buf_4
XFILLER_36_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5027__A2 _5025_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5983__B1 _4190_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4804__A _4804_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4250__A3 _4910_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4538__A1 _4937_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5735__B1 _4950_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6143__CLK _6205_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5635__A _5635_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_108_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3155__A _3162_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4710__A1 _4422_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4069__A3 _3830_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5266__A2 _5166_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4474__B1 _4742_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5974__B1 _5929_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output103_A _3111_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3985__C1 _3984_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3975__D _3975_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3737__C1 _3911_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4152__C _4152_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5726__B1 _5703_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5545__A _5545_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3752__A2 _3751_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5264__B _5643_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3504__A2 _3496_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4162__C1 _3580_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3065__A _3065_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4200_ input6/X _4200_/B VGND VGND VPWR VPWR _4201_/A sky130_fd_sc_hd__and2b_1
X_5180_ _4871_/Y _5706_/C _5179_/X _4998_/X VGND VGND VPWR VPWR _5180_/Y sky130_fd_sc_hd__a31oi_4
XFILLER_122_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4131_ _4061_/X _3904_/X _3663_/C VGND VGND VPWR VPWR _4131_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5711__C _5745_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4062_ _3967_/X _3524_/X _4061_/X VGND VGND VPWR VPWR _4062_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5662__C1 _5661_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4465__B1 _4341_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3013_ _6025_/Q _6157_/Q _3021_/S VGND VGND VPWR VPWR _3014_/A sky130_fd_sc_hd__mux2_1
XANTENNA__6016__CLK _6197_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4327__C _4358_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3004__S _3010_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4768__B2 _4766_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4768__A1 _4732_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4624__A _4819_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4964_ _4964_/A VGND VGND VPWR VPWR _4964_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5965__B1 _5734_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3915_ _3799_/A _3583_/C _3594_/A _3914_/Y VGND VGND VPWR VPWR _3915_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3976__C1 _3838_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6166__CLK _6203_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4895_ _4895_/A VGND VGND VPWR VPWR _5240_/D sky130_fd_sc_hd__buf_4
XANTENNA__5980__A3 _5959_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5717__B1 _5106_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3991__A2 _3593_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3846_ _4126_/B _3733_/Y _3843_/Y _3845_/X VGND VGND VPWR VPWR _3846_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5193__A1 _5118_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3777_ _3775_/Y _3776_/Y _3562_/X VGND VGND VPWR VPWR _3777_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4940__A1 _4680_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5516_ _4806_/Y _5433_/X _5504_/A VGND VGND VPWR VPWR _5516_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5447_ _5545_/A VGND VGND VPWR VPWR _5447_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_105_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4299__A3 _4308_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5378_ _5376_/Y _5377_/Y _5288_/X VGND VGND VPWR VPWR _5378_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4329_ _4601_/A VGND VGND VPWR VPWR _4329_/X sky130_fd_sc_hd__buf_2
XANTENNA__5248__A2 _5003_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3703__A _3703_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5799__A3 _5973_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5200__A2_N _5040_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5956__B1 _5163_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4223__A3 _5648_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3431__A1 _3428_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6171__D _6171_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5708__B1 _5707_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5184__A1 _5048_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2989__A _5294_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3734__A2 _3733_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input64_A memory_dmem_request_put[90] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4144__C1 _3537_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5892__C1 _4875_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6039__CLK _6074_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5239__A2 _5008_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3613__A _3613_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5304__S _5306_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6189__CLK _6205_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3670__A1 _3659_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3982__A_N _4088_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4444__A _4549_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5947__B1 _5163_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3986__C _4088_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5411__A2 _5409_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ _3700_/A VGND VGND VPWR VPWR _3701_/A sky130_fd_sc_hd__buf_4
XANTENNA__6081__D _6081_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4680_ _4680_/A VGND VGND VPWR VPWR _4680_/X sky130_fd_sc_hd__buf_2
XANTENNA__3973__A2 _3972_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3631_ _3631_/A VGND VGND VPWR VPWR _3631_/X sky130_fd_sc_hd__buf_2
XANTENNA__4922__A1 _5976_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5706__C _5706_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3562_ _3562_/A VGND VGND VPWR VPWR _3562_/X sky130_fd_sc_hd__buf_2
XANTENNA__3725__A2 _3718_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5275__A _5275_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4922__B2 _4708_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5301_ _5301_/A VGND VGND VPWR VPWR _6066_/D sky130_fd_sc_hd__clkbuf_1
X_3493_ _3606_/A VGND VGND VPWR VPWR _3592_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5478__A2 _5046_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5232_ _5230_/X _5231_/X _4765_/X VGND VGND VPWR VPWR _5232_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5883__C1 _5878_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4619__A _5188_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4150__A2 _3549_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5163_ _5163_/A VGND VGND VPWR VPWR _5163_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3523__A _3588_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4114_ _3319_/X _4112_/X _4113_/X VGND VGND VPWR VPWR _4114_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5094_ _5090_/X _5444_/A _5092_/X _5093_/X VGND VGND VPWR VPWR _5094_/X sky130_fd_sc_hd__a211o_1
XFILLER_83_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4045_ _3764_/X _4042_/X _4043_/X _3975_/C _4044_/Y VGND VGND VPWR VPWR _4045_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_56_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3110__A0 _6059_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4989__A1 _5392_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3661__A1 _3659_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5650__A2 _4511_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4354__A _4354_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5938__B1 _5756_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3949__C1 _3369_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5996_ _5570_/X _5994_/Y _5995_/X _5388_/A VGND VGND VPWR VPWR _6200_/D sky130_fd_sc_hd__a211o_1
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4947_ _4552_/X _4945_/X _5018_/C _4538_/X VGND VGND VPWR VPWR _4947_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4073__B _4073_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4071__D1 _4070_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4878_ _4878_/A _4878_/B _4878_/C _4878_/D VGND VGND VPWR VPWR _4878_/Y sky130_fd_sc_hd__nand4_4
XANTENNA__3964__A2 _3194_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3829_ _4074_/B VGND VGND VPWR VPWR _3829_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4913__A1 _6131_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4529__A _4578_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4677__B1 _4676_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4141__A2 _4140_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3433__A _3904_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4994__C_N _4200_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6166__D _6166_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3101__A0 _6056_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3652__A1 _3512_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5641__A2 _5640_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4264__A _4268_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5079__B _5079_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5929__B1 _5928_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3955__A2 _3975_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5157__A1 _5150_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4904__A1 _4881_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4132__A2 _4129_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4439__A _4926_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3343__A _3343_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6076__D _6076_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4174__A _4174_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5850_ _4726_/A _5706_/C _5148_/C _4541_/A VGND VGND VPWR VPWR _5850_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5935__A3 _5080_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5781_ _4924_/X _5063_/X _5064_/X _5780_/Y _4794_/X VGND VGND VPWR VPWR _5781_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__5396__B2 _4518_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2993_ _2993_/A VGND VGND VPWR VPWR _2993_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4801_ _5968_/C VGND VGND VPWR VPWR _4801_/X sky130_fd_sc_hd__clkbuf_4
X_4732_ _4732_/A _4732_/B _4732_/C VGND VGND VPWR VPWR _4732_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__3946__A2 _3895_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4663_ _5757_/B _5263_/A _4657_/X _4662_/X _5756_/A VGND VGND VPWR VPWR _4664_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_119_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3518__A _4034_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3614_ _3614_/A VGND VGND VPWR VPWR _3666_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5699__A2 _5698_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6204__CLK _6204_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4594_ _4668_/A _5000_/A _5029_/A _5021_/A _4744_/A VGND VGND VPWR VPWR _4594_/X
+ sky130_fd_sc_hd__o41a_1
X_3545_ _3773_/A _4092_/C _3967_/A _3700_/A VGND VGND VPWR VPWR _4036_/B sky130_fd_sc_hd__and4_1
XANTENNA__4371__A2 _4362_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3476_ _3476_/A _3476_/B _3476_/C _3476_/D VGND VGND VPWR VPWR _3476_/X sky130_fd_sc_hd__or4_4
XANTENNA__5733__A _5955_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5215_ _5836_/A _5213_/X _5214_/X VGND VGND VPWR VPWR _5215_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5320__A1 _6075_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4349__A _4769_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3253__A _3858_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6195_ _6196_/CLK _6195_/D VGND VGND VPWR VPWR _6195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5871__A2 _5865_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5146_ _5680_/A _4739_/X _4668_/X _4726_/A _5145_/X VGND VGND VPWR VPWR _5150_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5077_ _4945_/X _5076_/X _4823_/X _4824_/X _4943_/Y VGND VGND VPWR VPWR _5077_/Y
+ sky130_fd_sc_hd__a2111oi_2
XFILLER_84_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4028_ _3679_/X _4042_/C _3444_/X _3902_/A _4048_/A VGND VGND VPWR VPWR _4028_/Y
+ sky130_fd_sc_hd__a221oi_1
XANTENNA__5084__B1 _4393_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4831__B1 _4829_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3634__A1 _3343_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5979_ _5061_/X _5062_/X _5063_/X _4898_/Y VGND VGND VPWR VPWR _5979_/Y sky130_fd_sc_hd__o22ai_2
XFILLER_52_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4595__C1 _4594_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3937__A2 _3626_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5792__D1 _5752_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5139__A1 _4859_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3428__A _3902_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_119_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4898__B1 _4897_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3570__B1 _3600_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5643__A _5643_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4114__A2 _4112_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5311__A1 _6071_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5847__C1 _5846_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2986__B _2986_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4259__A _4259_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3163__A _3513_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5862__A2 _5859_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_85_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input27_A memory_dmem_request_put[53] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5075__B1 _4875_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_85_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4822__B1 _4937_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3625__A1 _3613_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_71_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5378__A1 _5376_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5917__A3 _5179_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3928__A2 _3895_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3389__B1 _3657_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5783__D1 _5752_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4050__A1 _3626_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5537__B _5568_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4441__B _4769_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3338__A _3835_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4889__B1 _4420_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output95_A _3095_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3330_ _3330_/A VGND VGND VPWR VPWR _3802_/B sky130_fd_sc_hd__buf_2
XANTENNA__5553__A _5988_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5838__C1 _5837_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3261_ _3461_/B _3311_/B VGND VGND VPWR VPWR _3657_/B sky130_fd_sc_hd__or2b_2
X_5000_ _5000_/A VGND VGND VPWR VPWR _5944_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__3073__A _3073_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4169__A _4169_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5302__A1 _6067_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5853__A2 _5899_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3192_ _3343_/A VGND VGND VPWR VPWR _3195_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5066__B1 _5060_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4813__B1 _4924_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3616__A1 _3406_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5902_ _4858_/Y _4859_/X _5901_/Y VGND VGND VPWR VPWR _5902_/Y sky130_fd_sc_hd__o21ai_1
X_5833_ _4332_/X _5018_/A _5148_/D _5761_/A _4328_/X VGND VGND VPWR VPWR _5833_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_62_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5369__A1 _4520_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5764_ _5722_/Y _5763_/X _5228_/X VGND VGND VPWR VPWR _5764_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4041__A1 _3679_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2976_ _6100_/Q VGND VGND VPWR VPWR _5998_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3248__A _3315_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5695_ _4404_/X _4405_/X _4296_/X _4668_/A VGND VGND VPWR VPWR _5695_/X sky130_fd_sc_hd__o22a_1
X_4715_ _5646_/A VGND VGND VPWR VPWR _4715_/X sky130_fd_sc_hd__clkbuf_2
X_4646_ _4854_/A VGND VGND VPWR VPWR _4917_/A sky130_fd_sc_hd__clkbuf_4
X_4577_ _5067_/A VGND VGND VPWR VPWR _5034_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__5136__A4 _5148_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3552__B1 _3600_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5463__A _5545_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3528_ _3528_/A VGND VGND VPWR VPWR _3537_/A sky130_fd_sc_hd__buf_2
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3459_ _3983_/C VGND VGND VPWR VPWR _4042_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_97_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3414__C _3708_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5844__A2 _4927_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3855__A1 _3846_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6178_ _6207_/CLK _6178_/D VGND VGND VPWR VPWR _6178_/Q sky130_fd_sc_hd__dfxtp_1
X_5129_ _4984_/X _5757_/C _5757_/D _6120_/Q _4987_/X VGND VGND VPWR VPWR _5129_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3711__A _3711_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5057__B1 _4252_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4807__A _4807_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4032__B2 _3891_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4032__A1 _4031_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4583__A2 _4576_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3158__A _3609_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5780__A1 _5880_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3791__B1 _3707_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4335__A2 _4362_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2997__A _2997_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4099__A1 _3668_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5835__A2 _4945_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3846__A1 _4126_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3621__A _3621_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4717__A _4717_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output133_A _3040_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5599__A1 _6027_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5548__A _5548_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6012__A2 _6205_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4452__A _4533_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4023__A1 _3536_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4171__B _4171_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5771__A1 _5751_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5771__B2 _5770_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3782__B1 _3528_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4500_ _6142_/Q _6141_/Q VGND VGND VPWR VPWR _4501_/A sky130_fd_sc_hd__or2_1
X_5480_ _5480_/A _5501_/B VGND VGND VPWR VPWR _5481_/A sky130_fd_sc_hd__and2_1
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4431_ _5706_/A VGND VGND VPWR VPWR _4431_/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__5283__A _5285_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4731__C1 _4730_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4362_ _4362_/A VGND VGND VPWR VPWR _4362_/X sky130_fd_sc_hd__buf_2
XFILLER_112_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4293_ _4293_/A _4293_/B VGND VGND VPWR VPWR _4293_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3515__B _3515_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3313_ _3382_/D VGND VGND VPWR VPWR _3767_/B sky130_fd_sc_hd__clkbuf_4
X_6101_ _6145_/CLK _6101_/D VGND VGND VPWR VPWR _6101_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5826__A2 _5899_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3244_ _3315_/A VGND VGND VPWR VPWR _3781_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_86_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ _6202_/CLK _6032_/D VGND VGND VPWR VPWR _6032_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3837__B2 _3836_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3837__A1 _3830_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3175_ _3440_/B VGND VGND VPWR VPWR _3870_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5039__B1 _4995_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3250__B _3366_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4262__A1 _4301_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4065__C _4092_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6003__A2 _5291_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4014__A1 _3343_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4362__A _4362_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5816_ _4952_/B _5814_/Y _5815_/Y _5725_/C VGND VGND VPWR VPWR _5816_/Y sky130_fd_sc_hd__o211ai_2
XFILLER_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5762__A1 _4362_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5747_ _5709_/Y _5708_/Y _5746_/Y _5237_/A VGND VGND VPWR VPWR _5747_/X sky130_fd_sc_hd__o211a_1
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4970__C1 _4969_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5678_ _6110_/Q _4721_/X _5677_/X VGND VGND VPWR VPWR _5678_/X sky130_fd_sc_hd__a21o_1
X_4629_ _4629_/A VGND VGND VPWR VPWR _4629_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3425__B _3631_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6072__CLK _6074_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5640__B _6098_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4537__A _4585_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3441__A _3873_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6174__D _6174_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5450__B1 _5439_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4005__A1 _3299_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4272__A _4301_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5202__B1 _5042_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5753__A1 _4328_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4961__C1 _4960_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3516__B1 _3748_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5505__A1 _4522_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3335__B _4074_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput93 _3091_/X VGND VGND VPWR VPWR memory_dmem_response_get[14] sky130_fd_sc_hd__buf_2
XANTENNA__5808__A2 _5166_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5550__B _5568_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3819__A1 _3818_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4447__A _4869_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4492__A1 _4474_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5036__A3 _5030_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6084__D _6084_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4980_ _4716_/X _4513_/X input40/X _4977_/X _4979_/X VGND VGND VPWR VPWR _4980_/Y
+ sky130_fd_sc_hd__o311ai_4
XANTENNA__5441__B1 _5398_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4795__A2 _5829_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3931_ _3867_/X _3881_/B _3195_/A _3308_/X VGND VGND VPWR VPWR _3931_/Y sky130_fd_sc_hd__a31oi_1
XANTENNA__3452__C1 _3450_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5278__A _6063_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5992__A1 _6200_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3862_ _3862_/A VGND VGND VPWR VPWR _4039_/B sky130_fd_sc_hd__buf_2
XFILLER_32_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4182__A _4231_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4547__A2 _4754_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5601_ _6160_/Q _6028_/Q _5605_/S VGND VGND VPWR VPWR _5602_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4910__A _4910_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5532_ _5532_/A VGND VGND VPWR VPWR _6135_/D sky130_fd_sc_hd__clkbuf_1
X_3793_ _3673_/Y _3293_/X _3767_/X _3674_/X VGND VGND VPWR VPWR _3793_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5725__B _5725_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3526__A _3526_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3770__A3 _3762_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5463_ _5545_/A VGND VGND VPWR VPWR _5540_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4414_ _4414_/A VGND VGND VPWR VPWR _5976_/A sky130_fd_sc_hd__clkbuf_4
X_5394_ _5420_/A VGND VGND VPWR VPWR _5395_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4345_ _4345_/A VGND VGND VPWR VPWR _4345_/X sky130_fd_sc_hd__buf_4
XANTENNA__6095__CLK _6204_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4276_ _4769_/C VGND VGND VPWR VPWR _5211_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5460__B _5468_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3261__A _3461_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3227_ _3437_/A _3606_/A VGND VGND VPWR VPWR _3500_/A sky130_fd_sc_hd__nand2_2
XFILLER_86_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4357__A _4738_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6015_ _6015_/A VGND VGND VPWR VPWR _6207_/D sky130_fd_sc_hd__clkbuf_1
X_3158_ _3609_/B VGND VGND VPWR VPWR _3647_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3089_ _3089_/A VGND VGND VPWR VPWR _3089_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5188__A _5188_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5983__B2 _6196_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4092__A _4092_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3994__B1 _3711_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4538__A2 _4536_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5196__C1 _5195_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5735__A1 _5712_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3436__A _3802_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2986__A_N _5640_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6169__D _6169_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4710__A2 _4699_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5651__A _5811_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5120__C1 _5152_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4474__A1 _4852_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4267__A _4405_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3171__A _3353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5671__B1 _4498_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5098__A _5098_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5974__A1 _5756_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5974__B2 _5973_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3985__B1 _3623_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3110__S _3116_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5187__C1 _4675_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3737__B1 _3756_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5726__B2 _5725_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3752__A3 _3727_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3346__A _3711_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5264__C _6128_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4162__B1 _4161_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6079__D _6079_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4130_ _3583_/C _3515_/B _3551_/A _3700_/A VGND VGND VPWR VPWR _4130_/X sky130_fd_sc_hd__a31o_1
XFILLER_122_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5111__C1 _4572_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4061_ _4061_/A VGND VGND VPWR VPWR _4061_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4465__A1 _4340_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4177__A _4230_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5662__B1 _5031_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3012_ _3056_/S VGND VGND VPWR VPWR _3021_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__4327__D _4878_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4768__A2 _4746_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4963_ _4487_/Y _4959_/X _4891_/X _4961_/Y _4962_/X VGND VGND VPWR VPWR _4963_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__5965__A1 _5746_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3914_ _3780_/A _4092_/B _3382_/D _4073_/B VGND VGND VPWR VPWR _3914_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_51_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3976__B1 _3975_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4894_ _4843_/A _4565_/A _4887_/X _5034_/C _4551_/Y VGND VGND VPWR VPWR _4894_/X
+ sky130_fd_sc_hd__o2111a_4
XANTENNA__5717__A1 _4686_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5178__C1 _5188_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5717__B2 _4820_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3991__A3 _3703_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3845_ _3844_/X _3687_/Y _3534_/X _3293_/X _3301_/A VGND VGND VPWR VPWR _3845_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_20_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4640__A _4640_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5193__A2 _5711_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3776_ _3673_/Y _3674_/X _3479_/X VGND VGND VPWR VPWR _3776_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4940__A2 _4935_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5515_ _5515_/A VGND VGND VPWR VPWR _6129_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3256__A _3386_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5446_ input18/X _5437_/X _5439_/X input10/X VGND VGND VPWR VPWR _5677_/C sky130_fd_sc_hd__a22o_1
Xclkbuf_4_8_0_CLK clkbuf_4_9_0_CLK/A VGND VGND VPWR VPWR _6204_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_121_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4153__B1 _3643_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4299__A4 _4245_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5377_ _6097_/Q _5368_/X _5371_/A VGND VGND VPWR VPWR _5377_/Y sky130_fd_sc_hd__o21ai_1
X_4328_ _5667_/A VGND VGND VPWR VPWR _4328_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_86_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3900__B1 _3643_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5248__A3 _5003_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4259_ _4259_/A VGND VGND VPWR VPWR _4890_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input1_A EN_memory_dmem_request_put VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_101_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5653__B1 _5107_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3664__C1 _3663_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4815__A _4862_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6110__CLK _6204_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5956__A1 input15/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3431__A2 _3410_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5708__B2 _4924_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5646__A _5646_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4550__A _4769_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5184__A2 _5021_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4916__C1 _5034_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3166__A _3461_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4144__B1 _3369_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input57_A memory_dmem_request_put[83] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5381__A _6099_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5892__B1 _5891_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5239__A3 _5009_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3613__B _3613_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3105__S _3105_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5644__B1 _5643_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4725__A _4725_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3670__A2 _3673_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5320__S _5328_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4444__B _4884_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5947__A1 input14/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3986__D _4088_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3958__B1 _3992_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4080__C1 _3828_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3973__A3 _3821_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3630_ _3663_/C VGND VGND VPWR VPWR _4124_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__4907__C1 _4978_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4922__A2 _5971_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3561_ _3707_/A VGND VGND VPWR VPWR _3562_/A sky130_fd_sc_hd__buf_4
XANTENNA__3725__A3 _3721_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5275__B _5275_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3076__A _3076_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5300_ _6190_/Q _6066_/Q _5306_/S VGND VGND VPWR VPWR _5301_/A sky130_fd_sc_hd__mux2_1
X_3492_ _3959_/D VGND VGND VPWR VPWR _3492_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5231_ _5018_/C _5021_/A _5028_/X _5080_/X _4675_/X VGND VGND VPWR VPWR _5231_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_69_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5478__A3 _5445_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5883__B1 _4783_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4150__A3 _3831_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5162_ _5162_/A VGND VGND VPWR VPWR _5163_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4619__B _4619_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4113_ _3527_/C _3703_/A _4074_/C _3589_/B _3607_/X VGND VGND VPWR VPWR _4113_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__3894__C1 _3893_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5093_ _5093_/A VGND VGND VPWR VPWR _5093_/X sky130_fd_sc_hd__buf_2
XANTENNA__6133__CLK _6146_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3015__S _3021_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4044_ _4044_/A _4044_/B _4044_/C _3990_/X VGND VGND VPWR VPWR _4044_/Y sky130_fd_sc_hd__nor4b_1
XANTENNA__3646__C1 _3546_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3110__A1 _6088_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4989__A2 _5438_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3661__A2 _3660_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4354__B _4354_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5938__A1 _4657_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3949__B1 _3701_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5995_ _5984_/Y _5985_/Y _6200_/Q VGND VGND VPWR VPWR _5995_/X sky130_fd_sc_hd__o21a_1
XFILLER_24_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4946_ _4946_/A VGND VGND VPWR VPWR _5018_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__4073__C _4073_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4071__C1 _4069_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4877_ _5152_/C VGND VGND VPWR VPWR _5944_/C sky130_fd_sc_hd__buf_2
XANTENNA__3964__A3 _3767_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3828_ _3828_/A VGND VGND VPWR VPWR _3828_/X sky130_fd_sc_hd__buf_2
XANTENNA__5571__C1 _6197_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4913__A2 _4975_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3759_ _4002_/A _3759_/B _3816_/D VGND VGND VPWR VPWR _3759_/X sky130_fd_sc_hd__or3_1
XFILLER_121_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4677__A1 _5004_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5429_ _5429_/A _5468_/B VGND VGND VPWR VPWR _5430_/A sky130_fd_sc_hd__and2_1
XFILLER_114_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4141__A3 _3290_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4529__B _4734_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_114_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3637__C1 _3749_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3101__A1 _6084_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4545__A _5073_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4044__D_N _3990_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3652__A2 _4135_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5929__A1 _5235_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4264__B _4293_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5929__B2 _5145_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6182__D _6182_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5079__C _5079_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3955__A3 _3359_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4280__A _4860_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5157__A2 _5156_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5376__A _6098_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4904__A2 _4889_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4117__B1 _4102_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5865__B1 _5734_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4132__A3 _4130_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5315__S _5317_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3624__A _3806_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6000__A _6000_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6156__CLK _6197_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4800_ _4800_/A VGND VGND VPWR VPWR _5968_/C sky130_fd_sc_hd__buf_2
XANTENNA__6092__D _6092_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4174__B _4174_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5250__D1 _4461_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5780_ _5880_/A _5025_/Y _5145_/X _5779_/X VGND VGND VPWR VPWR _5780_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_61_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2992_ _6017_/Q _6148_/Q _2998_/S VGND VGND VPWR VPWR _2993_/A sky130_fd_sc_hd__mux2_1
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _4692_/X _4353_/X _4524_/X _4666_/A _4730_/Y VGND VGND VPWR VPWR _4732_/C
+ sky130_fd_sc_hd__o311a_1
XANTENNA__3946__A3 _3720_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4662_ _5167_/A _4672_/A _5680_/B _4661_/X VGND VGND VPWR VPWR _4662_/X sky130_fd_sc_hd__o211a_1
XANTENNA__4190__A _5646_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5286__A _6064_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5002__D1 _5001_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3613_ _3613_/A _3613_/B _3612_/X _3562_/A VGND VGND VPWR VPWR _3613_/X sky130_fd_sc_hd__or4bb_1
X_4593_ _5008_/A _5009_/A _4929_/A VGND VGND VPWR VPWR _5021_/A sky130_fd_sc_hd__a21oi_4
X_3544_ _3780_/A VGND VGND VPWR VPWR _3967_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4371__A3 _4308_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3475_ _3911_/A _3674_/C _3871_/A _3475_/D VGND VGND VPWR VPWR _3476_/D sky130_fd_sc_hd__and4b_1
XANTENNA__4108__B1 _3242_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5733__B _5733_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5856__B1 _4732_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5214_ _5211_/X _4754_/X _4750_/Y _4642_/A _5743_/B VGND VGND VPWR VPWR _5214_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_69_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3534__A _3756_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6194_ _6196_/CLK _6194_/D VGND VGND VPWR VPWR _6194_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5145_ _5145_/A VGND VGND VPWR VPWR _5145_/X sky130_fd_sc_hd__buf_4
XFILLER_57_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5608__A0 _6163_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5076_ _5710_/A VGND VGND VPWR VPWR _5076_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5084__A1 _5066_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3619__C1 _3281_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4365__A _4769_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4027_ _3549_/A _3871_/B _3482_/A _3574_/A _3659_/X VGND VGND VPWR VPWR _4027_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_84_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4831__A1 _5745_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3634__A2 _3631_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5978_ _5976_/X _4556_/X _5228_/X _5977_/X VGND VGND VPWR VPWR _5978_/Y sky130_fd_sc_hd__o211ai_2
X_4929_ _4929_/A _4929_/B _4929_/C VGND VGND VPWR VPWR _5098_/A sky130_fd_sc_hd__nor3_4
XANTENNA__4595__B1 _4591_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3937__A3 _3573_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5792__C1 _5720_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6029__CLK _6155_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5139__A2 _4333_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4898__A1 _5240_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5924__A _5924_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6179__CLK _6205_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3570__A1 _3592_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_79_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5643__B _5643_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5847__B1 _5905_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2986__C _2986_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6177__D _6177_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5862__A3 _5860_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5075__A1 _5074_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_85_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4275__A _4759_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3086__A0 _6185_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4822__B2 _5118_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4822__A1 _4362_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3625__A2 _3623_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5378__A2 _5377_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3389__A1 _3870_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5783__C1 _4874_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4050__A2 _3832_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3338__B _3499_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4889__A1 _4886_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3010__A0 _6024_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5553__B _5553_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output88_A _3059_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5838__B1 _5031_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3354__A _3838_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _3260_/A VGND VGND VPWR VPWR _4048_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__4169__B _4169_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6087__D _6087_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5853__A3 _5240_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3191_ _3841_/A VGND VGND VPWR VPWR _3343_/A sky130_fd_sc_hd__clkbuf_4
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5066__B2 _5065_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5066__A1 _4422_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4185__A _4405_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3077__A0 _6181_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5901_ _5895_/X _5897_/X _5898_/X _5900_/Y VGND VGND VPWR VPWR _5901_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_81_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4813__A1 _4290_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3616__A2 _4152_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4026__C1 _3157_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5832_ _5263_/A _4501_/X _5819_/A VGND VGND VPWR VPWR _5982_/C sky130_fd_sc_hd__a21oi_4
XANTENNA__5369__A2 _4859_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5763_ _5190_/X _5761_/Y _5762_/Y _4948_/A VGND VGND VPWR VPWR _5763_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4041__A2 _3347_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2975_ _6197_/Q VGND VGND VPWR VPWR _5998_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_4714_ _6048_/Q _4629_/X _4630_/X _4634_/X _4713_/Y VGND VGND VPWR VPWR _6048_/D
+ sky130_fd_sc_hd__o32a_1
XANTENNA__3248__B _3436_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5694_ _4858_/Y _4859_/X _5692_/Y _5693_/Y VGND VGND VPWR VPWR _5694_/X sky130_fd_sc_hd__o22a_1
X_4645_ _4612_/X _5721_/A _5004_/D _4642_/X _4644_/X VGND VGND VPWR VPWR _4645_/X
+ sky130_fd_sc_hd__o2111a_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5744__A _5744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4576_ _4480_/C _4668_/B _4852_/C _5029_/A VGND VGND VPWR VPWR _4576_/X sky130_fd_sc_hd__a31o_2
XANTENNA__3552__A1 _3956_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3527_ _3773_/A _3588_/B _3527_/C VGND VGND VPWR VPWR _3749_/D sky130_fd_sc_hd__and3_2
XFILLER_1_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3264__A _3754_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3458_ _3835_/A VGND VGND VPWR VPWR _3543_/B sky130_fd_sc_hd__buf_2
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3389_ _3870_/A _3557_/A _3657_/C _3581_/A VGND VGND VPWR VPWR _3522_/A sky130_fd_sc_hd__o211a_1
XANTENNA__5844__A3 _5712_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6177_ _6201_/CLK _6177_/D VGND VGND VPWR VPWR _6177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3855__A2 _3854_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5128_ _6055_/Q _5040_/X _5095_/Y _5127_/Y VGND VGND VPWR VPWR _6055_/D sky130_fd_sc_hd__a2bb2oi_1
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3711__B _3711_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5057__A1 _5052_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3068__A0 _6193_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5059_ _5058_/X _5944_/A _4420_/X _4563_/X _4568_/X VGND VGND VPWR VPWR _5059_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__6006__B1 _5292_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4823__A _5034_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4032__A2 _3787_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5780__A2 _5025_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3791__A1 _3783_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5517__C1 _5516_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4335__A3 _4246_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4740__B1 _4697_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3174__A _3387_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4099__A2 _3551_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5835__A3 _4353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3902__A _3902_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3846__A2 _3733_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3621__B _3679_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output126_A _3027_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5829__A _5829_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4733__A _4769_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6012__A3 _6179_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_1_1_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_2_3_0_CLK/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3349__A _4073_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4023__A2 _3524_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5771__A2 _5166_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3782__A1 _3781_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4430_ _4738_/A _4926_/C _4640_/A _4955_/A VGND VGND VPWR VPWR _5706_/A sky130_fd_sc_hd__o211ai_4
XANTENNA__5876__A1_N _6191_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4731__B1 _4666_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5283__B _6014_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4361_ _5976_/C _5018_/B _4353_/X _5140_/B _4360_/X VGND VGND VPWR VPWR _4361_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3084__A _3084_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6100_ _6197_/CLK _6100_/D VGND VGND VPWR VPWR _6100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3312_ _3383_/A VGND VGND VPWR VPWR _3382_/D sky130_fd_sc_hd__buf_2
X_4292_ _4738_/A VGND VGND VPWR VPWR _4347_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__3515__C _3653_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5826__A3 _4945_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_67_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3243_ _3211_/X _3215_/X _3239_/X _3241_/X _3242_/X VGND VGND VPWR VPWR _3243_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6031_ _6197_/CLK _6031_/D VGND VGND VPWR VPWR _6031_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3837__A2 _3517_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3174_ _3387_/B VGND VGND VPWR VPWR _3440_/B sky130_fd_sc_hd__buf_2
XFILLER_39_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5039__B2 _5038_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3250__C _3440_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4798__B1 _4723_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4643__A _4643_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4262__A2 _4260_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5815_ _5754_/Y _5796_/Y _4393_/X VGND VGND VPWR VPWR _5815_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6003__A3 _6009_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3259__A _3802_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4014__A2 _3475_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5747__C1 _5237_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5762__A2 _5013_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5746_ _5746_/A _5746_/B _5746_/C _5746_/D VGND VGND VPWR VPWR _5746_/Y sky130_fd_sc_hd__nand4_1
XFILLER_10_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4970__B1 _4964_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5677_ _5772_/A _5772_/B _5677_/C VGND VGND VPWR VPWR _5677_/X sky130_fd_sc_hd__and3_1
X_4628_ _6047_/Q _4190_/X _4523_/X _4627_/Y VGND VGND VPWR VPWR _6047_/D sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__5474__A _5508_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4559_ _4584_/A VGND VGND VPWR VPWR _5228_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__4722__B1 _4224_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3425__C _3780_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5640__C _6097_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4789__B1 _4739_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4553__A _4555_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5450__B2 input11/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5450__A1 input19/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3169__A _3278_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5738__C1 _5680_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4005__A2 _4124_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4272__B _4285_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5675__A2_N _5646_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5202__A1 input30/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5202__B2 input14/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6190__D _6190_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4410__C1 _4409_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5753__A2 _5020_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4961__B1 _4945_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3516__A1 _3512_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5505__A2 _5433_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4713__B1 _4712_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3108__S _3116_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3335__C _4074_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput94 _3093_/X VGND VGND VPWR VPWR memory_dmem_response_get[15] sky130_fd_sc_hd__buf_2
XANTENNA__4728__A _4728_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3632__A _3632_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3819__A2 _3775_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4492__A2 _4480_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4229__C1 _4228_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3930_ _4039_/B _3923_/Y _3925_/X _3929_/Y _3685_/X VGND VGND VPWR VPWR _3930_/Y
+ sky130_fd_sc_hd__a311oi_4
XFILLER_51_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5559__A _5559_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5441__A1 _4977_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5441__B2 _6109_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4795__A3 _4793_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3452__B1 _3421_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5278__B _5570_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5992__A2 _5286_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3861_ _3911_/B _3230_/X _3720_/X _4124_/B _3934_/B VGND VGND VPWR VPWR _3861_/Y
+ sky130_fd_sc_hd__a221oi_1
XANTENNA__4182__B _4231_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4401__C1 _4769_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3792_ _3816_/A _3806_/B _3792_/C _3792_/D VGND VGND VPWR VPWR _3792_/X sky130_fd_sc_hd__or4_1
X_5600_ _5600_/A VGND VGND VPWR VPWR _6159_/D sky130_fd_sc_hd__clkbuf_1
X_5531_ _5531_/A _5531_/B VGND VGND VPWR VPWR _5532_/A sky130_fd_sc_hd__and2_1
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3807__A _3807_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5294__A _5294_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_105_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5725__C _5725_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3507__A1 _3478_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5462_ input22/X _5437_/A _5439_/A input14/X VGND VGND VPWR VPWR _5772_/C sky130_fd_sc_hd__a22o_1
XANTENNA__4704__B1 _5188_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4413_ _4574_/A VGND VGND VPWR VPWR _5148_/D sky130_fd_sc_hd__buf_2
X_5393_ _5436_/A _5392_/X _4201_/A VGND VGND VPWR VPWR _5420_/A sky130_fd_sc_hd__o21a_2
X_4344_ _4780_/A VGND VGND VPWR VPWR _4345_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4638__A _4759_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_113_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4275_ _4759_/C VGND VGND VPWR VPWR _4769_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4468__C1 _4948_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6014_ _6014_/A _6014_/B _6014_/C VGND VGND VPWR VPWR _6015_/A sky130_fd_sc_hd__and3_1
X_3226_ _3226_/A VGND VGND VPWR VPWR _3606_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3157_ _3858_/A _3278_/A _3157_/C _3586_/A VGND VGND VPWR VPWR _3157_/X sky130_fd_sc_hd__or4_4
XANTENNA__3691__B1 _3624_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3088_ _6186_/Q _6078_/Q _3094_/S VGND VGND VPWR VPWR _3089_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5469__A _5469_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4373__A _4643_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5188__B _5188_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4092__B _4092_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3994__A1 _3614_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3994__B2 _3648_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4538__A3 _4297_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5196__B1 _4494_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5735__A2 _4556_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4943__B1 _5878_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5729_ _5811_/A _5729_/B VGND VGND VPWR VPWR _5729_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3717__A _4048_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3436__B _3436_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5651__B _5651_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_104_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5120__B1 _5667_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4474__A2 _4865_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5671__A1 _5664_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6185__D _6185_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3682__B1 _3749_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4283__A _4283_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5974__A2 _5757_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4631__C1 _4804_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3985__A1 _3962_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5187__B1 _4574_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3737__A1 _3519_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3737__B2 _3871_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4162__B2 _3517_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4162__A1 _4158_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_68_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4458__A _4533_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5111__B1 _5050_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4060_ _3335_/X _3847_/X _4059_/X _3868_/X VGND VGND VPWR VPWR _4060_/X sky130_fd_sc_hd__o31a_1
XANTENNA__4177__B _4230_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5662__A1 _5060_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4465__A2 _4209_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6095__D _6095_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3011_ _3011_/A VGND VGND VPWR VPWR _3011_/X sky130_fd_sc_hd__clkbuf_1
X_4962_ _4783_/X _4827_/A _4552_/X _4856_/A VGND VGND VPWR VPWR _4962_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5965__A2 _5963_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4893_ _5228_/A VGND VGND VPWR VPWR _5237_/A sky130_fd_sc_hd__buf_4
X_3913_ _3593_/D _3653_/A _4073_/A _3525_/X _4149_/A VGND VGND VPWR VPWR _3913_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3976__A1 _3701_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5178__B1 _5191_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3844_ _3893_/C VGND VGND VPWR VPWR _3844_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__5717__A2 _5152_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4925__B1 _4924_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5193__A3 _4697_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3537__A _3537_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3775_ _3815_/B _3765_/X _3774_/X _3764_/X VGND VGND VPWR VPWR _3775_/Y sky130_fd_sc_hd__a22oi_2
XANTENNA__6062__CLK _6201_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4940__A3 _5971_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5514_ _5514_/A _5531_/B VGND VGND VPWR VPWR _5515_/A sky130_fd_sc_hd__and2_1
XFILLER_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5445_ _5445_/A VGND VGND VPWR VPWR _5445_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4153__A1 _3761_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5350__A0 _6046_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_120_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3900__A1 _3859_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5376_ _6098_/Q _5381_/B VGND VGND VPWR VPWR _5376_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_113_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4368__A _4832_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3272__A _3272_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4327_ _4527_/C _4527_/D _4358_/A _4878_/D VGND VGND VPWR VPWR _5667_/A sky130_fd_sc_hd__and4_2
XFILLER_86_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4258_ _4696_/A VGND VGND VPWR VPWR _4259_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5653__A1 _4855_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3209_ _3754_/B VGND VGND VPWR VPWR _3864_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_28_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3664__B1 _3662_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4189_ _4189_/A VGND VGND VPWR VPWR _5646_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4815__B _4929_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5956__A2 _5431_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5169__B1 _4652_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4916__B1 _4699_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3447__A _3621_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4144__A1 _3910_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5892__A1 _4959_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4144__B2 _3603_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3352__C1 _3351_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5381__B _5381_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3182__A _3870_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_78_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5644__A1 _4975_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3910__A _3910_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3655__B1 _3654_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5601__S _5605_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3407__B1 _3374_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5947__A2 _5395_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3121__S _3127_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3958__A1 _3679_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4080__B1 _4076_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6085__CLK _6203_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4907__B1 _4906_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3357__A _3891_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3560_ _3548_/X _3554_/X _3628_/A _3559_/Y VGND VGND VPWR VPWR _3560_/X sky130_fd_sc_hd__a211o_1
XANTENNA__5275__C _6014_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5230_ _4353_/X _5123_/C _4487_/Y _5167_/A _5755_/C VGND VGND VPWR VPWR _5230_/X
+ sky130_fd_sc_hd__o221a_1
X_3491_ _3491_/A VGND VGND VPWR VPWR _3959_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_102_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5883__A1 _5211_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5291__B _6205_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5883__B2 _4680_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3894__B1 _3218_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4188__A _4188_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5161_ input29/X _4804_/X _5042_/A input13/X VGND VGND VPWR VPWR _5161_/X sky130_fd_sc_hd__a22o_1
XFILLER_96_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4619__C _4852_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4112_ _3557_/A _4042_/A _3648_/B _4152_/A VGND VGND VPWR VPWR _4112_/X sky130_fd_sc_hd__a22o_1
X_5092_ _5529_/A VGND VGND VPWR VPWR _5092_/X sky130_fd_sc_hd__buf_2
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4043_ _3967_/A _4042_/C _3279_/A _3648_/Y VGND VGND VPWR VPWR _4043_/X sky130_fd_sc_hd__o31a_1
XFILLER_83_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3646__B1 _3645_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4989__A3 _4193_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_92_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5938__A2 _5913_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5399__B1 _5398_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5994_ _5998_/C _5998_/B _5986_/Y VGND VGND VPWR VPWR _5994_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4945_ _4945_/A VGND VGND VPWR VPWR _4945_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_91_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4354__C _4358_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3949__A1 _4124_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4073__D _4073_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4071__B1 _3695_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4876_ _4876_/A VGND VGND VPWR VPWR _5152_/C sky130_fd_sc_hd__clkbuf_8
XANTENNA__4651__A _4780_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3827_ _5388_/B _6031_/Q _3826_/X VGND VGND VPWR VPWR _6031_/D sky130_fd_sc_hd__a21o_1
X_3758_ _3959_/D _3815_/B _3756_/X _3792_/C VGND VGND VPWR VPWR _3816_/D sky130_fd_sc_hd__a31o_1
XANTENNA__5571__B1 _6100_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3689_ _3658_/X _3680_/A _3688_/X VGND VGND VPWR VPWR _3689_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__5482__A _5482_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5428_ _5508_/A VGND VGND VPWR VPWR _5468_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3885__B1 _4042_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4677__A2 _4669_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5359_ _6049_/Q _6093_/Q _5361_/S VGND VGND VPWR VPWR _5360_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4834__C1 _4794_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3637__B1 _3636_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4264__C _4264_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5929__A2 _4967_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4062__B1 _4061_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_90_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4038__A2_N _4037_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5376__B _5381_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3177__A _3603_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3905__A _4092_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4117__A1 _4116_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_99_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5865__A1 _5863_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3116__S _3116_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5331__S _5339_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_CLK clkbuf_4_7_0_CLK/A VGND VGND VPWR VPWR _6074_/CLK sky130_fd_sc_hd__clkbuf_2
XANTENNA__5250__C1 _5152_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4053__B1 _3588_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2991_ _3060_/S _6013_/B _6060_/Q VGND VGND VPWR VPWR _2991_/X sky130_fd_sc_hd__o21a_2
X_4730_ _5078_/B _4488_/X _5687_/A _4923_/A VGND VGND VPWR VPWR _4730_/Y sky130_fd_sc_hd__o211ai_4
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4471__A _4926_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3800__B1 _3464_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4661_ _4661_/A VGND VGND VPWR VPWR _4661_/X sky130_fd_sc_hd__buf_4
XANTENNA__5286__B _5286_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5002__C1 _4998_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3612_ _3871_/A _4083_/B _3680_/A _3612_/D VGND VGND VPWR VPWR _3612_/X sky130_fd_sc_hd__or4_1
XANTENNA__3087__A _3087_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4592_ _4614_/A VGND VGND VPWR VPWR _4668_/A sky130_fd_sc_hd__clkbuf_2
X_3543_ _3847_/A _3543_/B VGND VGND VPWR VPWR _3543_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__4371__A4 _4309_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3815__A _3815_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_88_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3474_ _4092_/A VGND VGND VPWR VPWR _3871_/A sky130_fd_sc_hd__buf_4
XANTENNA__4108__A1 _4105_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5733__C _5813_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6100__CLK _6197_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5213_ _4580_/A _4878_/A _4815_/C _4862_/A VGND VGND VPWR VPWR _5213_/X sky130_fd_sc_hd__a31o_4
XANTENNA__5856__A1 _5850_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5856__B2 _5855_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6193_ _6196_/CLK _6193_/D VGND VGND VPWR VPWR _6193_/Q sky130_fd_sc_hd__dfxtp_1
X_5144_ _4243_/A _4362_/A _4247_/A _4364_/A _4555_/B VGND VGND VPWR VPWR _5145_/A
+ sky130_fd_sc_hd__o311a_2
XANTENNA__3026__S _3032_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_96_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5608__A1 _6031_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4646__A _4854_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5075_ _5074_/X _4959_/X _5058_/X _4875_/X VGND VGND VPWR VPWR _5075_/Y sky130_fd_sc_hd__o31ai_2
XANTENNA__3619__B1 _3868_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_84_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4026_ _3470_/X _4048_/B _3882_/C _4025_/Y _3157_/X VGND VGND VPWR VPWR _4026_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__5084__A2 _5072_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4831__A2 _4843_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4143__C_N _3645_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3634__A3 _3756_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5241__C1 _4824_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5977_ _5755_/A _5680_/A _4891_/X _4916_/X VGND VGND VPWR VPWR _5977_/X sky130_fd_sc_hd__a31o_1
XFILLER_52_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4381__A _4578_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4595__A1 _4666_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4928_ _4928_/A VGND VGND VPWR VPWR _5680_/C sky130_fd_sc_hd__buf_2
XANTENNA__5792__B1 _5782_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5139__A3 _4518_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4859_ _5757_/B _4859_/B _4859_/C _4859_/D VGND VGND VPWR VPWR _4859_/X sky130_fd_sc_hd__and4b_2
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4898__A2 _5240_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5924__B _5924_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3570__A2 _3956_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5643__C _6123_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_106_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5847__A1 _6102_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4556__A _4556_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5075__A2 _4959_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_75_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3086__A1 _6077_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4822__A2 _4363_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6193__D _6193_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5387__A _5387_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3389__A2 _3557_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4291__A _4759_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5783__B1 _5782_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4050__A3 _4089_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4889__A2 _5732_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5535__B1 _5491_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6123__CLK _6123_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5326__S _5328_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3010__A1 _6156_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6011__A _6011_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5838__A1 _4998_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3849__B1 _3647_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _3781_/A VGND VGND VPWR VPWR _3841_/A sky130_fd_sc_hd__buf_2
XFILLER_78_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3370__A _3904_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4466__A _4835_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_66_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5066__A2 _4423_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3077__A1 _6073_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5900_ _5006_/X _5026_/X _5899_/X _5235_/X VGND VGND VPWR VPWR _5900_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_81_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4813__A2 _4617_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4274__B1 _4273_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5831_ _5228_/X _5825_/Y _5828_/X _5830_/Y VGND VGND VPWR VPWR _5831_/Y sky130_fd_sc_hd__o22ai_4
XANTENNA__4026__B1 _4025_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5369__A3 _4859_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5223__C1 _5042_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5762_ _4362_/X _5013_/S _4364_/X _5107_/A _5152_/B VGND VGND VPWR VPWR _5762_/Y
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA__5774__B1 _5769_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5297__A _5365_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4041__A3 _3533_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4713_ _4664_/Y _4683_/Y _4952_/B _4712_/Y VGND VGND VPWR VPWR _4713_/Y sky130_fd_sc_hd__a31oi_2
X_5693_ _5720_/A _5720_/B _4856_/A _4563_/A VGND VGND VPWR VPWR _5693_/Y sky130_fd_sc_hd__a31oi_2
X_4644_ _4827_/A VGND VGND VPWR VPWR _4644_/X sky130_fd_sc_hd__clkbuf_4
X_4575_ _4878_/D VGND VGND VPWR VPWR _4852_/C sky130_fd_sc_hd__buf_2
XFILLER_116_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3552__A2 _3500_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3545__A _3773_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3526_ _3526_/A VGND VGND VPWR VPWR _3773_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3457_ _3457_/A VGND VGND VPWR VPWR _3457_/X sky130_fd_sc_hd__buf_4
X_3388_ _3582_/C _3802_/D VGND VGND VPWR VPWR _3581_/A sky130_fd_sc_hd__nor2_4
XFILLER_69_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6176_ _6176_/CLK _6176_/D VGND VGND VPWR VPWR _6176_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4376__A _4860_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5127_ _5127_/A _5127_/B _5220_/C VGND VGND VPWR VPWR _5127_/Y sky130_fd_sc_hd__nand3_4
XFILLER_57_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5058_ _5096_/A _4777_/X _4778_/X _5079_/C _5687_/B VGND VGND VPWR VPWR _5058_/X
+ sky130_fd_sc_hd__o311a_2
XANTENNA__5057__A2 _5056_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3280__A _3864_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3068__A1 _6069_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4009_ _4003_/Y _4005_/X _4008_/X _3479_/X _3577_/X VGND VGND VPWR VPWR _4009_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6006__A1 _6206_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4017__B1 _3161_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5765__B1 _5175_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5000__A _5000_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6146__CLK _6146_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4032__A3 _3763_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3791__A2 _3790_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5517__B1 _5447_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5890__A2_N _4878_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3455__A _3802_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4740__A1 _4707_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4335__A4 _4309_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6188__D _6188_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3902__B _4074_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input32_A memory_dmem_request_put[58] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3621__C _3621_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3190__A _3781_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4256__B1 _4255_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output119_A _3080_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5829__B _5829_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4008__B1 _4007_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6012__A4 _6013_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4023__A3 _3975_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3782__A2 _3380_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3365__A _3461_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4731__A1 _4692_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4360_ _4243_/X _4293_/B _4910_/A _4865_/C _4668_/B VGND VGND VPWR VPWR _4360_/X
+ sky130_fd_sc_hd__o311a_4
XANTENNA__5283__C _5283_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3311_ _3461_/A _3311_/B VGND VGND VPWR VPWR _3383_/A sky130_fd_sc_hd__and2_1
XANTENNA__6098__D _6098_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4291_ _4759_/C VGND VGND VPWR VPWR _4738_/A sky130_fd_sc_hd__buf_2
XANTENNA__3515__D _3797_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5580__A _5580_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3242_ _3707_/A VGND VGND VPWR VPWR _3242_/X sky130_fd_sc_hd__buf_2
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _6045_/CLK _6030_/D VGND VGND VPWR VPWR _6030_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4495__B1 _4494_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3837__A3 _3833_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3173_ _3161_/X _3170_/X _3359_/A VGND VGND VPWR VPWR _3173_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4196__A input7/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6019__CLK _6155_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_94_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4924__A _4924_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4798__B2 _4797_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5995__B1 _6200_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6169__CLK _6197_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5747__B1 _5746_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5814_ _5813_/Y _4964_/X _5735_/X VGND VGND VPWR VPWR _5814_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_35_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3259__B _3437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4014__A3 _3499_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5745_ _5745_/A _5745_/B _5745_/C VGND VGND VPWR VPWR _5746_/C sky130_fd_sc_hd__and3_2
XANTENNA__5755__A _5755_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4970__A1 _4958_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5983__A1_N _5970_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5676_ _5676_/A VGND VGND VPWR VPWR _5676_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4627_ _4558_/Y _4569_/X _4974_/C _4626_/X VGND VGND VPWR VPWR _4627_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__3275__A _3513_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4722__A1 _6129_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4558_ _4542_/X _4557_/X _4252_/X VGND VGND VPWR VPWR _4558_/Y sky130_fd_sc_hd__a21oi_4
X_4489_ _4769_/B VGND VGND VPWR VPWR _4929_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3509_ _3509_/A _3589_/B VGND VGND VPWR VPWR _3509_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__3930__C1 _3685_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ _6197_/CLK _6159_/D VGND VGND VPWR VPWR _6159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3830__B_N _3654_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5640__D _5640_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_85_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4789__B2 _5836_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4789__A1 _4786_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5450__A2 _5437_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5738__B1 _4385_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4005__A3 _3223_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5202__A2 _4804_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4410__B1 _4403_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5753__A3 _4708_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4961__A1 _5240_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3185__A _3442_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3516__A2 _3410_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4713__A1 _4664_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5910__B1 _4744_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3921__C1 _3920_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput84 _2987_/X VGND VGND VPWR VPWR RDY_memory_dmem_request_put sky130_fd_sc_hd__buf_2
Xoutput95 _3095_/X VGND VGND VPWR VPWR memory_dmem_response_get[16] sky130_fd_sc_hd__buf_2
XFILLER_95_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4229__B1 _5044_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4744__A _4744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5977__B1 _4916_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3988__C1 _3583_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5441__A2 _5412_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3452__A1 _3359_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3860_ _3860_/A VGND VGND VPWR VPWR _3934_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__4182__C _4231_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4401__B1 _4533_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_72_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3791_ _3783_/X _3790_/Y _3707_/X VGND VGND VPWR VPWR _3792_/D sky130_fd_sc_hd__a21oi_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5530_ _5523_/X _4285_/B _5529_/X _5491_/X _6135_/Q VGND VGND VPWR VPWR _5531_/A
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3807__B _3814_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5294__B input2/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5461_ _5461_/A VGND VGND VPWR VPWR _6113_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4412_ _4614_/A _4543_/A VGND VGND VPWR VPWR _4574_/A sky130_fd_sc_hd__nand2_4
XANTENNA__3095__A _3095_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4704__A1 _4483_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5901__B1 _5898_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3507__A2 _3505_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5392_ input7/X input8/X _5392_/C _5438_/D VGND VGND VPWR VPWR _5392_/X sky130_fd_sc_hd__and4b_1
XFILLER_99_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4343_ _4555_/B VGND VGND VPWR VPWR _4780_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4274_ _4266_/A _4272_/X _4273_/Y _4209_/A VGND VGND VPWR VPWR _4759_/C sky130_fd_sc_hd__o2bb2ai_4
XFILLER_100_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3225_ _3440_/A _3366_/A VGND VGND VPWR VPWR _3621_/A sky130_fd_sc_hd__or2_2
XANTENNA__5665__C1 _4589_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4468__B1 _4918_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6013_ _6207_/Q _6013_/B _6013_/C VGND VGND VPWR VPWR _6014_/C sky130_fd_sc_hd__nand3_1
XFILLER_100_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3156_ _3603_/D VGND VGND VPWR VPWR _3586_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3691__A1 _3684_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4654__A _4654_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3087_ _3087_/A VGND VGND VPWR VPWR _3087_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3979__C1 _4116_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5188__C _5188_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4092__C _4092_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3994__A2 _4149_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5196__A1 _5187_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4943__A1 _5755_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_109_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3989_ _3932_/Y _3720_/A _3319_/X _3802_/X VGND VGND VPWR VPWR _3989_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5735__A3 _5050_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5728_ _6112_/Q _4511_/X _5676_/A _5727_/X VGND VGND VPWR VPWR _5729_/B sky130_fd_sc_hd__o211a_1
X_5659_ _5018_/A _4864_/Y _4865_/Y _4422_/A _4699_/X VGND VGND VPWR VPWR _5661_/A
+ sky130_fd_sc_hd__a311oi_4
XFILLER_104_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_2_1_0_CLK/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5656__C1 _4420_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5120__A1 _5711_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4474__A3 _4472_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3238__A_N _3509_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3682__A1 _3668_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5671__A2 _5670_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4564__A _4788_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5959__B1 _4957_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4631__B1 _4718_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3985__A2 _3583_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5187__A1 _5755_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5187__B2 _5976_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3737__A2 _3847_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5395__A _5395_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3119__S _3127_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4147__C1 _3621_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5895__C1 _5755_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4739__A _4739_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4698__B1 _4819_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4162__A2 _4159_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3643__A _3643_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4458__B _5008_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5111__B2 _4890_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5111__A1 _4693_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4177__C _4230_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_76_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5662__A2 _5658_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3010_ _6024_/Q _6156_/Q _3010_/S VGND VGND VPWR VPWR _3011_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4622__B1 _4619_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4961_ _5240_/A _4754_/X _4945_/X _4960_/X VGND VGND VPWR VPWR _4961_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_64_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5965__A3 _5964_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4193__B _4225_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3912_ _3708_/A _3847_/C _3633_/A _3515_/B VGND VGND VPWR VPWR _4143_/A sky130_fd_sc_hd__o22a_1
X_4892_ _5976_/A _4840_/X _4891_/X _4541_/A VGND VGND VPWR VPWR _4892_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3976__A2 _3340_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5178__A1 _4772_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3843_ _3594_/X _3320_/Y _3699_/A _3842_/X VGND VGND VPWR VPWR _3843_/Y sky130_fd_sc_hd__a211oi_1
XANTENNA__4925__A1 _5123_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6207__CLK _6207_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3537__B _3537_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3774_ _3549_/X _3881_/B _3195_/A _3633_/Y VGND VGND VPWR VPWR _3774_/X sky130_fd_sc_hd__a31o_1
XFILLER_118_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5513_ _5495_/X _4720_/X _5498_/X _6129_/Q _5503_/A VGND VGND VPWR VPWR _5514_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_9_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4940__A4 _5878_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5444_ _5444_/A VGND VGND VPWR VPWR _5444_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4153__A2 _3572_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5350__A1 _6089_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4649__A _4649_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3553__A _3553_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3361__B1 _3208_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5375_ _5368_/X _5371_/Y _6011_/B _5374_/X VGND VGND VPWR VPWR _6097_/D sky130_fd_sc_hd__o211a_1
XFILLER_113_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4326_ _4354_/D VGND VGND VPWR VPWR _4878_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__3900__A2 _3653_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4257_ _4700_/A VGND VGND VPWR VPWR _4696_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5653__A2 _4673_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3208_ _3509_/A VGND VGND VPWR VPWR _3208_/X sky130_fd_sc_hd__buf_2
X_4188_ _4188_/A VGND VGND VPWR VPWR _4189_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3664__A1 _3536_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3139_ _3748_/A VGND VGND VPWR VPWR _3139_/X sky130_fd_sc_hd__buf_2
XANTENNA__4815__C _4815_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4613__B1 _4345_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5810__C1 _5809_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5169__A1 _4740_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4916__A1 _5013_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3728__A _3822_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3447__B _3527_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4129__C1 _3350_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4144__A2 _3299_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4559__A _4584_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3352__B1 _3340_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5892__A2 _5890_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6196__D _6196_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5644__A2 _5444_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3910__B _3910_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3655__A1 _3652_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3407__A1 _3403_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3958__A2 _4124_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4080__A1 _3300_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output101_A _3106_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4080__B2 _4079_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5122__A1_N _5116_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4907__A1 input23/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4907__B2 _4717_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6014__A _6014_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3490_ _3536_/A _3975_/B _3359_/C _3488_/X _3489_/X VGND VGND VPWR VPWR _3490_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_6_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3373__A _3966_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5883__A2 _5878_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3894__A1 _3178_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_5160_ _5822_/A VGND VGND VPWR VPWR _5166_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__5291__C _6179_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_110_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4111_ _3967_/A _3495_/X _3674_/C _4110_/Y VGND VGND VPWR VPWR _4111_/X sky130_fd_sc_hd__o31a_1
XFILLER_78_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5091_ _5162_/A VGND VGND VPWR VPWR _5529_/A sky130_fd_sc_hd__buf_2
XFILLER_110_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4042_ _4042_/A _4073_/A _4042_/C _4042_/D VGND VGND VPWR VPWR _4042_/X sky130_fd_sc_hd__or4_1
XFILLER_68_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3646__A1 _3548_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5399__B2 _6101_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5399__A1 input9/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5993_ _5998_/A _5571_/X _5410_/X VGND VGND VPWR VPWR _6199_/D sky130_fd_sc_hd__o21a_1
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4944_ _4680_/X _4761_/X _4878_/Y _4618_/X VGND VGND VPWR VPWR _4944_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4354__D _4354_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3949__A2 _3720_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4331__A1_N _4527_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4071__A1 _4067_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4875_ _4875_/A VGND VGND VPWR VPWR _4875_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3548__A _3571_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3826_ _3825_/Y _3638_/Y _3816_/B _3778_/X _3787_/X VGND VGND VPWR VPWR _3826_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_118_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_3757_ _3689_/Y _3663_/X _3282_/A VGND VGND VPWR VPWR _3792_/C sky130_fd_sc_hd__a21boi_4
XANTENNA__5571__A1 _6199_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5859__C1 _5944_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3688_ _3603_/X _3686_/X _3687_/Y VGND VGND VPWR VPWR _3688_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4379__A _4379_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3283__A _3934_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5427_ input15/X _5412_/X _5431_/B _5398_/X _6107_/Q VGND VGND VPWR VPWR _5429_/A
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3885__A1 _3773_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5358_ _5358_/A VGND VGND VPWR VPWR _6092_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4309_ _4309_/A VGND VGND VPWR VPWR _4309_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5289_ _5285_/X _5286_/Y _5288_/X VGND VGND VPWR VPWR _5289_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4834__B1 _4833_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3637__A1 _3524_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5003__A _5667_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_74_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4264__D _4309_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4062__A1 _3967_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3458__A _3835_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5011__B1 _4584_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4770__C1 _5005_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5673__A _5673_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5392__B input8/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input62_A memory_dmem_request_put[88] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4289__A _4578_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3193__A _3780_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4117__A2 _3699_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5865__A2 _5864_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output149_A _3014_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5612__S _5616_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4825__B1 _4824_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_65_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6052__CLK _6196_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6009__A _6009_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_73_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5250__B1 _5078_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4053__A1 _3910_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2990_ _6202_/Q _6205_/Q _6179_/Q VGND VGND VPWR VPWR _6013_/B sky130_fd_sc_hd__and3_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3368__A _3631_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3800__A1 _3799_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5691__A1_N _4570_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4660_ _5188_/D _4929_/B _4580_/A VGND VGND VPWR VPWR _4672_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__5002__B1 _4461_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3611_ _3611_/A VGND VGND VPWR VPWR _4083_/B sky130_fd_sc_hd__buf_2
X_4591_ _5971_/B _4437_/Y _4572_/X _4369_/Y VGND VGND VPWR VPWR _4591_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__3564__B1 _3528_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3542_ _3507_/Y _3540_/Y _3453_/X _6019_/Q _3541_/X VGND VGND VPWR VPWR _6019_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3473_ _3870_/B VGND VGND VPWR VPWR _3674_/C sky130_fd_sc_hd__buf_4
XANTENNA__4108__A2 _4107_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3815__B _3815_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4199__A _4717_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5212_ _5211_/X _4552_/X _4953_/X _5179_/A _5106_/X VGND VGND VPWR VPWR _5212_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__5856__A2 _5851_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_69_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6192_ _6196_/CLK _6192_/D VGND VGND VPWR VPWR _6192_/Q sky130_fd_sc_hd__dfxtp_1
X_5143_ _5097_/X _4459_/X _5743_/B _4945_/X _4420_/A VGND VGND VPWR VPWR _5150_/A
+ sky130_fd_sc_hd__a41o_1
XANTENNA__4927__A _4927_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5069__B1 _4387_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3831__A _3831_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5074_ _4865_/D _4865_/A _4946_/A _5078_/D VGND VGND VPWR VPWR _5074_/X sky130_fd_sc_hd__o211a_4
XANTENNA__4816__B1 _4819_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3619__A1 _3749_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4025_ _3895_/A _3457_/A _3205_/X _3911_/A VGND VGND VPWR VPWR _4025_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_64_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5241__B1 _4618_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5976_ _5976_/A _5976_/B _5976_/C VGND VGND VPWR VPWR _5976_/X sky130_fd_sc_hd__and3_1
XFILLER_80_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4595__A2 _4590_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4927_ _4927_/A VGND VGND VPWR VPWR _4927_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__3278__A _3278_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5792__A1 _4927_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_100_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4858_ _4859_/D _5203_/A _6139_/Q VGND VGND VPWR VPWR _4858_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_60_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3809_ _3766_/Y _3808_/Y _3492_/X VGND VGND VPWR VPWR _3809_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4789_ _4786_/X _5062_/A _4739_/A _5836_/A VGND VGND VPWR VPWR _4789_/X sky130_fd_sc_hd__o22a_2
XFILLER_4_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5493__A _5493_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4898__A3 _5878_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5847__A2 _4807_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__6075__CLK _6176_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5075__A3 _5058_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4572__A _4643_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5232__B1 _4765_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_70_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5783__A1 _5712_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3243__C1 _3242_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3188__A _3233_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5535__A1 _5523_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5535__B2 _6137_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4889__A3 _4888_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4743__C1 _4742_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6011__B _6011_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5838__A2 _5833_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3127__S _3127_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3849__A1 _4092_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4747__A _4747_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3651__A _3711_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5342__S _5350_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_93_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4274__B2 _4209_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5471__B1 _5256_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5578__A _5578_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5830_ _4875_/X _5018_/Y _5829_/X _5237_/A VGND VGND VPWR VPWR _5830_/Y sky130_fd_sc_hd__o31ai_2
XANTENNA__4026__A1 _3470_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4482__A _4482_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__5223__B1 _5431_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5761_ _5761_/A _5761_/B _5761_/C _5761_/D VGND VGND VPWR VPWR _5761_/Y sky130_fd_sc_hd__nand4_2
XANTENNA__5774__A1 _5676_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4712_ _4685_/X _4711_/X _4503_/A VGND VGND VPWR VPWR _4712_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3785__B1 _3784_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3098__A _3098_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5692_ _4771_/X _4773_/Y _4374_/X VGND VGND VPWR VPWR _5692_/Y sky130_fd_sc_hd__a21oi_1
X_4643_ _4643_/A VGND VGND VPWR VPWR _4827_/A sky130_fd_sc_hd__clkbuf_2
X_4574_ _4574_/A VGND VGND VPWR VPWR _4574_/X sky130_fd_sc_hd__buf_4
X_3525_ _3525_/A VGND VGND VPWR VPWR _3525_/X sky130_fd_sc_hd__buf_4
XANTENNA__3545__B _4092_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6098__CLK _6207_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_116_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3037__S _3043_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3456_ _3966_/C VGND VGND VPWR VPWR _3457_/A sky130_fd_sc_hd__clkbuf_4
X_3387_ _3311_/B _3387_/B VGND VGND VPWR VPWR _3802_/D sky130_fd_sc_hd__and2b_1
XFILLER_69_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4657__A _4657_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3561__A _3707_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6175_ _6201_/CLK _6175_/D VGND VGND VPWR VPWR _6175_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4376__B _4860_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_97_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5126_ _4252_/X _5124_/A _5124_/Y _5175_/A VGND VGND VPWR VPWR _5127_/B sky130_fd_sc_hd__o211ai_2
XFILLER_29_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5057_ _5052_/Y _5056_/Y _4252_/X VGND VGND VPWR VPWR _5057_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_57_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4008_ _3183_/X _3534_/X _4006_/Y _4007_/X VGND VGND VPWR VPWR _4008_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5462__B1 _5439_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6006__A2 _5382_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5214__B1 _5743_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4392__A _4767_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4017__A1 _3990_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_80_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5959_ _5680_/A _4891_/X _5755_/A _4957_/A VGND VGND VPWR VPWR _5959_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5765__A1 _5735_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3776__B1 _3479_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5517__A1 _6130_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4740__A2 _4350_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_6_0_CLK clkbuf_4_7_0_CLK/A VGND VGND VPWR VPWR _6202_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_121_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3621__D _3621_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input25_A memory_dmem_request_put[51] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4256__A1 _4307_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5398__A _5503_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5829__C _5829_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4008__A1 _3183_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5205__B1 _5013_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4023__A4 _3612_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5337__S _5339_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4731__A2 _4353_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output93_A _3091_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3310_ _3614_/A VGND VGND VPWR VPWR _3867_/A sky130_fd_sc_hd__clkbuf_4
X_4290_ _5211_/A _4815_/C _4259_/A _4725_/A VGND VGND VPWR VPWR _4290_/Y sky130_fd_sc_hd__o211ai_4
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4477__A _4759_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_98_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3381__A _4034_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3241_ _3476_/B VGND VGND VPWR VPWR _3241_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__4495__A1 _4469_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5692__B1 _4374_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3172_ _4044_/B _3282_/A VGND VGND VPWR VPWR _3359_/A sky130_fd_sc_hd__and2_2
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5995__A1 _5984_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5747__A1 _5709_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5813_ _5955_/D _5813_/B _5813_/C VGND VGND VPWR VPWR _5813_/Y sky130_fd_sc_hd__nand3_1
XFILLER_34_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3758__B1 _3792_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5744_ _5744_/A VGND VGND VPWR VPWR _5745_/B sky130_fd_sc_hd__buf_2
XFILLER_108_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5755__B _5755_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4970__A2 _4963_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5675_ _6181_/Q _5646_/X _5651_/Y _5674_/Y VGND VGND VPWR VPWR _6181_/D sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__3556__A _4105_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4626_ _4570_/Y _4571_/X _4596_/Y _4625_/Y VGND VGND VPWR VPWR _4626_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3275__B _3275_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4557_ _4457_/X _4548_/Y _4554_/X _4556_/X VGND VGND VPWR VPWR _4557_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4722__A2 _4975_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4488_ _4878_/A VGND VGND VPWR VPWR _4488_/X sky130_fd_sc_hd__buf_4
XANTENNA__3930__B1 _3929_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3508_ _3508_/A VGND VGND VPWR VPWR _3508_/X sky130_fd_sc_hd__buf_2
XFILLER_1_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3291__A _3387_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3439_ _4149_/D _3660_/B _4092_/D _3732_/D _3438_/X VGND VGND VPWR VPWR _3439_/X
+ sky130_fd_sc_hd__o41a_2
XANTENNA__4387__A _4642_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5683__B1 _5060_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _6201_/CLK _6158_/D VGND VGND VPWR VPWR _6158_/Q sky130_fd_sc_hd__dfxtp_1
X_5109_ _5140_/B _4735_/Y _5050_/Y _5048_/X VGND VGND VPWR VPWR _5109_/Y sky130_fd_sc_hd__a22oi_1
XANTENNA__3694__C1 _3522_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_6089_ _6176_/CLK _6089_/D VGND VGND VPWR VPWR _6089_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6113__CLK _6123_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4789__A2 _5062_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3997__B1 _3781_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_82_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5738__A1 _5903_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4005__A4 _4004_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6208__150 VGND VGND VPWR VPWR _6208__150/HI memory_imem_response_get[22] sky130_fd_sc_hd__conb_1
XFILLER_13_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4410__A1 _4398_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4850__A _4850_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__4961__A2 _4754_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5753__A4 _4891_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6199__D _6199_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_107_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5910__A1 _5020_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3516__A3 _3320_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4713__A2 _4683_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_122_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3921__B1 _3918_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4297__A _4527_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput85 _2991_/X VGND VGND VPWR VPWR RDY_memory_dmem_response_get sky130_fd_sc_hd__buf_2
XFILLER_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput96 _3098_/X VGND VGND VPWR VPWR memory_dmem_response_get[17] sky130_fd_sc_hd__buf_2
XFILLER_63_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5426__B1 _5528_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output131_A _2995_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4229__A1 _4716_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_91_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5977__A1 _5755_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3988__B1 _3537_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5441__A3 _5440_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3452__A2 _3408_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4182__D _4231_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4760__A _4876_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4401__A1 _4329_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_3790_ _3607_/X _3733_/Y _4146_/A VGND VGND VPWR VPWR _3790_/Y sky130_fd_sc_hd__o21ai_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__3185__B_N _3440_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3376__A _3749_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3807__C _4044_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5460_ _5460_/A _5468_/B VGND VGND VPWR VPWR _5461_/A sky130_fd_sc_hd__and2_1
XANTENNA__5294__C _6013_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_117_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_4411_ _4442_/A VGND VGND VPWR VPWR _4614_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4704__A2 _4485_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5901__A1 _5895_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__5901__B2 _5900_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_5391_ _5438_/D input7/X _4225_/A VGND VGND VPWR VPWR _5436_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__5591__A _5591_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__3912__B1 _3633_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4342_ _4340_/Y _5818_/S _4341_/Y VGND VGND VPWR VPWR _4555_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__5114__C1 _5113_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_4273_ _6135_/Q VGND VGND VPWR VPWR _4273_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_113_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3224_ _3226_/A VGND VGND VPWR VPWR _3366_/A sky130_fd_sc_hd__buf_2
XANTENNA__5665__B1 _4869_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4468__B2 _4464_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__4468__A1 _4459_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__6136__CLK _6146_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_6012_ _6202_/Q _6205_/Q _6179_/Q _6013_/C _6207_/Q VGND VGND VPWR VPWR _6014_/A
+ sky130_fd_sc_hd__a41o_1
.ends

