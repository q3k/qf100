magic
tech sky130A
magscale 1 2
timestamp 1647564177
<< obsli1 >>
rect 1104 2159 98808 37553
<< obsm1 >>
rect 474 1708 99530 37584
<< metal2 >>
rect 478 39200 534 40000
rect 1398 39200 1454 40000
rect 2318 39200 2374 40000
rect 3238 39200 3294 40000
rect 4250 39200 4306 40000
rect 5170 39200 5226 40000
rect 6090 39200 6146 40000
rect 7010 39200 7066 40000
rect 8022 39200 8078 40000
rect 8942 39200 8998 40000
rect 9862 39200 9918 40000
rect 10782 39200 10838 40000
rect 11794 39200 11850 40000
rect 12714 39200 12770 40000
rect 13634 39200 13690 40000
rect 14554 39200 14610 40000
rect 15566 39200 15622 40000
rect 16486 39200 16542 40000
rect 17406 39200 17462 40000
rect 18326 39200 18382 40000
rect 19338 39200 19394 40000
rect 20258 39200 20314 40000
rect 21178 39200 21234 40000
rect 22098 39200 22154 40000
rect 23110 39200 23166 40000
rect 24030 39200 24086 40000
rect 24950 39200 25006 40000
rect 25870 39200 25926 40000
rect 26882 39200 26938 40000
rect 27802 39200 27858 40000
rect 28722 39200 28778 40000
rect 29642 39200 29698 40000
rect 30654 39200 30710 40000
rect 31574 39200 31630 40000
rect 32494 39200 32550 40000
rect 33414 39200 33470 40000
rect 34426 39200 34482 40000
rect 35346 39200 35402 40000
rect 36266 39200 36322 40000
rect 37186 39200 37242 40000
rect 38198 39200 38254 40000
rect 39118 39200 39174 40000
rect 40038 39200 40094 40000
rect 40958 39200 41014 40000
rect 41970 39200 42026 40000
rect 42890 39200 42946 40000
rect 43810 39200 43866 40000
rect 44730 39200 44786 40000
rect 45742 39200 45798 40000
rect 46662 39200 46718 40000
rect 47582 39200 47638 40000
rect 48502 39200 48558 40000
rect 49514 39200 49570 40000
rect 50434 39200 50490 40000
rect 51354 39200 51410 40000
rect 52366 39200 52422 40000
rect 53286 39200 53342 40000
rect 54206 39200 54262 40000
rect 55126 39200 55182 40000
rect 56138 39200 56194 40000
rect 57058 39200 57114 40000
rect 57978 39200 58034 40000
rect 58898 39200 58954 40000
rect 59910 39200 59966 40000
rect 60830 39200 60886 40000
rect 61750 39200 61806 40000
rect 62670 39200 62726 40000
rect 63682 39200 63738 40000
rect 64602 39200 64658 40000
rect 65522 39200 65578 40000
rect 66442 39200 66498 40000
rect 67454 39200 67510 40000
rect 68374 39200 68430 40000
rect 69294 39200 69350 40000
rect 70214 39200 70270 40000
rect 71226 39200 71282 40000
rect 72146 39200 72202 40000
rect 73066 39200 73122 40000
rect 73986 39200 74042 40000
rect 74998 39200 75054 40000
rect 75918 39200 75974 40000
rect 76838 39200 76894 40000
rect 77758 39200 77814 40000
rect 78770 39200 78826 40000
rect 79690 39200 79746 40000
rect 80610 39200 80666 40000
rect 81530 39200 81586 40000
rect 82542 39200 82598 40000
rect 83462 39200 83518 40000
rect 84382 39200 84438 40000
rect 85302 39200 85358 40000
rect 86314 39200 86370 40000
rect 87234 39200 87290 40000
rect 88154 39200 88210 40000
rect 89074 39200 89130 40000
rect 90086 39200 90142 40000
rect 91006 39200 91062 40000
rect 91926 39200 91982 40000
rect 92846 39200 92902 40000
rect 93858 39200 93914 40000
rect 94778 39200 94834 40000
rect 95698 39200 95754 40000
rect 96618 39200 96674 40000
rect 97630 39200 97686 40000
rect 98550 39200 98606 40000
rect 99470 39200 99526 40000
rect 478 0 534 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 3238 0 3294 800
rect 4158 0 4214 800
rect 5078 0 5134 800
rect 5998 0 6054 800
rect 7010 0 7066 800
rect 7930 0 7986 800
rect 8850 0 8906 800
rect 9770 0 9826 800
rect 10690 0 10746 800
rect 11610 0 11666 800
rect 12622 0 12678 800
rect 13542 0 13598 800
rect 14462 0 14518 800
rect 15382 0 15438 800
rect 16302 0 16358 800
rect 17222 0 17278 800
rect 18234 0 18290 800
rect 19154 0 19210 800
rect 20074 0 20130 800
rect 20994 0 21050 800
rect 21914 0 21970 800
rect 22834 0 22890 800
rect 23754 0 23810 800
rect 24766 0 24822 800
rect 25686 0 25742 800
rect 26606 0 26662 800
rect 27526 0 27582 800
rect 28446 0 28502 800
rect 29366 0 29422 800
rect 30378 0 30434 800
rect 31298 0 31354 800
rect 32218 0 32274 800
rect 33138 0 33194 800
rect 34058 0 34114 800
rect 34978 0 35034 800
rect 35990 0 36046 800
rect 36910 0 36966 800
rect 37830 0 37886 800
rect 38750 0 38806 800
rect 39670 0 39726 800
rect 40590 0 40646 800
rect 41510 0 41566 800
rect 42522 0 42578 800
rect 43442 0 43498 800
rect 44362 0 44418 800
rect 45282 0 45338 800
rect 46202 0 46258 800
rect 47122 0 47178 800
rect 48134 0 48190 800
rect 49054 0 49110 800
rect 49974 0 50030 800
rect 50894 0 50950 800
rect 51814 0 51870 800
rect 52734 0 52790 800
rect 53746 0 53802 800
rect 54666 0 54722 800
rect 55586 0 55642 800
rect 56506 0 56562 800
rect 57426 0 57482 800
rect 58346 0 58402 800
rect 59358 0 59414 800
rect 60278 0 60334 800
rect 61198 0 61254 800
rect 62118 0 62174 800
rect 63038 0 63094 800
rect 63958 0 64014 800
rect 64878 0 64934 800
rect 65890 0 65946 800
rect 66810 0 66866 800
rect 67730 0 67786 800
rect 68650 0 68706 800
rect 69570 0 69626 800
rect 70490 0 70546 800
rect 71502 0 71558 800
rect 72422 0 72478 800
rect 73342 0 73398 800
rect 74262 0 74318 800
rect 75182 0 75238 800
rect 76102 0 76158 800
rect 77114 0 77170 800
rect 78034 0 78090 800
rect 78954 0 79010 800
rect 79874 0 79930 800
rect 80794 0 80850 800
rect 81714 0 81770 800
rect 82634 0 82690 800
rect 83646 0 83702 800
rect 84566 0 84622 800
rect 85486 0 85542 800
rect 86406 0 86462 800
rect 87326 0 87382 800
rect 88246 0 88302 800
rect 89258 0 89314 800
rect 90178 0 90234 800
rect 91098 0 91154 800
rect 92018 0 92074 800
rect 92938 0 92994 800
rect 93858 0 93914 800
rect 94870 0 94926 800
rect 95790 0 95846 800
rect 96710 0 96766 800
rect 97630 0 97686 800
rect 98550 0 98606 800
rect 99470 0 99526 800
<< obsm2 >>
rect 18 39144 422 39250
rect 590 39144 1342 39250
rect 1510 39144 2262 39250
rect 2430 39144 3182 39250
rect 3350 39144 4194 39250
rect 4362 39144 5114 39250
rect 5282 39144 6034 39250
rect 6202 39144 6954 39250
rect 7122 39144 7966 39250
rect 8134 39144 8886 39250
rect 9054 39144 9806 39250
rect 9974 39144 10726 39250
rect 10894 39144 11738 39250
rect 11906 39144 12658 39250
rect 12826 39144 13578 39250
rect 13746 39144 14498 39250
rect 14666 39144 15510 39250
rect 15678 39144 16430 39250
rect 16598 39144 17350 39250
rect 17518 39144 18270 39250
rect 18438 39144 19282 39250
rect 19450 39144 20202 39250
rect 20370 39144 21122 39250
rect 21290 39144 22042 39250
rect 22210 39144 23054 39250
rect 23222 39144 23974 39250
rect 24142 39144 24894 39250
rect 25062 39144 25814 39250
rect 25982 39144 26826 39250
rect 26994 39144 27746 39250
rect 27914 39144 28666 39250
rect 28834 39144 29586 39250
rect 29754 39144 30598 39250
rect 30766 39144 31518 39250
rect 31686 39144 32438 39250
rect 32606 39144 33358 39250
rect 33526 39144 34370 39250
rect 34538 39144 35290 39250
rect 35458 39144 36210 39250
rect 36378 39144 37130 39250
rect 37298 39144 38142 39250
rect 38310 39144 39062 39250
rect 39230 39144 39982 39250
rect 40150 39144 40902 39250
rect 41070 39144 41914 39250
rect 42082 39144 42834 39250
rect 43002 39144 43754 39250
rect 43922 39144 44674 39250
rect 44842 39144 45686 39250
rect 45854 39144 46606 39250
rect 46774 39144 47526 39250
rect 47694 39144 48446 39250
rect 48614 39144 49458 39250
rect 49626 39144 50378 39250
rect 50546 39144 51298 39250
rect 51466 39144 52310 39250
rect 52478 39144 53230 39250
rect 53398 39144 54150 39250
rect 54318 39144 55070 39250
rect 55238 39144 56082 39250
rect 56250 39144 57002 39250
rect 57170 39144 57922 39250
rect 58090 39144 58842 39250
rect 59010 39144 59854 39250
rect 60022 39144 60774 39250
rect 60942 39144 61694 39250
rect 61862 39144 62614 39250
rect 62782 39144 63626 39250
rect 63794 39144 64546 39250
rect 64714 39144 65466 39250
rect 65634 39144 66386 39250
rect 66554 39144 67398 39250
rect 67566 39144 68318 39250
rect 68486 39144 69238 39250
rect 69406 39144 70158 39250
rect 70326 39144 71170 39250
rect 71338 39144 72090 39250
rect 72258 39144 73010 39250
rect 73178 39144 73930 39250
rect 74098 39144 74942 39250
rect 75110 39144 75862 39250
rect 76030 39144 76782 39250
rect 76950 39144 77702 39250
rect 77870 39144 78714 39250
rect 78882 39144 79634 39250
rect 79802 39144 80554 39250
rect 80722 39144 81474 39250
rect 81642 39144 82486 39250
rect 82654 39144 83406 39250
rect 83574 39144 84326 39250
rect 84494 39144 85246 39250
rect 85414 39144 86258 39250
rect 86426 39144 87178 39250
rect 87346 39144 88098 39250
rect 88266 39144 89018 39250
rect 89186 39144 90030 39250
rect 90198 39144 90950 39250
rect 91118 39144 91870 39250
rect 92038 39144 92790 39250
rect 92958 39144 93802 39250
rect 93970 39144 94722 39250
rect 94890 39144 95642 39250
rect 95810 39144 96562 39250
rect 96730 39144 97574 39250
rect 97742 39144 98494 39250
rect 98662 39144 99414 39250
rect 18 856 99524 39144
rect 18 734 422 856
rect 590 734 1342 856
rect 1510 734 2262 856
rect 2430 734 3182 856
rect 3350 734 4102 856
rect 4270 734 5022 856
rect 5190 734 5942 856
rect 6110 734 6954 856
rect 7122 734 7874 856
rect 8042 734 8794 856
rect 8962 734 9714 856
rect 9882 734 10634 856
rect 10802 734 11554 856
rect 11722 734 12566 856
rect 12734 734 13486 856
rect 13654 734 14406 856
rect 14574 734 15326 856
rect 15494 734 16246 856
rect 16414 734 17166 856
rect 17334 734 18178 856
rect 18346 734 19098 856
rect 19266 734 20018 856
rect 20186 734 20938 856
rect 21106 734 21858 856
rect 22026 734 22778 856
rect 22946 734 23698 856
rect 23866 734 24710 856
rect 24878 734 25630 856
rect 25798 734 26550 856
rect 26718 734 27470 856
rect 27638 734 28390 856
rect 28558 734 29310 856
rect 29478 734 30322 856
rect 30490 734 31242 856
rect 31410 734 32162 856
rect 32330 734 33082 856
rect 33250 734 34002 856
rect 34170 734 34922 856
rect 35090 734 35934 856
rect 36102 734 36854 856
rect 37022 734 37774 856
rect 37942 734 38694 856
rect 38862 734 39614 856
rect 39782 734 40534 856
rect 40702 734 41454 856
rect 41622 734 42466 856
rect 42634 734 43386 856
rect 43554 734 44306 856
rect 44474 734 45226 856
rect 45394 734 46146 856
rect 46314 734 47066 856
rect 47234 734 48078 856
rect 48246 734 48998 856
rect 49166 734 49918 856
rect 50086 734 50838 856
rect 51006 734 51758 856
rect 51926 734 52678 856
rect 52846 734 53690 856
rect 53858 734 54610 856
rect 54778 734 55530 856
rect 55698 734 56450 856
rect 56618 734 57370 856
rect 57538 734 58290 856
rect 58458 734 59302 856
rect 59470 734 60222 856
rect 60390 734 61142 856
rect 61310 734 62062 856
rect 62230 734 62982 856
rect 63150 734 63902 856
rect 64070 734 64822 856
rect 64990 734 65834 856
rect 66002 734 66754 856
rect 66922 734 67674 856
rect 67842 734 68594 856
rect 68762 734 69514 856
rect 69682 734 70434 856
rect 70602 734 71446 856
rect 71614 734 72366 856
rect 72534 734 73286 856
rect 73454 734 74206 856
rect 74374 734 75126 856
rect 75294 734 76046 856
rect 76214 734 77058 856
rect 77226 734 77978 856
rect 78146 734 78898 856
rect 79066 734 79818 856
rect 79986 734 80738 856
rect 80906 734 81658 856
rect 81826 734 82578 856
rect 82746 734 83590 856
rect 83758 734 84510 856
rect 84678 734 85430 856
rect 85598 734 86350 856
rect 86518 734 87270 856
rect 87438 734 88190 856
rect 88358 734 89202 856
rect 89370 734 90122 856
rect 90290 734 91042 856
rect 91210 734 91962 856
rect 92130 734 92882 856
rect 93050 734 93802 856
rect 93970 734 94814 856
rect 94982 734 95734 856
rect 95902 734 96654 856
rect 96822 734 97574 856
rect 97742 734 98494 856
rect 98662 734 99414 856
<< metal3 >>
rect 0 20000 800 20120
<< obsm3 >>
rect 13 20200 96688 37569
rect 880 19920 96688 20200
rect 13 1667 96688 19920
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
rect 50288 2128 50608 37584
rect 65648 2128 65968 37584
rect 81008 2128 81328 37584
rect 96368 2128 96688 37584
<< obsm4 >>
rect 9627 8331 19488 13293
rect 19968 8331 34848 13293
rect 35328 8331 38581 13293
<< labels >>
rlabel metal2 s 478 0 534 800 6 CLK
port 1 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 RST_N
port 2 nsew signal input
rlabel metal4 s 19568 2128 19888 37584 6 VGND
port 3 nsew ground input
rlabel metal4 s 50288 2128 50608 37584 6 VGND
port 3 nsew ground input
rlabel metal4 s 81008 2128 81328 37584 6 VGND
port 3 nsew ground input
rlabel metal4 s 4208 2128 4528 37584 6 VPWR
port 4 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 VPWR
port 4 nsew power input
rlabel metal4 s 65648 2128 65968 37584 6 VPWR
port 4 nsew power input
rlabel metal4 s 96368 2128 96688 37584 6 VPWR
port 4 nsew power input
rlabel metal2 s 7930 0 7986 800 6 cpu_ack_o
port 5 nsew signal output
rlabel metal2 s 10690 0 10746 800 6 cpu_adr_i[0]
port 6 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 cpu_adr_i[10]
port 7 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 cpu_adr_i[11]
port 8 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 cpu_adr_i[12]
port 9 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 cpu_adr_i[13]
port 10 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 cpu_adr_i[14]
port 11 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 cpu_adr_i[15]
port 12 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 cpu_adr_i[16]
port 13 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 cpu_adr_i[17]
port 14 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 cpu_adr_i[18]
port 15 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 cpu_adr_i[19]
port 16 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 cpu_adr_i[1]
port 17 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 cpu_adr_i[20]
port 18 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 cpu_adr_i[21]
port 19 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 cpu_adr_i[22]
port 20 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 cpu_adr_i[23]
port 21 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 cpu_adr_i[24]
port 22 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 cpu_adr_i[25]
port 23 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 cpu_adr_i[26]
port 24 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 cpu_adr_i[27]
port 25 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 cpu_adr_i[28]
port 26 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 cpu_adr_i[29]
port 27 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 cpu_adr_i[2]
port 28 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 cpu_adr_i[30]
port 29 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 cpu_adr_i[31]
port 30 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 cpu_adr_i[3]
port 31 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 cpu_adr_i[4]
port 32 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 cpu_adr_i[5]
port 33 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 cpu_adr_i[6]
port 34 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 cpu_adr_i[7]
port 35 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 cpu_adr_i[8]
port 36 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 cpu_adr_i[9]
port 37 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 cpu_cyc_i
port 38 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 cpu_dat_i[0]
port 39 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 cpu_dat_i[10]
port 40 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 cpu_dat_i[11]
port 41 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 cpu_dat_i[12]
port 42 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 cpu_dat_i[13]
port 43 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 cpu_dat_i[14]
port 44 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 cpu_dat_i[15]
port 45 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 cpu_dat_i[16]
port 46 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 cpu_dat_i[17]
port 47 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 cpu_dat_i[18]
port 48 nsew signal input
rlabel metal2 s 76102 0 76158 800 6 cpu_dat_i[19]
port 49 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 cpu_dat_i[1]
port 50 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 cpu_dat_i[20]
port 51 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 cpu_dat_i[21]
port 52 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 cpu_dat_i[22]
port 53 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 cpu_dat_i[23]
port 54 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 cpu_dat_i[24]
port 55 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 cpu_dat_i[25]
port 56 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 cpu_dat_i[26]
port 57 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 cpu_dat_i[27]
port 58 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 cpu_dat_i[28]
port 59 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 cpu_dat_i[29]
port 60 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 cpu_dat_i[2]
port 61 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 cpu_dat_i[30]
port 62 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 cpu_dat_i[31]
port 63 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 cpu_dat_i[3]
port 64 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 cpu_dat_i[4]
port 65 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 cpu_dat_i[5]
port 66 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 cpu_dat_i[6]
port 67 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 cpu_dat_i[7]
port 68 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 cpu_dat_i[8]
port 69 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 cpu_dat_i[9]
port 70 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 cpu_dat_o[0]
port 71 nsew signal output
rlabel metal2 s 60278 0 60334 800 6 cpu_dat_o[10]
port 72 nsew signal output
rlabel metal2 s 62118 0 62174 800 6 cpu_dat_o[11]
port 73 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 cpu_dat_o[12]
port 74 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 cpu_dat_o[13]
port 75 nsew signal output
rlabel metal2 s 67730 0 67786 800 6 cpu_dat_o[14]
port 76 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 cpu_dat_o[15]
port 77 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 cpu_dat_o[16]
port 78 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 cpu_dat_o[17]
port 79 nsew signal output
rlabel metal2 s 75182 0 75238 800 6 cpu_dat_o[18]
port 80 nsew signal output
rlabel metal2 s 77114 0 77170 800 6 cpu_dat_o[19]
port 81 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 cpu_dat_o[1]
port 82 nsew signal output
rlabel metal2 s 78954 0 79010 800 6 cpu_dat_o[20]
port 83 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 cpu_dat_o[21]
port 84 nsew signal output
rlabel metal2 s 82634 0 82690 800 6 cpu_dat_o[22]
port 85 nsew signal output
rlabel metal2 s 84566 0 84622 800 6 cpu_dat_o[23]
port 86 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 cpu_dat_o[24]
port 87 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 cpu_dat_o[25]
port 88 nsew signal output
rlabel metal2 s 90178 0 90234 800 6 cpu_dat_o[26]
port 89 nsew signal output
rlabel metal2 s 92018 0 92074 800 6 cpu_dat_o[27]
port 90 nsew signal output
rlabel metal2 s 93858 0 93914 800 6 cpu_dat_o[28]
port 91 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 cpu_dat_o[29]
port 92 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 cpu_dat_o[2]
port 93 nsew signal output
rlabel metal2 s 97630 0 97686 800 6 cpu_dat_o[30]
port 94 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 cpu_dat_o[31]
port 95 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 cpu_dat_o[3]
port 96 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 cpu_dat_o[4]
port 97 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 cpu_dat_o[5]
port 98 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 cpu_dat_o[6]
port 99 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 cpu_dat_o[7]
port 100 nsew signal output
rlabel metal2 s 56506 0 56562 800 6 cpu_dat_o[8]
port 101 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 cpu_dat_o[9]
port 102 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 cpu_err_o
port 103 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 cpu_rty_o
port 104 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 cpu_sel_i[0]
port 105 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 cpu_sel_i[1]
port 106 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 cpu_sel_i[2]
port 107 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 cpu_sel_i[3]
port 108 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 cpu_stb_i
port 109 nsew signal input
rlabel metal3 s 0 20000 800 20120 6 cpu_we_i
port 110 nsew signal input
rlabel metal2 s 6090 39200 6146 40000 6 spi_ack_i
port 111 nsew signal input
rlabel metal2 s 8942 39200 8998 40000 6 spi_adr_o[0]
port 112 nsew signal output
rlabel metal2 s 18326 39200 18382 40000 6 spi_adr_o[10]
port 113 nsew signal output
rlabel metal2 s 19338 39200 19394 40000 6 spi_adr_o[11]
port 114 nsew signal output
rlabel metal2 s 20258 39200 20314 40000 6 spi_adr_o[12]
port 115 nsew signal output
rlabel metal2 s 21178 39200 21234 40000 6 spi_adr_o[13]
port 116 nsew signal output
rlabel metal2 s 22098 39200 22154 40000 6 spi_adr_o[14]
port 117 nsew signal output
rlabel metal2 s 23110 39200 23166 40000 6 spi_adr_o[15]
port 118 nsew signal output
rlabel metal2 s 24030 39200 24086 40000 6 spi_adr_o[16]
port 119 nsew signal output
rlabel metal2 s 24950 39200 25006 40000 6 spi_adr_o[17]
port 120 nsew signal output
rlabel metal2 s 25870 39200 25926 40000 6 spi_adr_o[18]
port 121 nsew signal output
rlabel metal2 s 26882 39200 26938 40000 6 spi_adr_o[19]
port 122 nsew signal output
rlabel metal2 s 9862 39200 9918 40000 6 spi_adr_o[1]
port 123 nsew signal output
rlabel metal2 s 27802 39200 27858 40000 6 spi_adr_o[20]
port 124 nsew signal output
rlabel metal2 s 28722 39200 28778 40000 6 spi_adr_o[21]
port 125 nsew signal output
rlabel metal2 s 29642 39200 29698 40000 6 spi_adr_o[22]
port 126 nsew signal output
rlabel metal2 s 30654 39200 30710 40000 6 spi_adr_o[23]
port 127 nsew signal output
rlabel metal2 s 31574 39200 31630 40000 6 spi_adr_o[24]
port 128 nsew signal output
rlabel metal2 s 32494 39200 32550 40000 6 spi_adr_o[25]
port 129 nsew signal output
rlabel metal2 s 33414 39200 33470 40000 6 spi_adr_o[26]
port 130 nsew signal output
rlabel metal2 s 34426 39200 34482 40000 6 spi_adr_o[27]
port 131 nsew signal output
rlabel metal2 s 35346 39200 35402 40000 6 spi_adr_o[28]
port 132 nsew signal output
rlabel metal2 s 36266 39200 36322 40000 6 spi_adr_o[29]
port 133 nsew signal output
rlabel metal2 s 10782 39200 10838 40000 6 spi_adr_o[2]
port 134 nsew signal output
rlabel metal2 s 37186 39200 37242 40000 6 spi_adr_o[30]
port 135 nsew signal output
rlabel metal2 s 38198 39200 38254 40000 6 spi_adr_o[31]
port 136 nsew signal output
rlabel metal2 s 11794 39200 11850 40000 6 spi_adr_o[3]
port 137 nsew signal output
rlabel metal2 s 12714 39200 12770 40000 6 spi_adr_o[4]
port 138 nsew signal output
rlabel metal2 s 13634 39200 13690 40000 6 spi_adr_o[5]
port 139 nsew signal output
rlabel metal2 s 14554 39200 14610 40000 6 spi_adr_o[6]
port 140 nsew signal output
rlabel metal2 s 15566 39200 15622 40000 6 spi_adr_o[7]
port 141 nsew signal output
rlabel metal2 s 16486 39200 16542 40000 6 spi_adr_o[8]
port 142 nsew signal output
rlabel metal2 s 17406 39200 17462 40000 6 spi_adr_o[9]
port 143 nsew signal output
rlabel metal2 s 478 39200 534 40000 6 spi_cyc_o
port 144 nsew signal output
rlabel metal2 s 39118 39200 39174 40000 6 spi_dat_i[0]
port 145 nsew signal input
rlabel metal2 s 57978 39200 58034 40000 6 spi_dat_i[10]
port 146 nsew signal input
rlabel metal2 s 59910 39200 59966 40000 6 spi_dat_i[11]
port 147 nsew signal input
rlabel metal2 s 61750 39200 61806 40000 6 spi_dat_i[12]
port 148 nsew signal input
rlabel metal2 s 63682 39200 63738 40000 6 spi_dat_i[13]
port 149 nsew signal input
rlabel metal2 s 65522 39200 65578 40000 6 spi_dat_i[14]
port 150 nsew signal input
rlabel metal2 s 67454 39200 67510 40000 6 spi_dat_i[15]
port 151 nsew signal input
rlabel metal2 s 69294 39200 69350 40000 6 spi_dat_i[16]
port 152 nsew signal input
rlabel metal2 s 71226 39200 71282 40000 6 spi_dat_i[17]
port 153 nsew signal input
rlabel metal2 s 73066 39200 73122 40000 6 spi_dat_i[18]
port 154 nsew signal input
rlabel metal2 s 74998 39200 75054 40000 6 spi_dat_i[19]
port 155 nsew signal input
rlabel metal2 s 40958 39200 41014 40000 6 spi_dat_i[1]
port 156 nsew signal input
rlabel metal2 s 76838 39200 76894 40000 6 spi_dat_i[20]
port 157 nsew signal input
rlabel metal2 s 78770 39200 78826 40000 6 spi_dat_i[21]
port 158 nsew signal input
rlabel metal2 s 80610 39200 80666 40000 6 spi_dat_i[22]
port 159 nsew signal input
rlabel metal2 s 82542 39200 82598 40000 6 spi_dat_i[23]
port 160 nsew signal input
rlabel metal2 s 84382 39200 84438 40000 6 spi_dat_i[24]
port 161 nsew signal input
rlabel metal2 s 86314 39200 86370 40000 6 spi_dat_i[25]
port 162 nsew signal input
rlabel metal2 s 88154 39200 88210 40000 6 spi_dat_i[26]
port 163 nsew signal input
rlabel metal2 s 90086 39200 90142 40000 6 spi_dat_i[27]
port 164 nsew signal input
rlabel metal2 s 91926 39200 91982 40000 6 spi_dat_i[28]
port 165 nsew signal input
rlabel metal2 s 93858 39200 93914 40000 6 spi_dat_i[29]
port 166 nsew signal input
rlabel metal2 s 42890 39200 42946 40000 6 spi_dat_i[2]
port 167 nsew signal input
rlabel metal2 s 95698 39200 95754 40000 6 spi_dat_i[30]
port 168 nsew signal input
rlabel metal2 s 97630 39200 97686 40000 6 spi_dat_i[31]
port 169 nsew signal input
rlabel metal2 s 44730 39200 44786 40000 6 spi_dat_i[3]
port 170 nsew signal input
rlabel metal2 s 46662 39200 46718 40000 6 spi_dat_i[4]
port 171 nsew signal input
rlabel metal2 s 48502 39200 48558 40000 6 spi_dat_i[5]
port 172 nsew signal input
rlabel metal2 s 50434 39200 50490 40000 6 spi_dat_i[6]
port 173 nsew signal input
rlabel metal2 s 52366 39200 52422 40000 6 spi_dat_i[7]
port 174 nsew signal input
rlabel metal2 s 54206 39200 54262 40000 6 spi_dat_i[8]
port 175 nsew signal input
rlabel metal2 s 56138 39200 56194 40000 6 spi_dat_i[9]
port 176 nsew signal input
rlabel metal2 s 40038 39200 40094 40000 6 spi_dat_o[0]
port 177 nsew signal output
rlabel metal2 s 58898 39200 58954 40000 6 spi_dat_o[10]
port 178 nsew signal output
rlabel metal2 s 60830 39200 60886 40000 6 spi_dat_o[11]
port 179 nsew signal output
rlabel metal2 s 62670 39200 62726 40000 6 spi_dat_o[12]
port 180 nsew signal output
rlabel metal2 s 64602 39200 64658 40000 6 spi_dat_o[13]
port 181 nsew signal output
rlabel metal2 s 66442 39200 66498 40000 6 spi_dat_o[14]
port 182 nsew signal output
rlabel metal2 s 68374 39200 68430 40000 6 spi_dat_o[15]
port 183 nsew signal output
rlabel metal2 s 70214 39200 70270 40000 6 spi_dat_o[16]
port 184 nsew signal output
rlabel metal2 s 72146 39200 72202 40000 6 spi_dat_o[17]
port 185 nsew signal output
rlabel metal2 s 73986 39200 74042 40000 6 spi_dat_o[18]
port 186 nsew signal output
rlabel metal2 s 75918 39200 75974 40000 6 spi_dat_o[19]
port 187 nsew signal output
rlabel metal2 s 41970 39200 42026 40000 6 spi_dat_o[1]
port 188 nsew signal output
rlabel metal2 s 77758 39200 77814 40000 6 spi_dat_o[20]
port 189 nsew signal output
rlabel metal2 s 79690 39200 79746 40000 6 spi_dat_o[21]
port 190 nsew signal output
rlabel metal2 s 81530 39200 81586 40000 6 spi_dat_o[22]
port 191 nsew signal output
rlabel metal2 s 83462 39200 83518 40000 6 spi_dat_o[23]
port 192 nsew signal output
rlabel metal2 s 85302 39200 85358 40000 6 spi_dat_o[24]
port 193 nsew signal output
rlabel metal2 s 87234 39200 87290 40000 6 spi_dat_o[25]
port 194 nsew signal output
rlabel metal2 s 89074 39200 89130 40000 6 spi_dat_o[26]
port 195 nsew signal output
rlabel metal2 s 91006 39200 91062 40000 6 spi_dat_o[27]
port 196 nsew signal output
rlabel metal2 s 92846 39200 92902 40000 6 spi_dat_o[28]
port 197 nsew signal output
rlabel metal2 s 94778 39200 94834 40000 6 spi_dat_o[29]
port 198 nsew signal output
rlabel metal2 s 43810 39200 43866 40000 6 spi_dat_o[2]
port 199 nsew signal output
rlabel metal2 s 96618 39200 96674 40000 6 spi_dat_o[30]
port 200 nsew signal output
rlabel metal2 s 98550 39200 98606 40000 6 spi_dat_o[31]
port 201 nsew signal output
rlabel metal2 s 45742 39200 45798 40000 6 spi_dat_o[3]
port 202 nsew signal output
rlabel metal2 s 47582 39200 47638 40000 6 spi_dat_o[4]
port 203 nsew signal output
rlabel metal2 s 49514 39200 49570 40000 6 spi_dat_o[5]
port 204 nsew signal output
rlabel metal2 s 51354 39200 51410 40000 6 spi_dat_o[6]
port 205 nsew signal output
rlabel metal2 s 53286 39200 53342 40000 6 spi_dat_o[7]
port 206 nsew signal output
rlabel metal2 s 55126 39200 55182 40000 6 spi_dat_o[8]
port 207 nsew signal output
rlabel metal2 s 57058 39200 57114 40000 6 spi_dat_o[9]
port 208 nsew signal output
rlabel metal2 s 7010 39200 7066 40000 6 spi_err_i
port 209 nsew signal input
rlabel metal2 s 8022 39200 8078 40000 6 spi_rty_i
port 210 nsew signal input
rlabel metal2 s 2318 39200 2374 40000 6 spi_sel_o[0]
port 211 nsew signal output
rlabel metal2 s 3238 39200 3294 40000 6 spi_sel_o[1]
port 212 nsew signal output
rlabel metal2 s 4250 39200 4306 40000 6 spi_sel_o[2]
port 213 nsew signal output
rlabel metal2 s 5170 39200 5226 40000 6 spi_sel_o[3]
port 214 nsew signal output
rlabel metal2 s 1398 39200 1454 40000 6 spi_stb_o
port 215 nsew signal output
rlabel metal2 s 99470 39200 99526 40000 6 spi_we_o
port 216 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 100000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8939158
string GDS_FILE /home/q3k/sky130/qf105/openlane/mkQF100Fabric/runs/mkQF100Fabric/results/finishing/mkQF100Fabric.magic.gds
string GDS_START 742466
<< end >>

