VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mkQF100FlashController
  CLASS BLOCK ;
  FOREIGN mkQF100FlashController ;
  ORIGIN 0.000 0.000 ;
  SIZE 617.125 BY 627.845 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END CLK
  PIN EN_serverA_request_put
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END EN_serverA_request_put
  PIN EN_serverA_response_get
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END EN_serverA_response_get
  PIN EN_serverB_request_put
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 4.120 617.125 4.720 ;
    END
  END EN_serverB_request_put
  PIN EN_serverB_response_get
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 12.960 617.125 13.560 ;
    END
  END EN_serverB_response_get
  PIN RDY_serverA_request_put
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END RDY_serverA_request_put
  PIN RDY_serverA_response_get
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END RDY_serverA_response_get
  PIN RDY_serverB_request_put
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 22.480 617.125 23.080 ;
    END
  END RDY_serverB_request_put
  PIN RDY_serverB_response_get
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 31.320 617.125 31.920 ;
    END
  END RDY_serverB_response_get
  PIN RST_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END RST_N
  PIN serverA_request_put[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END serverA_request_put[0]
  PIN serverA_request_put[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END serverA_request_put[10]
  PIN serverA_request_put[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END serverA_request_put[11]
  PIN serverA_request_put[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END serverA_request_put[12]
  PIN serverA_request_put[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END serverA_request_put[13]
  PIN serverA_request_put[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END serverA_request_put[14]
  PIN serverA_request_put[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END serverA_request_put[15]
  PIN serverA_request_put[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END serverA_request_put[16]
  PIN serverA_request_put[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END serverA_request_put[17]
  PIN serverA_request_put[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END serverA_request_put[18]
  PIN serverA_request_put[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END serverA_request_put[19]
  PIN serverA_request_put[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END serverA_request_put[1]
  PIN serverA_request_put[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 0.000 403.790 4.000 ;
    END
  END serverA_request_put[20]
  PIN serverA_request_put[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 0.000 421.730 4.000 ;
    END
  END serverA_request_put[21]
  PIN serverA_request_put[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END serverA_request_put[22]
  PIN serverA_request_put[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END serverA_request_put[23]
  PIN serverA_request_put[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 0.000 476.470 4.000 ;
    END
  END serverA_request_put[24]
  PIN serverA_request_put[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END serverA_request_put[25]
  PIN serverA_request_put[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.530 0.000 512.810 4.000 ;
    END
  END serverA_request_put[26]
  PIN serverA_request_put[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 0.000 530.750 4.000 ;
    END
  END serverA_request_put[27]
  PIN serverA_request_put[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.870 0.000 549.150 4.000 ;
    END
  END serverA_request_put[28]
  PIN serverA_request_put[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END serverA_request_put[29]
  PIN serverA_request_put[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END serverA_request_put[2]
  PIN serverA_request_put[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END serverA_request_put[30]
  PIN serverA_request_put[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 0.000 603.430 4.000 ;
    END
  END serverA_request_put[31]
  PIN serverA_request_put[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END serverA_request_put[3]
  PIN serverA_request_put[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END serverA_request_put[4]
  PIN serverA_request_put[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END serverA_request_put[5]
  PIN serverA_request_put[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END serverA_request_put[6]
  PIN serverA_request_put[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END serverA_request_put[7]
  PIN serverA_request_put[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END serverA_request_put[8]
  PIN serverA_request_put[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END serverA_request_put[9]
  PIN serverA_response_get[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END serverA_response_get[0]
  PIN serverA_response_get[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END serverA_response_get[10]
  PIN serverA_response_get[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END serverA_response_get[11]
  PIN serverA_response_get[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END serverA_response_get[12]
  PIN serverA_response_get[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END serverA_response_get[13]
  PIN serverA_response_get[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END serverA_response_get[14]
  PIN serverA_response_get[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END serverA_response_get[15]
  PIN serverA_response_get[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END serverA_response_get[16]
  PIN serverA_response_get[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END serverA_response_get[17]
  PIN serverA_response_get[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END serverA_response_get[18]
  PIN serverA_response_get[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 0.000 394.590 4.000 ;
    END
  END serverA_response_get[19]
  PIN serverA_response_get[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END serverA_response_get[1]
  PIN serverA_response_get[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END serverA_response_get[20]
  PIN serverA_response_get[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END serverA_response_get[21]
  PIN serverA_response_get[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END serverA_response_get[22]
  PIN serverA_response_get[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END serverA_response_get[23]
  PIN serverA_response_get[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 0.000 485.210 4.000 ;
    END
  END serverA_response_get[24]
  PIN serverA_response_get[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 0.000 503.610 4.000 ;
    END
  END serverA_response_get[25]
  PIN serverA_response_get[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 0.000 521.550 4.000 ;
    END
  END serverA_response_get[26]
  PIN serverA_response_get[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 0.000 539.950 4.000 ;
    END
  END serverA_response_get[27]
  PIN serverA_response_get[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END serverA_response_get[28]
  PIN serverA_response_get[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 0.000 576.290 4.000 ;
    END
  END serverA_response_get[29]
  PIN serverA_response_get[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END serverA_response_get[2]
  PIN serverA_response_get[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 0.000 594.230 4.000 ;
    END
  END serverA_response_get[30]
  PIN serverA_response_get[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 0.000 612.630 4.000 ;
    END
  END serverA_response_get[31]
  PIN serverA_response_get[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END serverA_response_get[3]
  PIN serverA_response_get[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END serverA_response_get[4]
  PIN serverA_response_get[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END serverA_response_get[5]
  PIN serverA_response_get[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END serverA_response_get[6]
  PIN serverA_response_get[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END serverA_response_get[7]
  PIN serverA_response_get[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END serverA_response_get[8]
  PIN serverA_response_get[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END serverA_response_get[9]
  PIN serverB_request_put[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 40.840 617.125 41.440 ;
    END
  END serverB_request_put[0]
  PIN serverB_request_put[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 225.120 617.125 225.720 ;
    END
  END serverB_request_put[10]
  PIN serverB_request_put[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 243.480 617.125 244.080 ;
    END
  END serverB_request_put[11]
  PIN serverB_request_put[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 262.520 617.125 263.120 ;
    END
  END serverB_request_put[12]
  PIN serverB_request_put[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 280.880 617.125 281.480 ;
    END
  END serverB_request_put[13]
  PIN serverB_request_put[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 299.240 617.125 299.840 ;
    END
  END serverB_request_put[14]
  PIN serverB_request_put[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 317.600 617.125 318.200 ;
    END
  END serverB_request_put[15]
  PIN serverB_request_put[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 335.960 617.125 336.560 ;
    END
  END serverB_request_put[16]
  PIN serverB_request_put[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 354.320 617.125 354.920 ;
    END
  END serverB_request_put[17]
  PIN serverB_request_put[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 372.680 617.125 373.280 ;
    END
  END serverB_request_put[18]
  PIN serverB_request_put[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 391.720 617.125 392.320 ;
    END
  END serverB_request_put[19]
  PIN serverB_request_put[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 59.200 617.125 59.800 ;
    END
  END serverB_request_put[1]
  PIN serverB_request_put[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 410.080 617.125 410.680 ;
    END
  END serverB_request_put[20]
  PIN serverB_request_put[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 428.440 617.125 429.040 ;
    END
  END serverB_request_put[21]
  PIN serverB_request_put[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 446.800 617.125 447.400 ;
    END
  END serverB_request_put[22]
  PIN serverB_request_put[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 465.160 617.125 465.760 ;
    END
  END serverB_request_put[23]
  PIN serverB_request_put[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 483.520 617.125 484.120 ;
    END
  END serverB_request_put[24]
  PIN serverB_request_put[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 501.880 617.125 502.480 ;
    END
  END serverB_request_put[25]
  PIN serverB_request_put[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 520.920 617.125 521.520 ;
    END
  END serverB_request_put[26]
  PIN serverB_request_put[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 539.280 617.125 539.880 ;
    END
  END serverB_request_put[27]
  PIN serverB_request_put[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 557.640 617.125 558.240 ;
    END
  END serverB_request_put[28]
  PIN serverB_request_put[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 576.000 617.125 576.600 ;
    END
  END serverB_request_put[29]
  PIN serverB_request_put[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 77.560 617.125 78.160 ;
    END
  END serverB_request_put[2]
  PIN serverB_request_put[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 594.360 617.125 594.960 ;
    END
  END serverB_request_put[30]
  PIN serverB_request_put[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 612.720 617.125 613.320 ;
    END
  END serverB_request_put[31]
  PIN serverB_request_put[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 95.920 617.125 96.520 ;
    END
  END serverB_request_put[3]
  PIN serverB_request_put[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 114.280 617.125 114.880 ;
    END
  END serverB_request_put[4]
  PIN serverB_request_put[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 133.320 617.125 133.920 ;
    END
  END serverB_request_put[5]
  PIN serverB_request_put[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 151.680 617.125 152.280 ;
    END
  END serverB_request_put[6]
  PIN serverB_request_put[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 170.040 617.125 170.640 ;
    END
  END serverB_request_put[7]
  PIN serverB_request_put[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 188.400 617.125 189.000 ;
    END
  END serverB_request_put[8]
  PIN serverB_request_put[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 206.760 617.125 207.360 ;
    END
  END serverB_request_put[9]
  PIN serverB_response_get[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 49.680 617.125 50.280 ;
    END
  END serverB_response_get[0]
  PIN serverB_response_get[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 234.640 617.125 235.240 ;
    END
  END serverB_response_get[10]
  PIN serverB_response_get[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 253.000 617.125 253.600 ;
    END
  END serverB_response_get[11]
  PIN serverB_response_get[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 271.360 617.125 271.960 ;
    END
  END serverB_response_get[12]
  PIN serverB_response_get[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 289.720 617.125 290.320 ;
    END
  END serverB_response_get[13]
  PIN serverB_response_get[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 308.080 617.125 308.680 ;
    END
  END serverB_response_get[14]
  PIN serverB_response_get[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 327.120 617.125 327.720 ;
    END
  END serverB_response_get[15]
  PIN serverB_response_get[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 345.480 617.125 346.080 ;
    END
  END serverB_response_get[16]
  PIN serverB_response_get[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 363.840 617.125 364.440 ;
    END
  END serverB_response_get[17]
  PIN serverB_response_get[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 382.200 617.125 382.800 ;
    END
  END serverB_response_get[18]
  PIN serverB_response_get[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 400.560 617.125 401.160 ;
    END
  END serverB_response_get[19]
  PIN serverB_response_get[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 68.720 617.125 69.320 ;
    END
  END serverB_response_get[1]
  PIN serverB_response_get[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 418.920 617.125 419.520 ;
    END
  END serverB_response_get[20]
  PIN serverB_response_get[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 437.280 617.125 437.880 ;
    END
  END serverB_response_get[21]
  PIN serverB_response_get[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 456.320 617.125 456.920 ;
    END
  END serverB_response_get[22]
  PIN serverB_response_get[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 474.680 617.125 475.280 ;
    END
  END serverB_response_get[23]
  PIN serverB_response_get[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 493.040 617.125 493.640 ;
    END
  END serverB_response_get[24]
  PIN serverB_response_get[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 511.400 617.125 512.000 ;
    END
  END serverB_response_get[25]
  PIN serverB_response_get[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 529.760 617.125 530.360 ;
    END
  END serverB_response_get[26]
  PIN serverB_response_get[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 548.120 617.125 548.720 ;
    END
  END serverB_response_get[27]
  PIN serverB_response_get[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 566.480 617.125 567.080 ;
    END
  END serverB_response_get[28]
  PIN serverB_response_get[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 585.520 617.125 586.120 ;
    END
  END serverB_response_get[29]
  PIN serverB_response_get[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 87.080 617.125 87.680 ;
    END
  END serverB_response_get[2]
  PIN serverB_response_get[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 603.880 617.125 604.480 ;
    END
  END serverB_response_get[30]
  PIN serverB_response_get[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 622.240 617.125 622.840 ;
    END
  END serverB_response_get[31]
  PIN serverB_response_get[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 105.440 617.125 106.040 ;
    END
  END serverB_response_get[3]
  PIN serverB_response_get[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 123.800 617.125 124.400 ;
    END
  END serverB_response_get[4]
  PIN serverB_response_get[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 142.160 617.125 142.760 ;
    END
  END serverB_response_get[5]
  PIN serverB_response_get[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 160.520 617.125 161.120 ;
    END
  END serverB_response_get[6]
  PIN serverB_response_get[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 178.880 617.125 179.480 ;
    END
  END serverB_response_get[7]
  PIN serverB_response_get[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 197.920 617.125 198.520 ;
    END
  END serverB_response_get[8]
  PIN serverB_response_get[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 613.125 216.280 617.125 216.880 ;
    END
  END serverB_response_get[9]
  PIN spi_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END spi_csb
  PIN spi_miso
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END spi_miso
  PIN spi_mosi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END spi_mosi
  PIN spi_mosi_oe
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 4.000 492.960 ;
    END
  END spi_mosi_oe
  PIN spi_sclk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END spi_sclk
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 614.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 614.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 614.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 614.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 614.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 614.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 614.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 614.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 611.340 614.805 ;
      LAYER met1 ;
        RECT 4.210 7.860 612.650 614.960 ;
      LAYER met2 ;
        RECT 4.240 4.280 612.620 622.725 ;
        RECT 4.790 4.000 12.690 4.280 ;
        RECT 13.530 4.000 21.890 4.280 ;
        RECT 22.730 4.000 31.090 4.280 ;
        RECT 31.930 4.000 39.830 4.280 ;
        RECT 40.670 4.000 49.030 4.280 ;
        RECT 49.870 4.000 58.230 4.280 ;
        RECT 59.070 4.000 67.430 4.280 ;
        RECT 68.270 4.000 76.170 4.280 ;
        RECT 77.010 4.000 85.370 4.280 ;
        RECT 86.210 4.000 94.570 4.280 ;
        RECT 95.410 4.000 103.770 4.280 ;
        RECT 104.610 4.000 112.510 4.280 ;
        RECT 113.350 4.000 121.710 4.280 ;
        RECT 122.550 4.000 130.910 4.280 ;
        RECT 131.750 4.000 140.110 4.280 ;
        RECT 140.950 4.000 148.850 4.280 ;
        RECT 149.690 4.000 158.050 4.280 ;
        RECT 158.890 4.000 167.250 4.280 ;
        RECT 168.090 4.000 175.990 4.280 ;
        RECT 176.830 4.000 185.190 4.280 ;
        RECT 186.030 4.000 194.390 4.280 ;
        RECT 195.230 4.000 203.590 4.280 ;
        RECT 204.430 4.000 212.330 4.280 ;
        RECT 213.170 4.000 221.530 4.280 ;
        RECT 222.370 4.000 230.730 4.280 ;
        RECT 231.570 4.000 239.930 4.280 ;
        RECT 240.770 4.000 248.670 4.280 ;
        RECT 249.510 4.000 257.870 4.280 ;
        RECT 258.710 4.000 267.070 4.280 ;
        RECT 267.910 4.000 276.270 4.280 ;
        RECT 277.110 4.000 285.010 4.280 ;
        RECT 285.850 4.000 294.210 4.280 ;
        RECT 295.050 4.000 303.410 4.280 ;
        RECT 304.250 4.000 312.610 4.280 ;
        RECT 313.450 4.000 321.350 4.280 ;
        RECT 322.190 4.000 330.550 4.280 ;
        RECT 331.390 4.000 339.750 4.280 ;
        RECT 340.590 4.000 348.490 4.280 ;
        RECT 349.330 4.000 357.690 4.280 ;
        RECT 358.530 4.000 366.890 4.280 ;
        RECT 367.730 4.000 376.090 4.280 ;
        RECT 376.930 4.000 384.830 4.280 ;
        RECT 385.670 4.000 394.030 4.280 ;
        RECT 394.870 4.000 403.230 4.280 ;
        RECT 404.070 4.000 412.430 4.280 ;
        RECT 413.270 4.000 421.170 4.280 ;
        RECT 422.010 4.000 430.370 4.280 ;
        RECT 431.210 4.000 439.570 4.280 ;
        RECT 440.410 4.000 448.770 4.280 ;
        RECT 449.610 4.000 457.510 4.280 ;
        RECT 458.350 4.000 466.710 4.280 ;
        RECT 467.550 4.000 475.910 4.280 ;
        RECT 476.750 4.000 484.650 4.280 ;
        RECT 485.490 4.000 493.850 4.280 ;
        RECT 494.690 4.000 503.050 4.280 ;
        RECT 503.890 4.000 512.250 4.280 ;
        RECT 513.090 4.000 520.990 4.280 ;
        RECT 521.830 4.000 530.190 4.280 ;
        RECT 531.030 4.000 539.390 4.280 ;
        RECT 540.230 4.000 548.590 4.280 ;
        RECT 549.430 4.000 557.330 4.280 ;
        RECT 558.170 4.000 566.530 4.280 ;
        RECT 567.370 4.000 575.730 4.280 ;
        RECT 576.570 4.000 584.930 4.280 ;
        RECT 585.770 4.000 593.670 4.280 ;
        RECT 594.510 4.000 602.870 4.280 ;
        RECT 603.710 4.000 612.070 4.280 ;
      LAYER met3 ;
        RECT 4.000 621.840 612.725 622.705 ;
        RECT 4.000 613.720 613.125 621.840 ;
        RECT 4.000 612.320 612.725 613.720 ;
        RECT 4.000 604.880 613.125 612.320 ;
        RECT 4.000 603.480 612.725 604.880 ;
        RECT 4.000 595.360 613.125 603.480 ;
        RECT 4.000 593.960 612.725 595.360 ;
        RECT 4.000 586.520 613.125 593.960 ;
        RECT 4.000 585.120 612.725 586.520 ;
        RECT 4.000 583.120 613.125 585.120 ;
        RECT 4.400 581.720 613.125 583.120 ;
        RECT 4.000 577.000 613.125 581.720 ;
        RECT 4.000 575.600 612.725 577.000 ;
        RECT 4.000 567.480 613.125 575.600 ;
        RECT 4.000 566.080 612.725 567.480 ;
        RECT 4.000 558.640 613.125 566.080 ;
        RECT 4.000 557.240 612.725 558.640 ;
        RECT 4.000 549.120 613.125 557.240 ;
        RECT 4.000 547.720 612.725 549.120 ;
        RECT 4.000 540.280 613.125 547.720 ;
        RECT 4.000 538.880 612.725 540.280 ;
        RECT 4.000 530.760 613.125 538.880 ;
        RECT 4.000 529.360 612.725 530.760 ;
        RECT 4.000 521.920 613.125 529.360 ;
        RECT 4.000 520.520 612.725 521.920 ;
        RECT 4.000 512.400 613.125 520.520 ;
        RECT 4.000 511.000 612.725 512.400 ;
        RECT 4.000 502.880 613.125 511.000 ;
        RECT 4.000 501.480 612.725 502.880 ;
        RECT 4.000 494.040 613.125 501.480 ;
        RECT 4.000 493.360 612.725 494.040 ;
        RECT 4.400 492.640 612.725 493.360 ;
        RECT 4.400 491.960 613.125 492.640 ;
        RECT 4.000 484.520 613.125 491.960 ;
        RECT 4.000 483.120 612.725 484.520 ;
        RECT 4.000 475.680 613.125 483.120 ;
        RECT 4.000 474.280 612.725 475.680 ;
        RECT 4.000 466.160 613.125 474.280 ;
        RECT 4.000 464.760 612.725 466.160 ;
        RECT 4.000 457.320 613.125 464.760 ;
        RECT 4.000 455.920 612.725 457.320 ;
        RECT 4.000 447.800 613.125 455.920 ;
        RECT 4.000 446.400 612.725 447.800 ;
        RECT 4.000 438.280 613.125 446.400 ;
        RECT 4.000 436.880 612.725 438.280 ;
        RECT 4.000 429.440 613.125 436.880 ;
        RECT 4.000 428.040 612.725 429.440 ;
        RECT 4.000 419.920 613.125 428.040 ;
        RECT 4.000 418.520 612.725 419.920 ;
        RECT 4.000 411.080 613.125 418.520 ;
        RECT 4.000 409.680 612.725 411.080 ;
        RECT 4.000 403.600 613.125 409.680 ;
        RECT 4.400 402.200 613.125 403.600 ;
        RECT 4.000 401.560 613.125 402.200 ;
        RECT 4.000 400.160 612.725 401.560 ;
        RECT 4.000 392.720 613.125 400.160 ;
        RECT 4.000 391.320 612.725 392.720 ;
        RECT 4.000 383.200 613.125 391.320 ;
        RECT 4.000 381.800 612.725 383.200 ;
        RECT 4.000 373.680 613.125 381.800 ;
        RECT 4.000 372.280 612.725 373.680 ;
        RECT 4.000 364.840 613.125 372.280 ;
        RECT 4.000 363.440 612.725 364.840 ;
        RECT 4.000 355.320 613.125 363.440 ;
        RECT 4.000 353.920 612.725 355.320 ;
        RECT 4.000 346.480 613.125 353.920 ;
        RECT 4.000 345.080 612.725 346.480 ;
        RECT 4.000 336.960 613.125 345.080 ;
        RECT 4.000 335.560 612.725 336.960 ;
        RECT 4.000 328.120 613.125 335.560 ;
        RECT 4.000 326.720 612.725 328.120 ;
        RECT 4.000 318.600 613.125 326.720 ;
        RECT 4.000 317.200 612.725 318.600 ;
        RECT 4.000 313.840 613.125 317.200 ;
        RECT 4.400 312.440 613.125 313.840 ;
        RECT 4.000 309.080 613.125 312.440 ;
        RECT 4.000 307.680 612.725 309.080 ;
        RECT 4.000 300.240 613.125 307.680 ;
        RECT 4.000 298.840 612.725 300.240 ;
        RECT 4.000 290.720 613.125 298.840 ;
        RECT 4.000 289.320 612.725 290.720 ;
        RECT 4.000 281.880 613.125 289.320 ;
        RECT 4.000 280.480 612.725 281.880 ;
        RECT 4.000 272.360 613.125 280.480 ;
        RECT 4.000 270.960 612.725 272.360 ;
        RECT 4.000 263.520 613.125 270.960 ;
        RECT 4.000 262.120 612.725 263.520 ;
        RECT 4.000 254.000 613.125 262.120 ;
        RECT 4.000 252.600 612.725 254.000 ;
        RECT 4.000 244.480 613.125 252.600 ;
        RECT 4.000 243.080 612.725 244.480 ;
        RECT 4.000 235.640 613.125 243.080 ;
        RECT 4.000 234.240 612.725 235.640 ;
        RECT 4.000 226.120 613.125 234.240 ;
        RECT 4.000 224.720 612.725 226.120 ;
        RECT 4.000 224.080 613.125 224.720 ;
        RECT 4.400 222.680 613.125 224.080 ;
        RECT 4.000 217.280 613.125 222.680 ;
        RECT 4.000 215.880 612.725 217.280 ;
        RECT 4.000 207.760 613.125 215.880 ;
        RECT 4.000 206.360 612.725 207.760 ;
        RECT 4.000 198.920 613.125 206.360 ;
        RECT 4.000 197.520 612.725 198.920 ;
        RECT 4.000 189.400 613.125 197.520 ;
        RECT 4.000 188.000 612.725 189.400 ;
        RECT 4.000 179.880 613.125 188.000 ;
        RECT 4.000 178.480 612.725 179.880 ;
        RECT 4.000 171.040 613.125 178.480 ;
        RECT 4.000 169.640 612.725 171.040 ;
        RECT 4.000 161.520 613.125 169.640 ;
        RECT 4.000 160.120 612.725 161.520 ;
        RECT 4.000 152.680 613.125 160.120 ;
        RECT 4.000 151.280 612.725 152.680 ;
        RECT 4.000 143.160 613.125 151.280 ;
        RECT 4.000 141.760 612.725 143.160 ;
        RECT 4.000 134.320 613.125 141.760 ;
        RECT 4.400 132.920 612.725 134.320 ;
        RECT 4.000 124.800 613.125 132.920 ;
        RECT 4.000 123.400 612.725 124.800 ;
        RECT 4.000 115.280 613.125 123.400 ;
        RECT 4.000 113.880 612.725 115.280 ;
        RECT 4.000 106.440 613.125 113.880 ;
        RECT 4.000 105.040 612.725 106.440 ;
        RECT 4.000 96.920 613.125 105.040 ;
        RECT 4.000 95.520 612.725 96.920 ;
        RECT 4.000 88.080 613.125 95.520 ;
        RECT 4.000 86.680 612.725 88.080 ;
        RECT 4.000 78.560 613.125 86.680 ;
        RECT 4.000 77.160 612.725 78.560 ;
        RECT 4.000 69.720 613.125 77.160 ;
        RECT 4.000 68.320 612.725 69.720 ;
        RECT 4.000 60.200 613.125 68.320 ;
        RECT 4.000 58.800 612.725 60.200 ;
        RECT 4.000 50.680 613.125 58.800 ;
        RECT 4.000 49.280 612.725 50.680 ;
        RECT 4.000 45.240 613.125 49.280 ;
        RECT 4.400 43.840 613.125 45.240 ;
        RECT 4.000 41.840 613.125 43.840 ;
        RECT 4.000 40.440 612.725 41.840 ;
        RECT 4.000 32.320 613.125 40.440 ;
        RECT 4.000 30.920 612.725 32.320 ;
        RECT 4.000 23.480 613.125 30.920 ;
        RECT 4.000 22.080 612.725 23.480 ;
        RECT 4.000 13.960 613.125 22.080 ;
        RECT 4.000 12.560 612.725 13.960 ;
        RECT 4.000 5.120 613.125 12.560 ;
        RECT 4.000 4.255 612.725 5.120 ;
      LAYER met4 ;
        RECT 19.615 19.215 20.640 594.145 ;
        RECT 23.040 19.215 97.440 594.145 ;
        RECT 99.840 19.215 174.240 594.145 ;
        RECT 176.640 19.215 251.040 594.145 ;
        RECT 253.440 19.215 327.840 594.145 ;
        RECT 330.240 19.215 404.640 594.145 ;
        RECT 407.040 19.215 481.440 594.145 ;
        RECT 483.840 19.215 558.240 594.145 ;
        RECT 560.640 19.215 604.145 594.145 ;
  END
END mkQF100FlashController
END LIBRARY

