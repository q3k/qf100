magic
tech sky130A
magscale 1 2
timestamp 1647601538
<< obsli1 >>
rect 1104 2159 166980 168113
<< obsm1 >>
rect 1026 1300 167058 168144
<< metal2 >>
rect 1030 169475 1086 170275
rect 3146 169475 3202 170275
rect 5354 169475 5410 170275
rect 7562 169475 7618 170275
rect 9678 169475 9734 170275
rect 11886 169475 11942 170275
rect 14094 169475 14150 170275
rect 16302 169475 16358 170275
rect 18418 169475 18474 170275
rect 20626 169475 20682 170275
rect 22834 169475 22890 170275
rect 25042 169475 25098 170275
rect 27158 169475 27214 170275
rect 29366 169475 29422 170275
rect 31574 169475 31630 170275
rect 33782 169475 33838 170275
rect 35898 169475 35954 170275
rect 38106 169475 38162 170275
rect 40314 169475 40370 170275
rect 42522 169475 42578 170275
rect 44638 169475 44694 170275
rect 46846 169475 46902 170275
rect 49054 169475 49110 170275
rect 51262 169475 51318 170275
rect 53378 169475 53434 170275
rect 55586 169475 55642 170275
rect 57794 169475 57850 170275
rect 59910 169475 59966 170275
rect 62118 169475 62174 170275
rect 64326 169475 64382 170275
rect 66534 169475 66590 170275
rect 68650 169475 68706 170275
rect 70858 169475 70914 170275
rect 73066 169475 73122 170275
rect 75274 169475 75330 170275
rect 77390 169475 77446 170275
rect 79598 169475 79654 170275
rect 81806 169475 81862 170275
rect 84014 169475 84070 170275
rect 86130 169475 86186 170275
rect 88338 169475 88394 170275
rect 90546 169475 90602 170275
rect 92754 169475 92810 170275
rect 94870 169475 94926 170275
rect 97078 169475 97134 170275
rect 99286 169475 99342 170275
rect 101494 169475 101550 170275
rect 103610 169475 103666 170275
rect 105818 169475 105874 170275
rect 108026 169475 108082 170275
rect 110234 169475 110290 170275
rect 112350 169475 112406 170275
rect 114558 169475 114614 170275
rect 116766 169475 116822 170275
rect 118882 169475 118938 170275
rect 121090 169475 121146 170275
rect 123298 169475 123354 170275
rect 125506 169475 125562 170275
rect 127622 169475 127678 170275
rect 129830 169475 129886 170275
rect 132038 169475 132094 170275
rect 134246 169475 134302 170275
rect 136362 169475 136418 170275
rect 138570 169475 138626 170275
rect 140778 169475 140834 170275
rect 142986 169475 143042 170275
rect 145102 169475 145158 170275
rect 147310 169475 147366 170275
rect 149518 169475 149574 170275
rect 151726 169475 151782 170275
rect 153842 169475 153898 170275
rect 156050 169475 156106 170275
rect 158258 169475 158314 170275
rect 160466 169475 160522 170275
rect 162582 169475 162638 170275
rect 164790 169475 164846 170275
rect 166998 169475 167054 170275
rect 9310 0 9366 800
rect 27986 0 28042 800
rect 46662 0 46718 800
rect 65338 0 65394 800
rect 84014 0 84070 800
rect 102690 0 102746 800
rect 121366 0 121422 800
rect 140042 0 140098 800
rect 158718 0 158774 800
<< obsm2 >>
rect 1142 169419 3090 169697
rect 3258 169419 5298 169697
rect 5466 169419 7506 169697
rect 7674 169419 9622 169697
rect 9790 169419 11830 169697
rect 11998 169419 14038 169697
rect 14206 169419 16246 169697
rect 16414 169419 18362 169697
rect 18530 169419 20570 169697
rect 20738 169419 22778 169697
rect 22946 169419 24986 169697
rect 25154 169419 27102 169697
rect 27270 169419 29310 169697
rect 29478 169419 31518 169697
rect 31686 169419 33726 169697
rect 33894 169419 35842 169697
rect 36010 169419 38050 169697
rect 38218 169419 40258 169697
rect 40426 169419 42466 169697
rect 42634 169419 44582 169697
rect 44750 169419 46790 169697
rect 46958 169419 48998 169697
rect 49166 169419 51206 169697
rect 51374 169419 53322 169697
rect 53490 169419 55530 169697
rect 55698 169419 57738 169697
rect 57906 169419 59854 169697
rect 60022 169419 62062 169697
rect 62230 169419 64270 169697
rect 64438 169419 66478 169697
rect 66646 169419 68594 169697
rect 68762 169419 70802 169697
rect 70970 169419 73010 169697
rect 73178 169419 75218 169697
rect 75386 169419 77334 169697
rect 77502 169419 79542 169697
rect 79710 169419 81750 169697
rect 81918 169419 83958 169697
rect 84126 169419 86074 169697
rect 86242 169419 88282 169697
rect 88450 169419 90490 169697
rect 90658 169419 92698 169697
rect 92866 169419 94814 169697
rect 94982 169419 97022 169697
rect 97190 169419 99230 169697
rect 99398 169419 101438 169697
rect 101606 169419 103554 169697
rect 103722 169419 105762 169697
rect 105930 169419 107970 169697
rect 108138 169419 110178 169697
rect 110346 169419 112294 169697
rect 112462 169419 114502 169697
rect 114670 169419 116710 169697
rect 116878 169419 118826 169697
rect 118994 169419 121034 169697
rect 121202 169419 123242 169697
rect 123410 169419 125450 169697
rect 125618 169419 127566 169697
rect 127734 169419 129774 169697
rect 129942 169419 131982 169697
rect 132150 169419 134190 169697
rect 134358 169419 136306 169697
rect 136474 169419 138514 169697
rect 138682 169419 140722 169697
rect 140890 169419 142930 169697
rect 143098 169419 145046 169697
rect 145214 169419 147254 169697
rect 147422 169419 149462 169697
rect 149630 169419 151670 169697
rect 151838 169419 153786 169697
rect 153954 169419 155994 169697
rect 156162 169419 158202 169697
rect 158370 169419 160410 169697
rect 160578 169419 162526 169697
rect 162694 169419 164734 169697
rect 164902 169419 166942 169697
rect 1032 856 167052 169419
rect 1032 575 9254 856
rect 9422 575 27930 856
rect 28098 575 46606 856
rect 46774 575 65282 856
rect 65450 575 83958 856
rect 84126 575 102634 856
rect 102802 575 121310 856
rect 121478 575 139986 856
rect 140154 575 158662 856
rect 158830 575 167052 856
<< metal3 >>
rect 0 169600 800 169720
rect 167331 169464 168131 169584
rect 0 168376 800 168496
rect 167331 167968 168131 168088
rect 0 167152 800 167272
rect 167331 166608 168131 166728
rect 0 165928 800 166048
rect 167331 165112 168131 165232
rect 0 164704 800 164824
rect 0 163480 800 163600
rect 167331 163616 168131 163736
rect 0 162256 800 162376
rect 167331 162256 168131 162376
rect 0 161032 800 161152
rect 167331 160760 168131 160880
rect 0 159944 800 160064
rect 167331 159400 168131 159520
rect 0 158720 800 158840
rect 167331 157904 168131 158024
rect 0 157496 800 157616
rect 0 156272 800 156392
rect 167331 156408 168131 156528
rect 0 155048 800 155168
rect 167331 155048 168131 155168
rect 0 153824 800 153944
rect 167331 153552 168131 153672
rect 0 152600 800 152720
rect 167331 152192 168131 152312
rect 0 151376 800 151496
rect 167331 150696 168131 150816
rect 0 150288 800 150408
rect 0 149064 800 149184
rect 167331 149200 168131 149320
rect 0 147840 800 147960
rect 167331 147840 168131 147960
rect 0 146616 800 146736
rect 167331 146344 168131 146464
rect 0 145392 800 145512
rect 167331 144984 168131 145104
rect 0 144168 800 144288
rect 167331 143488 168131 143608
rect 0 142944 800 143064
rect 167331 141992 168131 142112
rect 0 141720 800 141840
rect 0 140632 800 140752
rect 167331 140632 168131 140752
rect 0 139408 800 139528
rect 167331 139136 168131 139256
rect 0 138184 800 138304
rect 167331 137640 168131 137760
rect 0 136960 800 137080
rect 167331 136280 168131 136400
rect 0 135736 800 135856
rect 167331 134784 168131 134904
rect 0 134512 800 134632
rect 0 133288 800 133408
rect 167331 133424 168131 133544
rect 0 132064 800 132184
rect 167331 131928 168131 132048
rect 0 130840 800 130960
rect 167331 130432 168131 130552
rect 0 129752 800 129872
rect 167331 129072 168131 129192
rect 0 128528 800 128648
rect 167331 127576 168131 127696
rect 0 127304 800 127424
rect 0 126080 800 126200
rect 167331 126216 168131 126336
rect 0 124856 800 124976
rect 167331 124720 168131 124840
rect 0 123632 800 123752
rect 167331 123224 168131 123344
rect 0 122408 800 122528
rect 167331 121864 168131 121984
rect 0 121184 800 121304
rect 167331 120368 168131 120488
rect 0 120096 800 120216
rect 0 118872 800 118992
rect 167331 119008 168131 119128
rect 0 117648 800 117768
rect 167331 117512 168131 117632
rect 0 116424 800 116544
rect 167331 116016 168131 116136
rect 0 115200 800 115320
rect 167331 114656 168131 114776
rect 0 113976 800 114096
rect 167331 113160 168131 113280
rect 0 112752 800 112872
rect 0 111528 800 111648
rect 167331 111664 168131 111784
rect 0 110440 800 110560
rect 167331 110304 168131 110424
rect 0 109216 800 109336
rect 167331 108808 168131 108928
rect 0 107992 800 108112
rect 167331 107448 168131 107568
rect 0 106768 800 106888
rect 167331 105952 168131 106072
rect 0 105544 800 105664
rect 0 104320 800 104440
rect 167331 104456 168131 104576
rect 0 103096 800 103216
rect 167331 103096 168131 103216
rect 0 101872 800 101992
rect 167331 101600 168131 101720
rect 0 100648 800 100768
rect 167331 100240 168131 100360
rect 0 99560 800 99680
rect 167331 98744 168131 98864
rect 0 98336 800 98456
rect 0 97112 800 97232
rect 167331 97248 168131 97368
rect 0 95888 800 96008
rect 167331 95888 168131 96008
rect 0 94664 800 94784
rect 167331 94392 168131 94512
rect 0 93440 800 93560
rect 167331 93032 168131 93152
rect 0 92216 800 92336
rect 167331 91536 168131 91656
rect 0 90992 800 91112
rect 0 89904 800 90024
rect 167331 90040 168131 90160
rect 0 88680 800 88800
rect 167331 88680 168131 88800
rect 0 87456 800 87576
rect 167331 87184 168131 87304
rect 0 86232 800 86352
rect 167331 85824 168131 85944
rect 0 85008 800 85128
rect 167331 84328 168131 84448
rect 0 83784 800 83904
rect 167331 82832 168131 82952
rect 0 82560 800 82680
rect 0 81336 800 81456
rect 167331 81472 168131 81592
rect 0 80248 800 80368
rect 167331 79976 168131 80096
rect 0 79024 800 79144
rect 167331 78480 168131 78600
rect 0 77800 800 77920
rect 167331 77120 168131 77240
rect 0 76576 800 76696
rect 167331 75624 168131 75744
rect 0 75352 800 75472
rect 0 74128 800 74248
rect 167331 74264 168131 74384
rect 0 72904 800 73024
rect 167331 72768 168131 72888
rect 0 71680 800 71800
rect 167331 71272 168131 71392
rect 0 70592 800 70712
rect 167331 69912 168131 70032
rect 0 69368 800 69488
rect 167331 68416 168131 68536
rect 0 68144 800 68264
rect 0 66920 800 67040
rect 167331 67056 168131 67176
rect 0 65696 800 65816
rect 167331 65560 168131 65680
rect 0 64472 800 64592
rect 167331 64064 168131 64184
rect 0 63248 800 63368
rect 167331 62704 168131 62824
rect 0 62024 800 62144
rect 167331 61208 168131 61328
rect 0 60800 800 60920
rect 0 59712 800 59832
rect 167331 59848 168131 59968
rect 0 58488 800 58608
rect 167331 58352 168131 58472
rect 0 57264 800 57384
rect 167331 56856 168131 56976
rect 0 56040 800 56160
rect 167331 55496 168131 55616
rect 0 54816 800 54936
rect 167331 54000 168131 54120
rect 0 53592 800 53712
rect 0 52368 800 52488
rect 167331 52504 168131 52624
rect 0 51144 800 51264
rect 167331 51144 168131 51264
rect 0 50056 800 50176
rect 167331 49648 168131 49768
rect 0 48832 800 48952
rect 167331 48288 168131 48408
rect 0 47608 800 47728
rect 167331 46792 168131 46912
rect 0 46384 800 46504
rect 0 45160 800 45280
rect 167331 45296 168131 45416
rect 0 43936 800 44056
rect 167331 43936 168131 44056
rect 0 42712 800 42832
rect 167331 42440 168131 42560
rect 0 41488 800 41608
rect 167331 41080 168131 41200
rect 0 40400 800 40520
rect 167331 39584 168131 39704
rect 0 39176 800 39296
rect 0 37952 800 38072
rect 167331 38088 168131 38208
rect 0 36728 800 36848
rect 167331 36728 168131 36848
rect 0 35504 800 35624
rect 167331 35232 168131 35352
rect 0 34280 800 34400
rect 167331 33872 168131 33992
rect 0 33056 800 33176
rect 167331 32376 168131 32496
rect 0 31832 800 31952
rect 167331 30880 168131 31000
rect 0 30608 800 30728
rect 0 29520 800 29640
rect 167331 29520 168131 29640
rect 0 28296 800 28416
rect 167331 28024 168131 28144
rect 0 27072 800 27192
rect 167331 26528 168131 26648
rect 0 25848 800 25968
rect 167331 25168 168131 25288
rect 0 24624 800 24744
rect 167331 23672 168131 23792
rect 0 23400 800 23520
rect 0 22176 800 22296
rect 167331 22312 168131 22432
rect 0 20952 800 21072
rect 167331 20816 168131 20936
rect 0 19864 800 19984
rect 167331 19320 168131 19440
rect 0 18640 800 18760
rect 167331 17960 168131 18080
rect 0 17416 800 17536
rect 167331 16464 168131 16584
rect 0 16192 800 16312
rect 0 14968 800 15088
rect 167331 15104 168131 15224
rect 0 13744 800 13864
rect 167331 13608 168131 13728
rect 0 12520 800 12640
rect 167331 12112 168131 12232
rect 0 11296 800 11416
rect 167331 10752 168131 10872
rect 0 10208 800 10328
rect 167331 9256 168131 9376
rect 0 8984 800 9104
rect 0 7760 800 7880
rect 167331 7896 168131 8016
rect 0 6536 800 6656
rect 167331 6400 168131 6520
rect 0 5312 800 5432
rect 167331 4904 168131 5024
rect 0 4088 800 4208
rect 167331 3544 168131 3664
rect 0 2864 800 2984
rect 167331 2048 168131 2168
rect 0 1640 800 1760
rect 0 552 800 672
rect 167331 688 168131 808
<< obsm3 >>
rect 880 169664 167331 169693
rect 880 169520 167251 169664
rect 800 169384 167251 169520
rect 800 168576 167331 169384
rect 880 168296 167331 168576
rect 800 168168 167331 168296
rect 800 167888 167251 168168
rect 800 167352 167331 167888
rect 880 167072 167331 167352
rect 800 166808 167331 167072
rect 800 166528 167251 166808
rect 800 166128 167331 166528
rect 880 165848 167331 166128
rect 800 165312 167331 165848
rect 800 165032 167251 165312
rect 800 164904 167331 165032
rect 880 164624 167331 164904
rect 800 163816 167331 164624
rect 800 163680 167251 163816
rect 880 163536 167251 163680
rect 880 163400 167331 163536
rect 800 162456 167331 163400
rect 880 162176 167251 162456
rect 800 161232 167331 162176
rect 880 160960 167331 161232
rect 880 160952 167251 160960
rect 800 160680 167251 160952
rect 800 160144 167331 160680
rect 880 159864 167331 160144
rect 800 159600 167331 159864
rect 800 159320 167251 159600
rect 800 158920 167331 159320
rect 880 158640 167331 158920
rect 800 158104 167331 158640
rect 800 157824 167251 158104
rect 800 157696 167331 157824
rect 880 157416 167331 157696
rect 800 156608 167331 157416
rect 800 156472 167251 156608
rect 880 156328 167251 156472
rect 880 156192 167331 156328
rect 800 155248 167331 156192
rect 880 154968 167251 155248
rect 800 154024 167331 154968
rect 880 153752 167331 154024
rect 880 153744 167251 153752
rect 800 153472 167251 153744
rect 800 152800 167331 153472
rect 880 152520 167331 152800
rect 800 152392 167331 152520
rect 800 152112 167251 152392
rect 800 151576 167331 152112
rect 880 151296 167331 151576
rect 800 150896 167331 151296
rect 800 150616 167251 150896
rect 800 150488 167331 150616
rect 880 150208 167331 150488
rect 800 149400 167331 150208
rect 800 149264 167251 149400
rect 880 149120 167251 149264
rect 880 148984 167331 149120
rect 800 148040 167331 148984
rect 880 147760 167251 148040
rect 800 146816 167331 147760
rect 880 146544 167331 146816
rect 880 146536 167251 146544
rect 800 146264 167251 146536
rect 800 145592 167331 146264
rect 880 145312 167331 145592
rect 800 145184 167331 145312
rect 800 144904 167251 145184
rect 800 144368 167331 144904
rect 880 144088 167331 144368
rect 800 143688 167331 144088
rect 800 143408 167251 143688
rect 800 143144 167331 143408
rect 880 142864 167331 143144
rect 800 142192 167331 142864
rect 800 141920 167251 142192
rect 880 141912 167251 141920
rect 880 141640 167331 141912
rect 800 140832 167331 141640
rect 880 140552 167251 140832
rect 800 139608 167331 140552
rect 880 139336 167331 139608
rect 880 139328 167251 139336
rect 800 139056 167251 139328
rect 800 138384 167331 139056
rect 880 138104 167331 138384
rect 800 137840 167331 138104
rect 800 137560 167251 137840
rect 800 137160 167331 137560
rect 880 136880 167331 137160
rect 800 136480 167331 136880
rect 800 136200 167251 136480
rect 800 135936 167331 136200
rect 880 135656 167331 135936
rect 800 134984 167331 135656
rect 800 134712 167251 134984
rect 880 134704 167251 134712
rect 880 134432 167331 134704
rect 800 133624 167331 134432
rect 800 133488 167251 133624
rect 880 133344 167251 133488
rect 880 133208 167331 133344
rect 800 132264 167331 133208
rect 880 132128 167331 132264
rect 880 131984 167251 132128
rect 800 131848 167251 131984
rect 800 131040 167331 131848
rect 880 130760 167331 131040
rect 800 130632 167331 130760
rect 800 130352 167251 130632
rect 800 129952 167331 130352
rect 880 129672 167331 129952
rect 800 129272 167331 129672
rect 800 128992 167251 129272
rect 800 128728 167331 128992
rect 880 128448 167331 128728
rect 800 127776 167331 128448
rect 800 127504 167251 127776
rect 880 127496 167251 127504
rect 880 127224 167331 127496
rect 800 126416 167331 127224
rect 800 126280 167251 126416
rect 880 126136 167251 126280
rect 880 126000 167331 126136
rect 800 125056 167331 126000
rect 880 124920 167331 125056
rect 880 124776 167251 124920
rect 800 124640 167251 124776
rect 800 123832 167331 124640
rect 880 123552 167331 123832
rect 800 123424 167331 123552
rect 800 123144 167251 123424
rect 800 122608 167331 123144
rect 880 122328 167331 122608
rect 800 122064 167331 122328
rect 800 121784 167251 122064
rect 800 121384 167331 121784
rect 880 121104 167331 121384
rect 800 120568 167331 121104
rect 800 120296 167251 120568
rect 880 120288 167251 120296
rect 880 120016 167331 120288
rect 800 119208 167331 120016
rect 800 119072 167251 119208
rect 880 118928 167251 119072
rect 880 118792 167331 118928
rect 800 117848 167331 118792
rect 880 117712 167331 117848
rect 880 117568 167251 117712
rect 800 117432 167251 117568
rect 800 116624 167331 117432
rect 880 116344 167331 116624
rect 800 116216 167331 116344
rect 800 115936 167251 116216
rect 800 115400 167331 115936
rect 880 115120 167331 115400
rect 800 114856 167331 115120
rect 800 114576 167251 114856
rect 800 114176 167331 114576
rect 880 113896 167331 114176
rect 800 113360 167331 113896
rect 800 113080 167251 113360
rect 800 112952 167331 113080
rect 880 112672 167331 112952
rect 800 111864 167331 112672
rect 800 111728 167251 111864
rect 880 111584 167251 111728
rect 880 111448 167331 111584
rect 800 110640 167331 111448
rect 880 110504 167331 110640
rect 880 110360 167251 110504
rect 800 110224 167251 110360
rect 800 109416 167331 110224
rect 880 109136 167331 109416
rect 800 109008 167331 109136
rect 800 108728 167251 109008
rect 800 108192 167331 108728
rect 880 107912 167331 108192
rect 800 107648 167331 107912
rect 800 107368 167251 107648
rect 800 106968 167331 107368
rect 880 106688 167331 106968
rect 800 106152 167331 106688
rect 800 105872 167251 106152
rect 800 105744 167331 105872
rect 880 105464 167331 105744
rect 800 104656 167331 105464
rect 800 104520 167251 104656
rect 880 104376 167251 104520
rect 880 104240 167331 104376
rect 800 103296 167331 104240
rect 880 103016 167251 103296
rect 800 102072 167331 103016
rect 880 101800 167331 102072
rect 880 101792 167251 101800
rect 800 101520 167251 101792
rect 800 100848 167331 101520
rect 880 100568 167331 100848
rect 800 100440 167331 100568
rect 800 100160 167251 100440
rect 800 99760 167331 100160
rect 880 99480 167331 99760
rect 800 98944 167331 99480
rect 800 98664 167251 98944
rect 800 98536 167331 98664
rect 880 98256 167331 98536
rect 800 97448 167331 98256
rect 800 97312 167251 97448
rect 880 97168 167251 97312
rect 880 97032 167331 97168
rect 800 96088 167331 97032
rect 880 95808 167251 96088
rect 800 94864 167331 95808
rect 880 94592 167331 94864
rect 880 94584 167251 94592
rect 800 94312 167251 94584
rect 800 93640 167331 94312
rect 880 93360 167331 93640
rect 800 93232 167331 93360
rect 800 92952 167251 93232
rect 800 92416 167331 92952
rect 880 92136 167331 92416
rect 800 91736 167331 92136
rect 800 91456 167251 91736
rect 800 91192 167331 91456
rect 880 90912 167331 91192
rect 800 90240 167331 90912
rect 800 90104 167251 90240
rect 880 89960 167251 90104
rect 880 89824 167331 89960
rect 800 88880 167331 89824
rect 880 88600 167251 88880
rect 800 87656 167331 88600
rect 880 87384 167331 87656
rect 880 87376 167251 87384
rect 800 87104 167251 87376
rect 800 86432 167331 87104
rect 880 86152 167331 86432
rect 800 86024 167331 86152
rect 800 85744 167251 86024
rect 800 85208 167331 85744
rect 880 84928 167331 85208
rect 800 84528 167331 84928
rect 800 84248 167251 84528
rect 800 83984 167331 84248
rect 880 83704 167331 83984
rect 800 83032 167331 83704
rect 800 82760 167251 83032
rect 880 82752 167251 82760
rect 880 82480 167331 82752
rect 800 81672 167331 82480
rect 800 81536 167251 81672
rect 880 81392 167251 81536
rect 880 81256 167331 81392
rect 800 80448 167331 81256
rect 880 80176 167331 80448
rect 880 80168 167251 80176
rect 800 79896 167251 80168
rect 800 79224 167331 79896
rect 880 78944 167331 79224
rect 800 78680 167331 78944
rect 800 78400 167251 78680
rect 800 78000 167331 78400
rect 880 77720 167331 78000
rect 800 77320 167331 77720
rect 800 77040 167251 77320
rect 800 76776 167331 77040
rect 880 76496 167331 76776
rect 800 75824 167331 76496
rect 800 75552 167251 75824
rect 880 75544 167251 75552
rect 880 75272 167331 75544
rect 800 74464 167331 75272
rect 800 74328 167251 74464
rect 880 74184 167251 74328
rect 880 74048 167331 74184
rect 800 73104 167331 74048
rect 880 72968 167331 73104
rect 880 72824 167251 72968
rect 800 72688 167251 72824
rect 800 71880 167331 72688
rect 880 71600 167331 71880
rect 800 71472 167331 71600
rect 800 71192 167251 71472
rect 800 70792 167331 71192
rect 880 70512 167331 70792
rect 800 70112 167331 70512
rect 800 69832 167251 70112
rect 800 69568 167331 69832
rect 880 69288 167331 69568
rect 800 68616 167331 69288
rect 800 68344 167251 68616
rect 880 68336 167251 68344
rect 880 68064 167331 68336
rect 800 67256 167331 68064
rect 800 67120 167251 67256
rect 880 66976 167251 67120
rect 880 66840 167331 66976
rect 800 65896 167331 66840
rect 880 65760 167331 65896
rect 880 65616 167251 65760
rect 800 65480 167251 65616
rect 800 64672 167331 65480
rect 880 64392 167331 64672
rect 800 64264 167331 64392
rect 800 63984 167251 64264
rect 800 63448 167331 63984
rect 880 63168 167331 63448
rect 800 62904 167331 63168
rect 800 62624 167251 62904
rect 800 62224 167331 62624
rect 880 61944 167331 62224
rect 800 61408 167331 61944
rect 800 61128 167251 61408
rect 800 61000 167331 61128
rect 880 60720 167331 61000
rect 800 60048 167331 60720
rect 800 59912 167251 60048
rect 880 59768 167251 59912
rect 880 59632 167331 59768
rect 800 58688 167331 59632
rect 880 58552 167331 58688
rect 880 58408 167251 58552
rect 800 58272 167251 58408
rect 800 57464 167331 58272
rect 880 57184 167331 57464
rect 800 57056 167331 57184
rect 800 56776 167251 57056
rect 800 56240 167331 56776
rect 880 55960 167331 56240
rect 800 55696 167331 55960
rect 800 55416 167251 55696
rect 800 55016 167331 55416
rect 880 54736 167331 55016
rect 800 54200 167331 54736
rect 800 53920 167251 54200
rect 800 53792 167331 53920
rect 880 53512 167331 53792
rect 800 52704 167331 53512
rect 800 52568 167251 52704
rect 880 52424 167251 52568
rect 880 52288 167331 52424
rect 800 51344 167331 52288
rect 880 51064 167251 51344
rect 800 50256 167331 51064
rect 880 49976 167331 50256
rect 800 49848 167331 49976
rect 800 49568 167251 49848
rect 800 49032 167331 49568
rect 880 48752 167331 49032
rect 800 48488 167331 48752
rect 800 48208 167251 48488
rect 800 47808 167331 48208
rect 880 47528 167331 47808
rect 800 46992 167331 47528
rect 800 46712 167251 46992
rect 800 46584 167331 46712
rect 880 46304 167331 46584
rect 800 45496 167331 46304
rect 800 45360 167251 45496
rect 880 45216 167251 45360
rect 880 45080 167331 45216
rect 800 44136 167331 45080
rect 880 43856 167251 44136
rect 800 42912 167331 43856
rect 880 42640 167331 42912
rect 880 42632 167251 42640
rect 800 42360 167251 42632
rect 800 41688 167331 42360
rect 880 41408 167331 41688
rect 800 41280 167331 41408
rect 800 41000 167251 41280
rect 800 40600 167331 41000
rect 880 40320 167331 40600
rect 800 39784 167331 40320
rect 800 39504 167251 39784
rect 800 39376 167331 39504
rect 880 39096 167331 39376
rect 800 38288 167331 39096
rect 800 38152 167251 38288
rect 880 38008 167251 38152
rect 880 37872 167331 38008
rect 800 36928 167331 37872
rect 880 36648 167251 36928
rect 800 35704 167331 36648
rect 880 35432 167331 35704
rect 880 35424 167251 35432
rect 800 35152 167251 35424
rect 800 34480 167331 35152
rect 880 34200 167331 34480
rect 800 34072 167331 34200
rect 800 33792 167251 34072
rect 800 33256 167331 33792
rect 880 32976 167331 33256
rect 800 32576 167331 32976
rect 800 32296 167251 32576
rect 800 32032 167331 32296
rect 880 31752 167331 32032
rect 800 31080 167331 31752
rect 800 30808 167251 31080
rect 880 30800 167251 30808
rect 880 30528 167331 30800
rect 800 29720 167331 30528
rect 880 29440 167251 29720
rect 800 28496 167331 29440
rect 880 28224 167331 28496
rect 880 28216 167251 28224
rect 800 27944 167251 28216
rect 800 27272 167331 27944
rect 880 26992 167331 27272
rect 800 26728 167331 26992
rect 800 26448 167251 26728
rect 800 26048 167331 26448
rect 880 25768 167331 26048
rect 800 25368 167331 25768
rect 800 25088 167251 25368
rect 800 24824 167331 25088
rect 880 24544 167331 24824
rect 800 23872 167331 24544
rect 800 23600 167251 23872
rect 880 23592 167251 23600
rect 880 23320 167331 23592
rect 800 22512 167331 23320
rect 800 22376 167251 22512
rect 880 22232 167251 22376
rect 880 22096 167331 22232
rect 800 21152 167331 22096
rect 880 21016 167331 21152
rect 880 20872 167251 21016
rect 800 20736 167251 20872
rect 800 20064 167331 20736
rect 880 19784 167331 20064
rect 800 19520 167331 19784
rect 800 19240 167251 19520
rect 800 18840 167331 19240
rect 880 18560 167331 18840
rect 800 18160 167331 18560
rect 800 17880 167251 18160
rect 800 17616 167331 17880
rect 880 17336 167331 17616
rect 800 16664 167331 17336
rect 800 16392 167251 16664
rect 880 16384 167251 16392
rect 880 16112 167331 16384
rect 800 15304 167331 16112
rect 800 15168 167251 15304
rect 880 15024 167251 15168
rect 880 14888 167331 15024
rect 800 13944 167331 14888
rect 880 13808 167331 13944
rect 880 13664 167251 13808
rect 800 13528 167251 13664
rect 800 12720 167331 13528
rect 880 12440 167331 12720
rect 800 12312 167331 12440
rect 800 12032 167251 12312
rect 800 11496 167331 12032
rect 880 11216 167331 11496
rect 800 10952 167331 11216
rect 800 10672 167251 10952
rect 800 10408 167331 10672
rect 880 10128 167331 10408
rect 800 9456 167331 10128
rect 800 9184 167251 9456
rect 880 9176 167251 9184
rect 880 8904 167331 9176
rect 800 8096 167331 8904
rect 800 7960 167251 8096
rect 880 7816 167251 7960
rect 880 7680 167331 7816
rect 800 6736 167331 7680
rect 880 6600 167331 6736
rect 880 6456 167251 6600
rect 800 6320 167251 6456
rect 800 5512 167331 6320
rect 880 5232 167331 5512
rect 800 5104 167331 5232
rect 800 4824 167251 5104
rect 800 4288 167331 4824
rect 880 4008 167331 4288
rect 800 3744 167331 4008
rect 800 3464 167251 3744
rect 800 3064 167331 3464
rect 880 2784 167331 3064
rect 800 2248 167331 2784
rect 800 1968 167251 2248
rect 800 1840 167331 1968
rect 880 1560 167331 1840
rect 800 888 167331 1560
rect 800 752 167251 888
rect 880 608 167251 752
rect 880 579 167331 608
<< metal4 >>
rect 4208 2128 4528 168144
rect 19568 2128 19888 168144
rect 34928 2128 35248 168144
rect 50288 2128 50608 168144
rect 65648 2128 65968 168144
rect 81008 2128 81328 168144
rect 96368 2128 96688 168144
rect 111728 2128 112048 168144
rect 127088 2128 127408 168144
rect 142448 2128 142768 168144
rect 157808 2128 158128 168144
<< obsm4 >>
rect 1899 3979 4128 159629
rect 4608 3979 19488 159629
rect 19968 3979 34848 159629
rect 35328 3979 50208 159629
rect 50688 3979 65568 159629
rect 66048 3979 80928 159629
rect 81408 3979 96288 159629
rect 96768 3979 111648 159629
rect 112128 3979 127008 159629
rect 127488 3979 142368 159629
rect 142848 3979 157728 159629
rect 158208 3979 165541 159629
<< labels >>
rlabel metal3 s 167331 153552 168131 153672 6 CLK
port 1 nsew signal input
rlabel metal3 s 0 552 800 672 6 EN_dmem_client_request_get
port 2 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 EN_dmem_client_response_put
port 3 nsew signal input
rlabel metal2 s 1030 169475 1086 170275 6 EN_imem_client_request_get
port 4 nsew signal input
rlabel metal2 s 3146 169475 3202 170275 6 EN_imem_client_response_put
port 5 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 RDY_dmem_client_request_get
port 6 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 RDY_dmem_client_response_put
port 7 nsew signal output
rlabel metal2 s 5354 169475 5410 170275 6 RDY_imem_client_request_get
port 8 nsew signal output
rlabel metal2 s 7562 169475 7618 170275 6 RDY_imem_client_response_put
port 9 nsew signal output
rlabel metal2 s 149518 169475 149574 170275 6 RDY_readPC
port 10 nsew signal output
rlabel metal2 s 9310 0 9366 800 6 RST_N
port 11 nsew signal input
rlabel metal4 s 19568 2128 19888 168144 6 VGND
port 12 nsew ground input
rlabel metal4 s 50288 2128 50608 168144 6 VGND
port 12 nsew ground input
rlabel metal4 s 81008 2128 81328 168144 6 VGND
port 12 nsew ground input
rlabel metal4 s 111728 2128 112048 168144 6 VGND
port 12 nsew ground input
rlabel metal4 s 142448 2128 142768 168144 6 VGND
port 12 nsew ground input
rlabel metal4 s 4208 2128 4528 168144 6 VPWR
port 13 nsew power input
rlabel metal4 s 34928 2128 35248 168144 6 VPWR
port 13 nsew power input
rlabel metal4 s 65648 2128 65968 168144 6 VPWR
port 13 nsew power input
rlabel metal4 s 96368 2128 96688 168144 6 VPWR
port 13 nsew power input
rlabel metal4 s 127088 2128 127408 168144 6 VPWR
port 13 nsew power input
rlabel metal4 s 157808 2128 158128 168144 6 VPWR
port 13 nsew power input
rlabel metal3 s 0 5312 800 5432 6 dmem_client_request_get[0]
port 14 nsew signal output
rlabel metal3 s 0 29520 800 29640 6 dmem_client_request_get[10]
port 15 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 dmem_client_request_get[11]
port 16 nsew signal output
rlabel metal3 s 0 34280 800 34400 6 dmem_client_request_get[12]
port 17 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 dmem_client_request_get[13]
port 18 nsew signal output
rlabel metal3 s 0 39176 800 39296 6 dmem_client_request_get[14]
port 19 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 dmem_client_request_get[15]
port 20 nsew signal output
rlabel metal3 s 0 43936 800 44056 6 dmem_client_request_get[16]
port 21 nsew signal output
rlabel metal3 s 0 46384 800 46504 6 dmem_client_request_get[17]
port 22 nsew signal output
rlabel metal3 s 0 48832 800 48952 6 dmem_client_request_get[18]
port 23 nsew signal output
rlabel metal3 s 0 51144 800 51264 6 dmem_client_request_get[19]
port 24 nsew signal output
rlabel metal3 s 0 7760 800 7880 6 dmem_client_request_get[1]
port 25 nsew signal output
rlabel metal3 s 0 53592 800 53712 6 dmem_client_request_get[20]
port 26 nsew signal output
rlabel metal3 s 0 56040 800 56160 6 dmem_client_request_get[21]
port 27 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 dmem_client_request_get[22]
port 28 nsew signal output
rlabel metal3 s 0 60800 800 60920 6 dmem_client_request_get[23]
port 29 nsew signal output
rlabel metal3 s 0 63248 800 63368 6 dmem_client_request_get[24]
port 30 nsew signal output
rlabel metal3 s 0 65696 800 65816 6 dmem_client_request_get[25]
port 31 nsew signal output
rlabel metal3 s 0 68144 800 68264 6 dmem_client_request_get[26]
port 32 nsew signal output
rlabel metal3 s 0 70592 800 70712 6 dmem_client_request_get[27]
port 33 nsew signal output
rlabel metal3 s 0 72904 800 73024 6 dmem_client_request_get[28]
port 34 nsew signal output
rlabel metal3 s 0 75352 800 75472 6 dmem_client_request_get[29]
port 35 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 dmem_client_request_get[2]
port 36 nsew signal output
rlabel metal3 s 0 77800 800 77920 6 dmem_client_request_get[30]
port 37 nsew signal output
rlabel metal3 s 0 80248 800 80368 6 dmem_client_request_get[31]
port 38 nsew signal output
rlabel metal3 s 0 82560 800 82680 6 dmem_client_request_get[32]
port 39 nsew signal output
rlabel metal3 s 0 83784 800 83904 6 dmem_client_request_get[33]
port 40 nsew signal output
rlabel metal3 s 0 85008 800 85128 6 dmem_client_request_get[34]
port 41 nsew signal output
rlabel metal3 s 0 86232 800 86352 6 dmem_client_request_get[35]
port 42 nsew signal output
rlabel metal3 s 0 87456 800 87576 6 dmem_client_request_get[36]
port 43 nsew signal output
rlabel metal3 s 0 88680 800 88800 6 dmem_client_request_get[37]
port 44 nsew signal output
rlabel metal3 s 0 89904 800 90024 6 dmem_client_request_get[38]
port 45 nsew signal output
rlabel metal3 s 0 90992 800 91112 6 dmem_client_request_get[39]
port 46 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 dmem_client_request_get[3]
port 47 nsew signal output
rlabel metal3 s 0 92216 800 92336 6 dmem_client_request_get[40]
port 48 nsew signal output
rlabel metal3 s 0 93440 800 93560 6 dmem_client_request_get[41]
port 49 nsew signal output
rlabel metal3 s 0 94664 800 94784 6 dmem_client_request_get[42]
port 50 nsew signal output
rlabel metal3 s 0 95888 800 96008 6 dmem_client_request_get[43]
port 51 nsew signal output
rlabel metal3 s 0 97112 800 97232 6 dmem_client_request_get[44]
port 52 nsew signal output
rlabel metal3 s 0 98336 800 98456 6 dmem_client_request_get[45]
port 53 nsew signal output
rlabel metal3 s 0 99560 800 99680 6 dmem_client_request_get[46]
port 54 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 dmem_client_request_get[47]
port 55 nsew signal output
rlabel metal3 s 0 101872 800 101992 6 dmem_client_request_get[48]
port 56 nsew signal output
rlabel metal3 s 0 103096 800 103216 6 dmem_client_request_get[49]
port 57 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 dmem_client_request_get[4]
port 58 nsew signal output
rlabel metal3 s 0 104320 800 104440 6 dmem_client_request_get[50]
port 59 nsew signal output
rlabel metal3 s 0 105544 800 105664 6 dmem_client_request_get[51]
port 60 nsew signal output
rlabel metal3 s 0 106768 800 106888 6 dmem_client_request_get[52]
port 61 nsew signal output
rlabel metal3 s 0 107992 800 108112 6 dmem_client_request_get[53]
port 62 nsew signal output
rlabel metal3 s 0 109216 800 109336 6 dmem_client_request_get[54]
port 63 nsew signal output
rlabel metal3 s 0 110440 800 110560 6 dmem_client_request_get[55]
port 64 nsew signal output
rlabel metal3 s 0 111528 800 111648 6 dmem_client_request_get[56]
port 65 nsew signal output
rlabel metal3 s 0 112752 800 112872 6 dmem_client_request_get[57]
port 66 nsew signal output
rlabel metal3 s 0 113976 800 114096 6 dmem_client_request_get[58]
port 67 nsew signal output
rlabel metal3 s 0 115200 800 115320 6 dmem_client_request_get[59]
port 68 nsew signal output
rlabel metal3 s 0 17416 800 17536 6 dmem_client_request_get[5]
port 69 nsew signal output
rlabel metal3 s 0 116424 800 116544 6 dmem_client_request_get[60]
port 70 nsew signal output
rlabel metal3 s 0 117648 800 117768 6 dmem_client_request_get[61]
port 71 nsew signal output
rlabel metal3 s 0 118872 800 118992 6 dmem_client_request_get[62]
port 72 nsew signal output
rlabel metal3 s 0 120096 800 120216 6 dmem_client_request_get[63]
port 73 nsew signal output
rlabel metal3 s 0 121184 800 121304 6 dmem_client_request_get[64]
port 74 nsew signal output
rlabel metal3 s 0 122408 800 122528 6 dmem_client_request_get[65]
port 75 nsew signal output
rlabel metal3 s 0 123632 800 123752 6 dmem_client_request_get[66]
port 76 nsew signal output
rlabel metal3 s 0 124856 800 124976 6 dmem_client_request_get[67]
port 77 nsew signal output
rlabel metal3 s 0 126080 800 126200 6 dmem_client_request_get[68]
port 78 nsew signal output
rlabel metal3 s 0 127304 800 127424 6 dmem_client_request_get[69]
port 79 nsew signal output
rlabel metal3 s 0 19864 800 19984 6 dmem_client_request_get[6]
port 80 nsew signal output
rlabel metal3 s 0 128528 800 128648 6 dmem_client_request_get[70]
port 81 nsew signal output
rlabel metal3 s 0 129752 800 129872 6 dmem_client_request_get[71]
port 82 nsew signal output
rlabel metal3 s 0 130840 800 130960 6 dmem_client_request_get[72]
port 83 nsew signal output
rlabel metal3 s 0 132064 800 132184 6 dmem_client_request_get[73]
port 84 nsew signal output
rlabel metal3 s 0 133288 800 133408 6 dmem_client_request_get[74]
port 85 nsew signal output
rlabel metal3 s 0 134512 800 134632 6 dmem_client_request_get[75]
port 86 nsew signal output
rlabel metal3 s 0 135736 800 135856 6 dmem_client_request_get[76]
port 87 nsew signal output
rlabel metal3 s 0 136960 800 137080 6 dmem_client_request_get[77]
port 88 nsew signal output
rlabel metal3 s 0 138184 800 138304 6 dmem_client_request_get[78]
port 89 nsew signal output
rlabel metal3 s 0 139408 800 139528 6 dmem_client_request_get[79]
port 90 nsew signal output
rlabel metal3 s 0 22176 800 22296 6 dmem_client_request_get[7]
port 91 nsew signal output
rlabel metal3 s 0 140632 800 140752 6 dmem_client_request_get[80]
port 92 nsew signal output
rlabel metal3 s 0 141720 800 141840 6 dmem_client_request_get[81]
port 93 nsew signal output
rlabel metal3 s 0 142944 800 143064 6 dmem_client_request_get[82]
port 94 nsew signal output
rlabel metal3 s 0 144168 800 144288 6 dmem_client_request_get[83]
port 95 nsew signal output
rlabel metal3 s 0 145392 800 145512 6 dmem_client_request_get[84]
port 96 nsew signal output
rlabel metal3 s 0 146616 800 146736 6 dmem_client_request_get[85]
port 97 nsew signal output
rlabel metal3 s 0 147840 800 147960 6 dmem_client_request_get[86]
port 98 nsew signal output
rlabel metal3 s 0 149064 800 149184 6 dmem_client_request_get[87]
port 99 nsew signal output
rlabel metal3 s 0 150288 800 150408 6 dmem_client_request_get[88]
port 100 nsew signal output
rlabel metal3 s 0 151376 800 151496 6 dmem_client_request_get[89]
port 101 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 dmem_client_request_get[8]
port 102 nsew signal output
rlabel metal3 s 0 152600 800 152720 6 dmem_client_request_get[90]
port 103 nsew signal output
rlabel metal3 s 0 153824 800 153944 6 dmem_client_request_get[91]
port 104 nsew signal output
rlabel metal3 s 0 155048 800 155168 6 dmem_client_request_get[92]
port 105 nsew signal output
rlabel metal3 s 0 156272 800 156392 6 dmem_client_request_get[93]
port 106 nsew signal output
rlabel metal3 s 0 157496 800 157616 6 dmem_client_request_get[94]
port 107 nsew signal output
rlabel metal3 s 0 158720 800 158840 6 dmem_client_request_get[95]
port 108 nsew signal output
rlabel metal3 s 0 159944 800 160064 6 dmem_client_request_get[96]
port 109 nsew signal output
rlabel metal3 s 0 161032 800 161152 6 dmem_client_request_get[97]
port 110 nsew signal output
rlabel metal3 s 0 162256 800 162376 6 dmem_client_request_get[98]
port 111 nsew signal output
rlabel metal3 s 0 163480 800 163600 6 dmem_client_request_get[99]
port 112 nsew signal output
rlabel metal3 s 0 27072 800 27192 6 dmem_client_request_get[9]
port 113 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 dmem_client_response_put[0]
port 114 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 dmem_client_response_put[10]
port 115 nsew signal input
rlabel metal3 s 0 33056 800 33176 6 dmem_client_response_put[11]
port 116 nsew signal input
rlabel metal3 s 0 35504 800 35624 6 dmem_client_response_put[12]
port 117 nsew signal input
rlabel metal3 s 0 37952 800 38072 6 dmem_client_response_put[13]
port 118 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 dmem_client_response_put[14]
port 119 nsew signal input
rlabel metal3 s 0 42712 800 42832 6 dmem_client_response_put[15]
port 120 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 dmem_client_response_put[16]
port 121 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 dmem_client_response_put[17]
port 122 nsew signal input
rlabel metal3 s 0 50056 800 50176 6 dmem_client_response_put[18]
port 123 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 dmem_client_response_put[19]
port 124 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 dmem_client_response_put[1]
port 125 nsew signal input
rlabel metal3 s 0 54816 800 54936 6 dmem_client_response_put[20]
port 126 nsew signal input
rlabel metal3 s 0 57264 800 57384 6 dmem_client_response_put[21]
port 127 nsew signal input
rlabel metal3 s 0 59712 800 59832 6 dmem_client_response_put[22]
port 128 nsew signal input
rlabel metal3 s 0 62024 800 62144 6 dmem_client_response_put[23]
port 129 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 dmem_client_response_put[24]
port 130 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 dmem_client_response_put[25]
port 131 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 dmem_client_response_put[26]
port 132 nsew signal input
rlabel metal3 s 0 71680 800 71800 6 dmem_client_response_put[27]
port 133 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 dmem_client_response_put[28]
port 134 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 dmem_client_response_put[29]
port 135 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 dmem_client_response_put[2]
port 136 nsew signal input
rlabel metal3 s 0 79024 800 79144 6 dmem_client_response_put[30]
port 137 nsew signal input
rlabel metal3 s 0 81336 800 81456 6 dmem_client_response_put[31]
port 138 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 dmem_client_response_put[3]
port 139 nsew signal input
rlabel metal3 s 0 16192 800 16312 6 dmem_client_response_put[4]
port 140 nsew signal input
rlabel metal3 s 0 18640 800 18760 6 dmem_client_response_put[5]
port 141 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 dmem_client_response_put[6]
port 142 nsew signal input
rlabel metal3 s 0 23400 800 23520 6 dmem_client_response_put[7]
port 143 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 dmem_client_response_put[8]
port 144 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 dmem_client_response_put[9]
port 145 nsew signal input
rlabel metal2 s 9678 169475 9734 170275 6 imem_client_request_get[0]
port 146 nsew signal output
rlabel metal2 s 53378 169475 53434 170275 6 imem_client_request_get[10]
port 147 nsew signal output
rlabel metal2 s 57794 169475 57850 170275 6 imem_client_request_get[11]
port 148 nsew signal output
rlabel metal2 s 62118 169475 62174 170275 6 imem_client_request_get[12]
port 149 nsew signal output
rlabel metal2 s 66534 169475 66590 170275 6 imem_client_request_get[13]
port 150 nsew signal output
rlabel metal2 s 70858 169475 70914 170275 6 imem_client_request_get[14]
port 151 nsew signal output
rlabel metal2 s 75274 169475 75330 170275 6 imem_client_request_get[15]
port 152 nsew signal output
rlabel metal2 s 79598 169475 79654 170275 6 imem_client_request_get[16]
port 153 nsew signal output
rlabel metal2 s 84014 169475 84070 170275 6 imem_client_request_get[17]
port 154 nsew signal output
rlabel metal2 s 88338 169475 88394 170275 6 imem_client_request_get[18]
port 155 nsew signal output
rlabel metal2 s 92754 169475 92810 170275 6 imem_client_request_get[19]
port 156 nsew signal output
rlabel metal2 s 14094 169475 14150 170275 6 imem_client_request_get[1]
port 157 nsew signal output
rlabel metal2 s 97078 169475 97134 170275 6 imem_client_request_get[20]
port 158 nsew signal output
rlabel metal2 s 101494 169475 101550 170275 6 imem_client_request_get[21]
port 159 nsew signal output
rlabel metal2 s 105818 169475 105874 170275 6 imem_client_request_get[22]
port 160 nsew signal output
rlabel metal2 s 110234 169475 110290 170275 6 imem_client_request_get[23]
port 161 nsew signal output
rlabel metal2 s 114558 169475 114614 170275 6 imem_client_request_get[24]
port 162 nsew signal output
rlabel metal2 s 118882 169475 118938 170275 6 imem_client_request_get[25]
port 163 nsew signal output
rlabel metal2 s 123298 169475 123354 170275 6 imem_client_request_get[26]
port 164 nsew signal output
rlabel metal2 s 127622 169475 127678 170275 6 imem_client_request_get[27]
port 165 nsew signal output
rlabel metal2 s 132038 169475 132094 170275 6 imem_client_request_get[28]
port 166 nsew signal output
rlabel metal2 s 136362 169475 136418 170275 6 imem_client_request_get[29]
port 167 nsew signal output
rlabel metal2 s 18418 169475 18474 170275 6 imem_client_request_get[2]
port 168 nsew signal output
rlabel metal2 s 140778 169475 140834 170275 6 imem_client_request_get[30]
port 169 nsew signal output
rlabel metal2 s 145102 169475 145158 170275 6 imem_client_request_get[31]
port 170 nsew signal output
rlabel metal2 s 22834 169475 22890 170275 6 imem_client_request_get[3]
port 171 nsew signal output
rlabel metal2 s 27158 169475 27214 170275 6 imem_client_request_get[4]
port 172 nsew signal output
rlabel metal2 s 31574 169475 31630 170275 6 imem_client_request_get[5]
port 173 nsew signal output
rlabel metal2 s 35898 169475 35954 170275 6 imem_client_request_get[6]
port 174 nsew signal output
rlabel metal2 s 40314 169475 40370 170275 6 imem_client_request_get[7]
port 175 nsew signal output
rlabel metal2 s 44638 169475 44694 170275 6 imem_client_request_get[8]
port 176 nsew signal output
rlabel metal2 s 49054 169475 49110 170275 6 imem_client_request_get[9]
port 177 nsew signal output
rlabel metal2 s 11886 169475 11942 170275 6 imem_client_response_put[0]
port 178 nsew signal input
rlabel metal2 s 55586 169475 55642 170275 6 imem_client_response_put[10]
port 179 nsew signal input
rlabel metal2 s 59910 169475 59966 170275 6 imem_client_response_put[11]
port 180 nsew signal input
rlabel metal2 s 64326 169475 64382 170275 6 imem_client_response_put[12]
port 181 nsew signal input
rlabel metal2 s 68650 169475 68706 170275 6 imem_client_response_put[13]
port 182 nsew signal input
rlabel metal2 s 73066 169475 73122 170275 6 imem_client_response_put[14]
port 183 nsew signal input
rlabel metal2 s 77390 169475 77446 170275 6 imem_client_response_put[15]
port 184 nsew signal input
rlabel metal2 s 81806 169475 81862 170275 6 imem_client_response_put[16]
port 185 nsew signal input
rlabel metal2 s 86130 169475 86186 170275 6 imem_client_response_put[17]
port 186 nsew signal input
rlabel metal2 s 90546 169475 90602 170275 6 imem_client_response_put[18]
port 187 nsew signal input
rlabel metal2 s 94870 169475 94926 170275 6 imem_client_response_put[19]
port 188 nsew signal input
rlabel metal2 s 16302 169475 16358 170275 6 imem_client_response_put[1]
port 189 nsew signal input
rlabel metal2 s 99286 169475 99342 170275 6 imem_client_response_put[20]
port 190 nsew signal input
rlabel metal2 s 103610 169475 103666 170275 6 imem_client_response_put[21]
port 191 nsew signal input
rlabel metal2 s 108026 169475 108082 170275 6 imem_client_response_put[22]
port 192 nsew signal input
rlabel metal2 s 112350 169475 112406 170275 6 imem_client_response_put[23]
port 193 nsew signal input
rlabel metal2 s 116766 169475 116822 170275 6 imem_client_response_put[24]
port 194 nsew signal input
rlabel metal2 s 121090 169475 121146 170275 6 imem_client_response_put[25]
port 195 nsew signal input
rlabel metal2 s 125506 169475 125562 170275 6 imem_client_response_put[26]
port 196 nsew signal input
rlabel metal2 s 129830 169475 129886 170275 6 imem_client_response_put[27]
port 197 nsew signal input
rlabel metal2 s 134246 169475 134302 170275 6 imem_client_response_put[28]
port 198 nsew signal input
rlabel metal2 s 138570 169475 138626 170275 6 imem_client_response_put[29]
port 199 nsew signal input
rlabel metal2 s 20626 169475 20682 170275 6 imem_client_response_put[2]
port 200 nsew signal input
rlabel metal2 s 142986 169475 143042 170275 6 imem_client_response_put[30]
port 201 nsew signal input
rlabel metal2 s 147310 169475 147366 170275 6 imem_client_response_put[31]
port 202 nsew signal input
rlabel metal2 s 25042 169475 25098 170275 6 imem_client_response_put[3]
port 203 nsew signal input
rlabel metal2 s 29366 169475 29422 170275 6 imem_client_response_put[4]
port 204 nsew signal input
rlabel metal2 s 33782 169475 33838 170275 6 imem_client_response_put[5]
port 205 nsew signal input
rlabel metal2 s 38106 169475 38162 170275 6 imem_client_response_put[6]
port 206 nsew signal input
rlabel metal2 s 42522 169475 42578 170275 6 imem_client_response_put[7]
port 207 nsew signal input
rlabel metal2 s 46846 169475 46902 170275 6 imem_client_response_put[8]
port 208 nsew signal input
rlabel metal2 s 51262 169475 51318 170275 6 imem_client_response_put[9]
port 209 nsew signal input
rlabel metal2 s 151726 169475 151782 170275 6 readPC[0]
port 210 nsew signal output
rlabel metal3 s 167331 157904 168131 158024 6 readPC[10]
port 211 nsew signal output
rlabel metal3 s 167331 159400 168131 159520 6 readPC[11]
port 212 nsew signal output
rlabel metal3 s 167331 160760 168131 160880 6 readPC[12]
port 213 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 readPC[13]
port 214 nsew signal output
rlabel metal2 s 84014 0 84070 800 6 readPC[14]
port 215 nsew signal output
rlabel metal2 s 158258 169475 158314 170275 6 readPC[15]
port 216 nsew signal output
rlabel metal2 s 160466 169475 160522 170275 6 readPC[16]
port 217 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 readPC[17]
port 218 nsew signal output
rlabel metal3 s 167331 162256 168131 162376 6 readPC[18]
port 219 nsew signal output
rlabel metal3 s 167331 163616 168131 163736 6 readPC[19]
port 220 nsew signal output
rlabel metal3 s 167331 155048 168131 155168 6 readPC[1]
port 221 nsew signal output
rlabel metal3 s 0 168376 800 168496 6 readPC[20]
port 222 nsew signal output
rlabel metal3 s 0 169600 800 169720 6 readPC[21]
port 223 nsew signal output
rlabel metal2 s 162582 169475 162638 170275 6 readPC[22]
port 224 nsew signal output
rlabel metal2 s 121366 0 121422 800 6 readPC[23]
port 225 nsew signal output
rlabel metal3 s 167331 165112 168131 165232 6 readPC[24]
port 226 nsew signal output
rlabel metal2 s 140042 0 140098 800 6 readPC[25]
port 227 nsew signal output
rlabel metal3 s 167331 166608 168131 166728 6 readPC[26]
port 228 nsew signal output
rlabel metal2 s 164790 169475 164846 170275 6 readPC[27]
port 229 nsew signal output
rlabel metal2 s 166998 169475 167054 170275 6 readPC[28]
port 230 nsew signal output
rlabel metal2 s 158718 0 158774 800 6 readPC[29]
port 231 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 readPC[2]
port 232 nsew signal output
rlabel metal3 s 167331 167968 168131 168088 6 readPC[30]
port 233 nsew signal output
rlabel metal3 s 167331 169464 168131 169584 6 readPC[31]
port 234 nsew signal output
rlabel metal2 s 153842 169475 153898 170275 6 readPC[3]
port 235 nsew signal output
rlabel metal3 s 0 164704 800 164824 6 readPC[4]
port 236 nsew signal output
rlabel metal2 s 156050 169475 156106 170275 6 readPC[5]
port 237 nsew signal output
rlabel metal3 s 167331 156408 168131 156528 6 readPC[6]
port 238 nsew signal output
rlabel metal3 s 0 165928 800 166048 6 readPC[7]
port 239 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 readPC[8]
port 240 nsew signal output
rlabel metal3 s 0 167152 800 167272 6 readPC[9]
port 241 nsew signal output
rlabel metal3 s 167331 688 168131 808 6 sysmem_client_ack_i
port 242 nsew signal input
rlabel metal3 s 167331 9256 168131 9376 6 sysmem_client_adr_o[0]
port 243 nsew signal output
rlabel metal3 s 167331 58352 168131 58472 6 sysmem_client_adr_o[10]
port 244 nsew signal output
rlabel metal3 s 167331 62704 168131 62824 6 sysmem_client_adr_o[11]
port 245 nsew signal output
rlabel metal3 s 167331 67056 168131 67176 6 sysmem_client_adr_o[12]
port 246 nsew signal output
rlabel metal3 s 167331 71272 168131 71392 6 sysmem_client_adr_o[13]
port 247 nsew signal output
rlabel metal3 s 167331 75624 168131 75744 6 sysmem_client_adr_o[14]
port 248 nsew signal output
rlabel metal3 s 167331 79976 168131 80096 6 sysmem_client_adr_o[15]
port 249 nsew signal output
rlabel metal3 s 167331 84328 168131 84448 6 sysmem_client_adr_o[16]
port 250 nsew signal output
rlabel metal3 s 167331 88680 168131 88800 6 sysmem_client_adr_o[17]
port 251 nsew signal output
rlabel metal3 s 167331 93032 168131 93152 6 sysmem_client_adr_o[18]
port 252 nsew signal output
rlabel metal3 s 167331 97248 168131 97368 6 sysmem_client_adr_o[19]
port 253 nsew signal output
rlabel metal3 s 167331 15104 168131 15224 6 sysmem_client_adr_o[1]
port 254 nsew signal output
rlabel metal3 s 167331 101600 168131 101720 6 sysmem_client_adr_o[20]
port 255 nsew signal output
rlabel metal3 s 167331 105952 168131 106072 6 sysmem_client_adr_o[21]
port 256 nsew signal output
rlabel metal3 s 167331 110304 168131 110424 6 sysmem_client_adr_o[22]
port 257 nsew signal output
rlabel metal3 s 167331 114656 168131 114776 6 sysmem_client_adr_o[23]
port 258 nsew signal output
rlabel metal3 s 167331 119008 168131 119128 6 sysmem_client_adr_o[24]
port 259 nsew signal output
rlabel metal3 s 167331 123224 168131 123344 6 sysmem_client_adr_o[25]
port 260 nsew signal output
rlabel metal3 s 167331 127576 168131 127696 6 sysmem_client_adr_o[26]
port 261 nsew signal output
rlabel metal3 s 167331 131928 168131 132048 6 sysmem_client_adr_o[27]
port 262 nsew signal output
rlabel metal3 s 167331 136280 168131 136400 6 sysmem_client_adr_o[28]
port 263 nsew signal output
rlabel metal3 s 167331 140632 168131 140752 6 sysmem_client_adr_o[29]
port 264 nsew signal output
rlabel metal3 s 167331 20816 168131 20936 6 sysmem_client_adr_o[2]
port 265 nsew signal output
rlabel metal3 s 167331 144984 168131 145104 6 sysmem_client_adr_o[30]
port 266 nsew signal output
rlabel metal3 s 167331 149200 168131 149320 6 sysmem_client_adr_o[31]
port 267 nsew signal output
rlabel metal3 s 167331 26528 168131 26648 6 sysmem_client_adr_o[3]
port 268 nsew signal output
rlabel metal3 s 167331 32376 168131 32496 6 sysmem_client_adr_o[4]
port 269 nsew signal output
rlabel metal3 s 167331 36728 168131 36848 6 sysmem_client_adr_o[5]
port 270 nsew signal output
rlabel metal3 s 167331 41080 168131 41200 6 sysmem_client_adr_o[6]
port 271 nsew signal output
rlabel metal3 s 167331 45296 168131 45416 6 sysmem_client_adr_o[7]
port 272 nsew signal output
rlabel metal3 s 167331 49648 168131 49768 6 sysmem_client_adr_o[8]
port 273 nsew signal output
rlabel metal3 s 167331 54000 168131 54120 6 sysmem_client_adr_o[9]
port 274 nsew signal output
rlabel metal3 s 167331 2048 168131 2168 6 sysmem_client_cyc_o
port 275 nsew signal output
rlabel metal3 s 167331 10752 168131 10872 6 sysmem_client_dat_i[0]
port 276 nsew signal input
rlabel metal3 s 167331 59848 168131 59968 6 sysmem_client_dat_i[10]
port 277 nsew signal input
rlabel metal3 s 167331 64064 168131 64184 6 sysmem_client_dat_i[11]
port 278 nsew signal input
rlabel metal3 s 167331 68416 168131 68536 6 sysmem_client_dat_i[12]
port 279 nsew signal input
rlabel metal3 s 167331 72768 168131 72888 6 sysmem_client_dat_i[13]
port 280 nsew signal input
rlabel metal3 s 167331 77120 168131 77240 6 sysmem_client_dat_i[14]
port 281 nsew signal input
rlabel metal3 s 167331 81472 168131 81592 6 sysmem_client_dat_i[15]
port 282 nsew signal input
rlabel metal3 s 167331 85824 168131 85944 6 sysmem_client_dat_i[16]
port 283 nsew signal input
rlabel metal3 s 167331 90040 168131 90160 6 sysmem_client_dat_i[17]
port 284 nsew signal input
rlabel metal3 s 167331 94392 168131 94512 6 sysmem_client_dat_i[18]
port 285 nsew signal input
rlabel metal3 s 167331 98744 168131 98864 6 sysmem_client_dat_i[19]
port 286 nsew signal input
rlabel metal3 s 167331 16464 168131 16584 6 sysmem_client_dat_i[1]
port 287 nsew signal input
rlabel metal3 s 167331 103096 168131 103216 6 sysmem_client_dat_i[20]
port 288 nsew signal input
rlabel metal3 s 167331 107448 168131 107568 6 sysmem_client_dat_i[21]
port 289 nsew signal input
rlabel metal3 s 167331 111664 168131 111784 6 sysmem_client_dat_i[22]
port 290 nsew signal input
rlabel metal3 s 167331 116016 168131 116136 6 sysmem_client_dat_i[23]
port 291 nsew signal input
rlabel metal3 s 167331 120368 168131 120488 6 sysmem_client_dat_i[24]
port 292 nsew signal input
rlabel metal3 s 167331 124720 168131 124840 6 sysmem_client_dat_i[25]
port 293 nsew signal input
rlabel metal3 s 167331 129072 168131 129192 6 sysmem_client_dat_i[26]
port 294 nsew signal input
rlabel metal3 s 167331 133424 168131 133544 6 sysmem_client_dat_i[27]
port 295 nsew signal input
rlabel metal3 s 167331 137640 168131 137760 6 sysmem_client_dat_i[28]
port 296 nsew signal input
rlabel metal3 s 167331 141992 168131 142112 6 sysmem_client_dat_i[29]
port 297 nsew signal input
rlabel metal3 s 167331 22312 168131 22432 6 sysmem_client_dat_i[2]
port 298 nsew signal input
rlabel metal3 s 167331 146344 168131 146464 6 sysmem_client_dat_i[30]
port 299 nsew signal input
rlabel metal3 s 167331 150696 168131 150816 6 sysmem_client_dat_i[31]
port 300 nsew signal input
rlabel metal3 s 167331 28024 168131 28144 6 sysmem_client_dat_i[3]
port 301 nsew signal input
rlabel metal3 s 167331 33872 168131 33992 6 sysmem_client_dat_i[4]
port 302 nsew signal input
rlabel metal3 s 167331 38088 168131 38208 6 sysmem_client_dat_i[5]
port 303 nsew signal input
rlabel metal3 s 167331 42440 168131 42560 6 sysmem_client_dat_i[6]
port 304 nsew signal input
rlabel metal3 s 167331 46792 168131 46912 6 sysmem_client_dat_i[7]
port 305 nsew signal input
rlabel metal3 s 167331 51144 168131 51264 6 sysmem_client_dat_i[8]
port 306 nsew signal input
rlabel metal3 s 167331 55496 168131 55616 6 sysmem_client_dat_i[9]
port 307 nsew signal input
rlabel metal3 s 167331 12112 168131 12232 6 sysmem_client_dat_o[0]
port 308 nsew signal output
rlabel metal3 s 167331 61208 168131 61328 6 sysmem_client_dat_o[10]
port 309 nsew signal output
rlabel metal3 s 167331 65560 168131 65680 6 sysmem_client_dat_o[11]
port 310 nsew signal output
rlabel metal3 s 167331 69912 168131 70032 6 sysmem_client_dat_o[12]
port 311 nsew signal output
rlabel metal3 s 167331 74264 168131 74384 6 sysmem_client_dat_o[13]
port 312 nsew signal output
rlabel metal3 s 167331 78480 168131 78600 6 sysmem_client_dat_o[14]
port 313 nsew signal output
rlabel metal3 s 167331 82832 168131 82952 6 sysmem_client_dat_o[15]
port 314 nsew signal output
rlabel metal3 s 167331 87184 168131 87304 6 sysmem_client_dat_o[16]
port 315 nsew signal output
rlabel metal3 s 167331 91536 168131 91656 6 sysmem_client_dat_o[17]
port 316 nsew signal output
rlabel metal3 s 167331 95888 168131 96008 6 sysmem_client_dat_o[18]
port 317 nsew signal output
rlabel metal3 s 167331 100240 168131 100360 6 sysmem_client_dat_o[19]
port 318 nsew signal output
rlabel metal3 s 167331 17960 168131 18080 6 sysmem_client_dat_o[1]
port 319 nsew signal output
rlabel metal3 s 167331 104456 168131 104576 6 sysmem_client_dat_o[20]
port 320 nsew signal output
rlabel metal3 s 167331 108808 168131 108928 6 sysmem_client_dat_o[21]
port 321 nsew signal output
rlabel metal3 s 167331 113160 168131 113280 6 sysmem_client_dat_o[22]
port 322 nsew signal output
rlabel metal3 s 167331 117512 168131 117632 6 sysmem_client_dat_o[23]
port 323 nsew signal output
rlabel metal3 s 167331 121864 168131 121984 6 sysmem_client_dat_o[24]
port 324 nsew signal output
rlabel metal3 s 167331 126216 168131 126336 6 sysmem_client_dat_o[25]
port 325 nsew signal output
rlabel metal3 s 167331 130432 168131 130552 6 sysmem_client_dat_o[26]
port 326 nsew signal output
rlabel metal3 s 167331 134784 168131 134904 6 sysmem_client_dat_o[27]
port 327 nsew signal output
rlabel metal3 s 167331 139136 168131 139256 6 sysmem_client_dat_o[28]
port 328 nsew signal output
rlabel metal3 s 167331 143488 168131 143608 6 sysmem_client_dat_o[29]
port 329 nsew signal output
rlabel metal3 s 167331 23672 168131 23792 6 sysmem_client_dat_o[2]
port 330 nsew signal output
rlabel metal3 s 167331 147840 168131 147960 6 sysmem_client_dat_o[30]
port 331 nsew signal output
rlabel metal3 s 167331 152192 168131 152312 6 sysmem_client_dat_o[31]
port 332 nsew signal output
rlabel metal3 s 167331 29520 168131 29640 6 sysmem_client_dat_o[3]
port 333 nsew signal output
rlabel metal3 s 167331 35232 168131 35352 6 sysmem_client_dat_o[4]
port 334 nsew signal output
rlabel metal3 s 167331 39584 168131 39704 6 sysmem_client_dat_o[5]
port 335 nsew signal output
rlabel metal3 s 167331 43936 168131 44056 6 sysmem_client_dat_o[6]
port 336 nsew signal output
rlabel metal3 s 167331 48288 168131 48408 6 sysmem_client_dat_o[7]
port 337 nsew signal output
rlabel metal3 s 167331 52504 168131 52624 6 sysmem_client_dat_o[8]
port 338 nsew signal output
rlabel metal3 s 167331 56856 168131 56976 6 sysmem_client_dat_o[9]
port 339 nsew signal output
rlabel metal3 s 167331 3544 168131 3664 6 sysmem_client_err_i
port 340 nsew signal input
rlabel metal3 s 167331 4904 168131 5024 6 sysmem_client_rty_i
port 341 nsew signal input
rlabel metal3 s 167331 13608 168131 13728 6 sysmem_client_sel_o[0]
port 342 nsew signal output
rlabel metal3 s 167331 19320 168131 19440 6 sysmem_client_sel_o[1]
port 343 nsew signal output
rlabel metal3 s 167331 25168 168131 25288 6 sysmem_client_sel_o[2]
port 344 nsew signal output
rlabel metal3 s 167331 30880 168131 31000 6 sysmem_client_sel_o[3]
port 345 nsew signal output
rlabel metal3 s 167331 6400 168131 6520 6 sysmem_client_stb_o
port 346 nsew signal output
rlabel metal3 s 167331 7896 168131 8016 6 sysmem_client_we_o
port 347 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 168131 170275
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 73379078
string GDS_FILE /home/q3k/sky130/qf105/openlane/mkLanaiCPU/runs/mkLanaiCPU/results/finishing/mkLanaiCPU.magic.gds
string GDS_START 1533176
<< end >>

