VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mkQF100Memory
  CLASS BLOCK ;
  FOREIGN mkQF100Memory ;
  ORIGIN 0.000 0.000 ;
  SIZE 319.240 BY 329.960 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 0.000 0.830 4.000 ;
    END
  END CLK
  PIN EN_memory_dmem_request_put
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END EN_memory_dmem_request_put
  PIN EN_memory_dmem_response_get
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 4.000 ;
    END
  END EN_memory_dmem_response_get
  PIN EN_memory_imem_request_put
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END EN_memory_imem_request_put
  PIN EN_memory_imem_response_get
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END EN_memory_imem_response_get
  PIN RDY_memory_dmem_request_put
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END RDY_memory_dmem_request_put
  PIN RDY_memory_dmem_response_get
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END RDY_memory_dmem_response_get
  PIN RDY_memory_imem_request_put
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END RDY_memory_imem_request_put
  PIN RDY_memory_imem_response_get
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END RDY_memory_imem_response_get
  PIN RST_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END RST_N
  PIN memory_dmem_request_put[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END memory_dmem_request_put[0]
  PIN memory_dmem_request_put[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END memory_dmem_request_put[10]
  PIN memory_dmem_request_put[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END memory_dmem_request_put[11]
  PIN memory_dmem_request_put[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END memory_dmem_request_put[12]
  PIN memory_dmem_request_put[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END memory_dmem_request_put[13]
  PIN memory_dmem_request_put[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END memory_dmem_request_put[14]
  PIN memory_dmem_request_put[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END memory_dmem_request_put[15]
  PIN memory_dmem_request_put[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END memory_dmem_request_put[16]
  PIN memory_dmem_request_put[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END memory_dmem_request_put[17]
  PIN memory_dmem_request_put[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END memory_dmem_request_put[18]
  PIN memory_dmem_request_put[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END memory_dmem_request_put[19]
  PIN memory_dmem_request_put[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END memory_dmem_request_put[1]
  PIN memory_dmem_request_put[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END memory_dmem_request_put[20]
  PIN memory_dmem_request_put[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END memory_dmem_request_put[21]
  PIN memory_dmem_request_put[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END memory_dmem_request_put[22]
  PIN memory_dmem_request_put[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END memory_dmem_request_put[23]
  PIN memory_dmem_request_put[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END memory_dmem_request_put[24]
  PIN memory_dmem_request_put[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END memory_dmem_request_put[25]
  PIN memory_dmem_request_put[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END memory_dmem_request_put[26]
  PIN memory_dmem_request_put[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END memory_dmem_request_put[27]
  PIN memory_dmem_request_put[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END memory_dmem_request_put[28]
  PIN memory_dmem_request_put[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END memory_dmem_request_put[29]
  PIN memory_dmem_request_put[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END memory_dmem_request_put[2]
  PIN memory_dmem_request_put[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END memory_dmem_request_put[30]
  PIN memory_dmem_request_put[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END memory_dmem_request_put[31]
  PIN memory_dmem_request_put[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END memory_dmem_request_put[32]
  PIN memory_dmem_request_put[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END memory_dmem_request_put[33]
  PIN memory_dmem_request_put[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END memory_dmem_request_put[34]
  PIN memory_dmem_request_put[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END memory_dmem_request_put[35]
  PIN memory_dmem_request_put[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 4.000 ;
    END
  END memory_dmem_request_put[36]
  PIN memory_dmem_request_put[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END memory_dmem_request_put[37]
  PIN memory_dmem_request_put[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END memory_dmem_request_put[38]
  PIN memory_dmem_request_put[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END memory_dmem_request_put[39]
  PIN memory_dmem_request_put[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END memory_dmem_request_put[3]
  PIN memory_dmem_request_put[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END memory_dmem_request_put[40]
  PIN memory_dmem_request_put[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END memory_dmem_request_put[41]
  PIN memory_dmem_request_put[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END memory_dmem_request_put[42]
  PIN memory_dmem_request_put[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END memory_dmem_request_put[43]
  PIN memory_dmem_request_put[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END memory_dmem_request_put[44]
  PIN memory_dmem_request_put[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END memory_dmem_request_put[45]
  PIN memory_dmem_request_put[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 0.000 236.350 4.000 ;
    END
  END memory_dmem_request_put[46]
  PIN memory_dmem_request_put[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END memory_dmem_request_put[47]
  PIN memory_dmem_request_put[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 4.000 ;
    END
  END memory_dmem_request_put[48]
  PIN memory_dmem_request_put[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END memory_dmem_request_put[49]
  PIN memory_dmem_request_put[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END memory_dmem_request_put[4]
  PIN memory_dmem_request_put[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END memory_dmem_request_put[50]
  PIN memory_dmem_request_put[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END memory_dmem_request_put[51]
  PIN memory_dmem_request_put[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END memory_dmem_request_put[52]
  PIN memory_dmem_request_put[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END memory_dmem_request_put[53]
  PIN memory_dmem_request_put[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END memory_dmem_request_put[54]
  PIN memory_dmem_request_put[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END memory_dmem_request_put[55]
  PIN memory_dmem_request_put[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END memory_dmem_request_put[56]
  PIN memory_dmem_request_put[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END memory_dmem_request_put[57]
  PIN memory_dmem_request_put[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END memory_dmem_request_put[58]
  PIN memory_dmem_request_put[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END memory_dmem_request_put[59]
  PIN memory_dmem_request_put[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END memory_dmem_request_put[5]
  PIN memory_dmem_request_put[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END memory_dmem_request_put[60]
  PIN memory_dmem_request_put[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 0.000 259.350 4.000 ;
    END
  END memory_dmem_request_put[61]
  PIN memory_dmem_request_put[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END memory_dmem_request_put[62]
  PIN memory_dmem_request_put[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END memory_dmem_request_put[63]
  PIN memory_dmem_request_put[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END memory_dmem_request_put[64]
  PIN memory_dmem_request_put[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END memory_dmem_request_put[65]
  PIN memory_dmem_request_put[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END memory_dmem_request_put[66]
  PIN memory_dmem_request_put[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END memory_dmem_request_put[67]
  PIN memory_dmem_request_put[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END memory_dmem_request_put[68]
  PIN memory_dmem_request_put[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END memory_dmem_request_put[69]
  PIN memory_dmem_request_put[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END memory_dmem_request_put[6]
  PIN memory_dmem_request_put[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END memory_dmem_request_put[70]
  PIN memory_dmem_request_put[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END memory_dmem_request_put[71]
  PIN memory_dmem_request_put[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END memory_dmem_request_put[72]
  PIN memory_dmem_request_put[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END memory_dmem_request_put[73]
  PIN memory_dmem_request_put[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END memory_dmem_request_put[74]
  PIN memory_dmem_request_put[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END memory_dmem_request_put[75]
  PIN memory_dmem_request_put[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END memory_dmem_request_put[76]
  PIN memory_dmem_request_put[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 0.000 284.190 4.000 ;
    END
  END memory_dmem_request_put[77]
  PIN memory_dmem_request_put[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END memory_dmem_request_put[78]
  PIN memory_dmem_request_put[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END memory_dmem_request_put[79]
  PIN memory_dmem_request_put[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END memory_dmem_request_put[7]
  PIN memory_dmem_request_put[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END memory_dmem_request_put[80]
  PIN memory_dmem_request_put[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END memory_dmem_request_put[81]
  PIN memory_dmem_request_put[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END memory_dmem_request_put[82]
  PIN memory_dmem_request_put[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END memory_dmem_request_put[83]
  PIN memory_dmem_request_put[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END memory_dmem_request_put[84]
  PIN memory_dmem_request_put[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END memory_dmem_request_put[85]
  PIN memory_dmem_request_put[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 0.000 297.990 4.000 ;
    END
  END memory_dmem_request_put[86]
  PIN memory_dmem_request_put[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END memory_dmem_request_put[87]
  PIN memory_dmem_request_put[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END memory_dmem_request_put[88]
  PIN memory_dmem_request_put[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END memory_dmem_request_put[89]
  PIN memory_dmem_request_put[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END memory_dmem_request_put[8]
  PIN memory_dmem_request_put[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END memory_dmem_request_put[90]
  PIN memory_dmem_request_put[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END memory_dmem_request_put[91]
  PIN memory_dmem_request_put[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END memory_dmem_request_put[92]
  PIN memory_dmem_request_put[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END memory_dmem_request_put[93]
  PIN memory_dmem_request_put[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END memory_dmem_request_put[94]
  PIN memory_dmem_request_put[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END memory_dmem_request_put[95]
  PIN memory_dmem_request_put[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END memory_dmem_request_put[96]
  PIN memory_dmem_request_put[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END memory_dmem_request_put[97]
  PIN memory_dmem_request_put[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END memory_dmem_request_put[98]
  PIN memory_dmem_request_put[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END memory_dmem_request_put[99]
  PIN memory_dmem_request_put[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END memory_dmem_request_put[9]
  PIN memory_dmem_response_get[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END memory_dmem_response_get[0]
  PIN memory_dmem_response_get[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END memory_dmem_response_get[10]
  PIN memory_dmem_response_get[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END memory_dmem_response_get[11]
  PIN memory_dmem_response_get[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END memory_dmem_response_get[12]
  PIN memory_dmem_response_get[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END memory_dmem_response_get[13]
  PIN memory_dmem_response_get[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END memory_dmem_response_get[14]
  PIN memory_dmem_response_get[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END memory_dmem_response_get[15]
  PIN memory_dmem_response_get[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END memory_dmem_response_get[16]
  PIN memory_dmem_response_get[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END memory_dmem_response_get[17]
  PIN memory_dmem_response_get[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END memory_dmem_response_get[18]
  PIN memory_dmem_response_get[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END memory_dmem_response_get[19]
  PIN memory_dmem_response_get[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END memory_dmem_response_get[1]
  PIN memory_dmem_response_get[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END memory_dmem_response_get[20]
  PIN memory_dmem_response_get[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END memory_dmem_response_get[21]
  PIN memory_dmem_response_get[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END memory_dmem_response_get[22]
  PIN memory_dmem_response_get[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END memory_dmem_response_get[23]
  PIN memory_dmem_response_get[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END memory_dmem_response_get[24]
  PIN memory_dmem_response_get[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END memory_dmem_response_get[25]
  PIN memory_dmem_response_get[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END memory_dmem_response_get[26]
  PIN memory_dmem_response_get[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END memory_dmem_response_get[27]
  PIN memory_dmem_response_get[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END memory_dmem_response_get[28]
  PIN memory_dmem_response_get[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END memory_dmem_response_get[29]
  PIN memory_dmem_response_get[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END memory_dmem_response_get[2]
  PIN memory_dmem_response_get[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END memory_dmem_response_get[30]
  PIN memory_dmem_response_get[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END memory_dmem_response_get[31]
  PIN memory_dmem_response_get[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END memory_dmem_response_get[3]
  PIN memory_dmem_response_get[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END memory_dmem_response_get[4]
  PIN memory_dmem_response_get[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END memory_dmem_response_get[5]
  PIN memory_dmem_response_get[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END memory_dmem_response_get[6]
  PIN memory_dmem_response_get[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END memory_dmem_response_get[7]
  PIN memory_dmem_response_get[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END memory_dmem_response_get[8]
  PIN memory_dmem_response_get[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 4.000 ;
    END
  END memory_dmem_response_get[9]
  PIN memory_imem_request_put[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END memory_imem_request_put[0]
  PIN memory_imem_request_put[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END memory_imem_request_put[10]
  PIN memory_imem_request_put[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END memory_imem_request_put[11]
  PIN memory_imem_request_put[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END memory_imem_request_put[12]
  PIN memory_imem_request_put[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END memory_imem_request_put[13]
  PIN memory_imem_request_put[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END memory_imem_request_put[14]
  PIN memory_imem_request_put[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END memory_imem_request_put[15]
  PIN memory_imem_request_put[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 4.000 ;
    END
  END memory_imem_request_put[16]
  PIN memory_imem_request_put[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END memory_imem_request_put[17]
  PIN memory_imem_request_put[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END memory_imem_request_put[18]
  PIN memory_imem_request_put[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END memory_imem_request_put[19]
  PIN memory_imem_request_put[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END memory_imem_request_put[1]
  PIN memory_imem_request_put[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END memory_imem_request_put[20]
  PIN memory_imem_request_put[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END memory_imem_request_put[21]
  PIN memory_imem_request_put[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END memory_imem_request_put[22]
  PIN memory_imem_request_put[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END memory_imem_request_put[23]
  PIN memory_imem_request_put[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END memory_imem_request_put[24]
  PIN memory_imem_request_put[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END memory_imem_request_put[25]
  PIN memory_imem_request_put[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END memory_imem_request_put[26]
  PIN memory_imem_request_put[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END memory_imem_request_put[27]
  PIN memory_imem_request_put[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END memory_imem_request_put[28]
  PIN memory_imem_request_put[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END memory_imem_request_put[29]
  PIN memory_imem_request_put[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END memory_imem_request_put[2]
  PIN memory_imem_request_put[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END memory_imem_request_put[30]
  PIN memory_imem_request_put[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END memory_imem_request_put[31]
  PIN memory_imem_request_put[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END memory_imem_request_put[3]
  PIN memory_imem_request_put[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END memory_imem_request_put[4]
  PIN memory_imem_request_put[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END memory_imem_request_put[5]
  PIN memory_imem_request_put[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END memory_imem_request_put[6]
  PIN memory_imem_request_put[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END memory_imem_request_put[7]
  PIN memory_imem_request_put[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END memory_imem_request_put[8]
  PIN memory_imem_request_put[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END memory_imem_request_put[9]
  PIN memory_imem_response_get[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END memory_imem_response_get[0]
  PIN memory_imem_response_get[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END memory_imem_response_get[10]
  PIN memory_imem_response_get[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END memory_imem_response_get[11]
  PIN memory_imem_response_get[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END memory_imem_response_get[12]
  PIN memory_imem_response_get[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END memory_imem_response_get[13]
  PIN memory_imem_response_get[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END memory_imem_response_get[14]
  PIN memory_imem_response_get[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END memory_imem_response_get[15]
  PIN memory_imem_response_get[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END memory_imem_response_get[16]
  PIN memory_imem_response_get[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END memory_imem_response_get[17]
  PIN memory_imem_response_get[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END memory_imem_response_get[18]
  PIN memory_imem_response_get[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END memory_imem_response_get[19]
  PIN memory_imem_response_get[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END memory_imem_response_get[1]
  PIN memory_imem_response_get[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END memory_imem_response_get[20]
  PIN memory_imem_response_get[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END memory_imem_response_get[21]
  PIN memory_imem_response_get[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END memory_imem_response_get[22]
  PIN memory_imem_response_get[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END memory_imem_response_get[23]
  PIN memory_imem_response_get[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END memory_imem_response_get[24]
  PIN memory_imem_response_get[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END memory_imem_response_get[25]
  PIN memory_imem_response_get[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END memory_imem_response_get[26]
  PIN memory_imem_response_get[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END memory_imem_response_get[27]
  PIN memory_imem_response_get[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END memory_imem_response_get[28]
  PIN memory_imem_response_get[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END memory_imem_response_get[29]
  PIN memory_imem_response_get[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END memory_imem_response_get[2]
  PIN memory_imem_response_get[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END memory_imem_response_get[30]
  PIN memory_imem_response_get[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END memory_imem_response_get[31]
  PIN memory_imem_response_get[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END memory_imem_response_get[3]
  PIN memory_imem_response_get[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END memory_imem_response_get[4]
  PIN memory_imem_response_get[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END memory_imem_response_get[5]
  PIN memory_imem_response_get[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END memory_imem_response_get[6]
  PIN memory_imem_response_get[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END memory_imem_response_get[7]
  PIN memory_imem_response_get[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END memory_imem_response_get[8]
  PIN memory_imem_response_get[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END memory_imem_response_get[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 318.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 318.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 318.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 318.480 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 313.260 318.325 ;
      LAYER met1 ;
        RECT 0.530 4.460 318.250 318.480 ;
      LAYER met2 ;
        RECT 0.560 4.280 318.220 318.480 ;
        RECT 1.110 3.670 1.650 4.280 ;
        RECT 2.490 3.670 3.030 4.280 ;
        RECT 3.870 3.670 4.870 4.280 ;
        RECT 5.710 3.670 6.250 4.280 ;
        RECT 7.090 3.670 7.630 4.280 ;
        RECT 8.470 3.670 9.470 4.280 ;
        RECT 10.310 3.670 10.850 4.280 ;
        RECT 11.690 3.670 12.230 4.280 ;
        RECT 13.070 3.670 14.070 4.280 ;
        RECT 14.910 3.670 15.450 4.280 ;
        RECT 16.290 3.670 17.290 4.280 ;
        RECT 18.130 3.670 18.670 4.280 ;
        RECT 19.510 3.670 20.050 4.280 ;
        RECT 20.890 3.670 21.890 4.280 ;
        RECT 22.730 3.670 23.270 4.280 ;
        RECT 24.110 3.670 24.650 4.280 ;
        RECT 25.490 3.670 26.490 4.280 ;
        RECT 27.330 3.670 27.870 4.280 ;
        RECT 28.710 3.670 29.710 4.280 ;
        RECT 30.550 3.670 31.090 4.280 ;
        RECT 31.930 3.670 32.470 4.280 ;
        RECT 33.310 3.670 34.310 4.280 ;
        RECT 35.150 3.670 35.690 4.280 ;
        RECT 36.530 3.670 37.070 4.280 ;
        RECT 37.910 3.670 38.910 4.280 ;
        RECT 39.750 3.670 40.290 4.280 ;
        RECT 41.130 3.670 41.670 4.280 ;
        RECT 42.510 3.670 43.510 4.280 ;
        RECT 44.350 3.670 44.890 4.280 ;
        RECT 45.730 3.670 46.730 4.280 ;
        RECT 47.570 3.670 48.110 4.280 ;
        RECT 48.950 3.670 49.490 4.280 ;
        RECT 50.330 3.670 51.330 4.280 ;
        RECT 52.170 3.670 52.710 4.280 ;
        RECT 53.550 3.670 54.090 4.280 ;
        RECT 54.930 3.670 55.930 4.280 ;
        RECT 56.770 3.670 57.310 4.280 ;
        RECT 58.150 3.670 59.150 4.280 ;
        RECT 59.990 3.670 60.530 4.280 ;
        RECT 61.370 3.670 61.910 4.280 ;
        RECT 62.750 3.670 63.750 4.280 ;
        RECT 64.590 3.670 65.130 4.280 ;
        RECT 65.970 3.670 66.510 4.280 ;
        RECT 67.350 3.670 68.350 4.280 ;
        RECT 69.190 3.670 69.730 4.280 ;
        RECT 70.570 3.670 71.110 4.280 ;
        RECT 71.950 3.670 72.950 4.280 ;
        RECT 73.790 3.670 74.330 4.280 ;
        RECT 75.170 3.670 76.170 4.280 ;
        RECT 77.010 3.670 77.550 4.280 ;
        RECT 78.390 3.670 78.930 4.280 ;
        RECT 79.770 3.670 80.770 4.280 ;
        RECT 81.610 3.670 82.150 4.280 ;
        RECT 82.990 3.670 83.530 4.280 ;
        RECT 84.370 3.670 85.370 4.280 ;
        RECT 86.210 3.670 86.750 4.280 ;
        RECT 87.590 3.670 88.590 4.280 ;
        RECT 89.430 3.670 89.970 4.280 ;
        RECT 90.810 3.670 91.350 4.280 ;
        RECT 92.190 3.670 93.190 4.280 ;
        RECT 94.030 3.670 94.570 4.280 ;
        RECT 95.410 3.670 95.950 4.280 ;
        RECT 96.790 3.670 97.790 4.280 ;
        RECT 98.630 3.670 99.170 4.280 ;
        RECT 100.010 3.670 100.550 4.280 ;
        RECT 101.390 3.670 102.390 4.280 ;
        RECT 103.230 3.670 103.770 4.280 ;
        RECT 104.610 3.670 105.610 4.280 ;
        RECT 106.450 3.670 106.990 4.280 ;
        RECT 107.830 3.670 108.370 4.280 ;
        RECT 109.210 3.670 110.210 4.280 ;
        RECT 111.050 3.670 111.590 4.280 ;
        RECT 112.430 3.670 112.970 4.280 ;
        RECT 113.810 3.670 114.810 4.280 ;
        RECT 115.650 3.670 116.190 4.280 ;
        RECT 117.030 3.670 118.030 4.280 ;
        RECT 118.870 3.670 119.410 4.280 ;
        RECT 120.250 3.670 120.790 4.280 ;
        RECT 121.630 3.670 122.630 4.280 ;
        RECT 123.470 3.670 124.010 4.280 ;
        RECT 124.850 3.670 125.390 4.280 ;
        RECT 126.230 3.670 127.230 4.280 ;
        RECT 128.070 3.670 128.610 4.280 ;
        RECT 129.450 3.670 129.990 4.280 ;
        RECT 130.830 3.670 131.830 4.280 ;
        RECT 132.670 3.670 133.210 4.280 ;
        RECT 134.050 3.670 135.050 4.280 ;
        RECT 135.890 3.670 136.430 4.280 ;
        RECT 137.270 3.670 137.810 4.280 ;
        RECT 138.650 3.670 139.650 4.280 ;
        RECT 140.490 3.670 141.030 4.280 ;
        RECT 141.870 3.670 142.410 4.280 ;
        RECT 143.250 3.670 144.250 4.280 ;
        RECT 145.090 3.670 145.630 4.280 ;
        RECT 146.470 3.670 147.470 4.280 ;
        RECT 148.310 3.670 148.850 4.280 ;
        RECT 149.690 3.670 150.230 4.280 ;
        RECT 151.070 3.670 152.070 4.280 ;
        RECT 152.910 3.670 153.450 4.280 ;
        RECT 154.290 3.670 154.830 4.280 ;
        RECT 155.670 3.670 156.670 4.280 ;
        RECT 157.510 3.670 158.050 4.280 ;
        RECT 158.890 3.670 159.890 4.280 ;
        RECT 160.730 3.670 161.270 4.280 ;
        RECT 162.110 3.670 162.650 4.280 ;
        RECT 163.490 3.670 164.490 4.280 ;
        RECT 165.330 3.670 165.870 4.280 ;
        RECT 166.710 3.670 167.250 4.280 ;
        RECT 168.090 3.670 169.090 4.280 ;
        RECT 169.930 3.670 170.470 4.280 ;
        RECT 171.310 3.670 171.850 4.280 ;
        RECT 172.690 3.670 173.690 4.280 ;
        RECT 174.530 3.670 175.070 4.280 ;
        RECT 175.910 3.670 176.910 4.280 ;
        RECT 177.750 3.670 178.290 4.280 ;
        RECT 179.130 3.670 179.670 4.280 ;
        RECT 180.510 3.670 181.510 4.280 ;
        RECT 182.350 3.670 182.890 4.280 ;
        RECT 183.730 3.670 184.270 4.280 ;
        RECT 185.110 3.670 186.110 4.280 ;
        RECT 186.950 3.670 187.490 4.280 ;
        RECT 188.330 3.670 189.330 4.280 ;
        RECT 190.170 3.670 190.710 4.280 ;
        RECT 191.550 3.670 192.090 4.280 ;
        RECT 192.930 3.670 193.930 4.280 ;
        RECT 194.770 3.670 195.310 4.280 ;
        RECT 196.150 3.670 196.690 4.280 ;
        RECT 197.530 3.670 198.530 4.280 ;
        RECT 199.370 3.670 199.910 4.280 ;
        RECT 200.750 3.670 201.290 4.280 ;
        RECT 202.130 3.670 203.130 4.280 ;
        RECT 203.970 3.670 204.510 4.280 ;
        RECT 205.350 3.670 206.350 4.280 ;
        RECT 207.190 3.670 207.730 4.280 ;
        RECT 208.570 3.670 209.110 4.280 ;
        RECT 209.950 3.670 210.950 4.280 ;
        RECT 211.790 3.670 212.330 4.280 ;
        RECT 213.170 3.670 213.710 4.280 ;
        RECT 214.550 3.670 215.550 4.280 ;
        RECT 216.390 3.670 216.930 4.280 ;
        RECT 217.770 3.670 218.770 4.280 ;
        RECT 219.610 3.670 220.150 4.280 ;
        RECT 220.990 3.670 221.530 4.280 ;
        RECT 222.370 3.670 223.370 4.280 ;
        RECT 224.210 3.670 224.750 4.280 ;
        RECT 225.590 3.670 226.130 4.280 ;
        RECT 226.970 3.670 227.970 4.280 ;
        RECT 228.810 3.670 229.350 4.280 ;
        RECT 230.190 3.670 230.730 4.280 ;
        RECT 231.570 3.670 232.570 4.280 ;
        RECT 233.410 3.670 233.950 4.280 ;
        RECT 234.790 3.670 235.790 4.280 ;
        RECT 236.630 3.670 237.170 4.280 ;
        RECT 238.010 3.670 238.550 4.280 ;
        RECT 239.390 3.670 240.390 4.280 ;
        RECT 241.230 3.670 241.770 4.280 ;
        RECT 242.610 3.670 243.150 4.280 ;
        RECT 243.990 3.670 244.990 4.280 ;
        RECT 245.830 3.670 246.370 4.280 ;
        RECT 247.210 3.670 248.210 4.280 ;
        RECT 249.050 3.670 249.590 4.280 ;
        RECT 250.430 3.670 250.970 4.280 ;
        RECT 251.810 3.670 252.810 4.280 ;
        RECT 253.650 3.670 254.190 4.280 ;
        RECT 255.030 3.670 255.570 4.280 ;
        RECT 256.410 3.670 257.410 4.280 ;
        RECT 258.250 3.670 258.790 4.280 ;
        RECT 259.630 3.670 260.170 4.280 ;
        RECT 261.010 3.670 262.010 4.280 ;
        RECT 262.850 3.670 263.390 4.280 ;
        RECT 264.230 3.670 265.230 4.280 ;
        RECT 266.070 3.670 266.610 4.280 ;
        RECT 267.450 3.670 267.990 4.280 ;
        RECT 268.830 3.670 269.830 4.280 ;
        RECT 270.670 3.670 271.210 4.280 ;
        RECT 272.050 3.670 272.590 4.280 ;
        RECT 273.430 3.670 274.430 4.280 ;
        RECT 275.270 3.670 275.810 4.280 ;
        RECT 276.650 3.670 277.650 4.280 ;
        RECT 278.490 3.670 279.030 4.280 ;
        RECT 279.870 3.670 280.410 4.280 ;
        RECT 281.250 3.670 282.250 4.280 ;
        RECT 283.090 3.670 283.630 4.280 ;
        RECT 284.470 3.670 285.010 4.280 ;
        RECT 285.850 3.670 286.850 4.280 ;
        RECT 287.690 3.670 288.230 4.280 ;
        RECT 289.070 3.670 289.610 4.280 ;
        RECT 290.450 3.670 291.450 4.280 ;
        RECT 292.290 3.670 292.830 4.280 ;
        RECT 293.670 3.670 294.670 4.280 ;
        RECT 295.510 3.670 296.050 4.280 ;
        RECT 296.890 3.670 297.430 4.280 ;
        RECT 298.270 3.670 299.270 4.280 ;
        RECT 300.110 3.670 300.650 4.280 ;
        RECT 301.490 3.670 302.030 4.280 ;
        RECT 302.870 3.670 303.870 4.280 ;
        RECT 304.710 3.670 305.250 4.280 ;
        RECT 306.090 3.670 307.090 4.280 ;
        RECT 307.930 3.670 308.470 4.280 ;
        RECT 309.310 3.670 309.850 4.280 ;
        RECT 310.690 3.670 311.690 4.280 ;
        RECT 312.530 3.670 313.070 4.280 ;
        RECT 313.910 3.670 314.450 4.280 ;
        RECT 315.290 3.670 316.290 4.280 ;
        RECT 317.130 3.670 317.670 4.280 ;
      LAYER met3 ;
        RECT 3.030 10.715 315.955 318.405 ;
      LAYER met4 ;
        RECT 3.055 11.735 20.640 303.105 ;
        RECT 23.040 11.735 97.440 303.105 ;
        RECT 99.840 11.735 174.240 303.105 ;
        RECT 176.640 11.735 251.040 303.105 ;
        RECT 253.440 11.735 312.505 303.105 ;
  END
END mkQF100Memory
END LIBRARY

