magic
tech sky130A
magscale 1 2
timestamp 1647707691
<< obsli1 >>
rect 1104 2159 98808 57681
<< obsm1 >>
rect 198 1300 99714 58200
<< metal2 >>
rect 202 59200 258 60000
rect 662 59200 718 60000
rect 1122 59200 1178 60000
rect 1582 59200 1638 60000
rect 2042 59200 2098 60000
rect 2502 59200 2558 60000
rect 2962 59200 3018 60000
rect 3422 59200 3478 60000
rect 3974 59200 4030 60000
rect 4434 59200 4490 60000
rect 4894 59200 4950 60000
rect 5354 59200 5410 60000
rect 5814 59200 5870 60000
rect 6274 59200 6330 60000
rect 6734 59200 6790 60000
rect 7194 59200 7250 60000
rect 7746 59200 7802 60000
rect 8206 59200 8262 60000
rect 8666 59200 8722 60000
rect 9126 59200 9182 60000
rect 9586 59200 9642 60000
rect 10046 59200 10102 60000
rect 10506 59200 10562 60000
rect 10966 59200 11022 60000
rect 11518 59200 11574 60000
rect 11978 59200 12034 60000
rect 12438 59200 12494 60000
rect 12898 59200 12954 60000
rect 13358 59200 13414 60000
rect 13818 59200 13874 60000
rect 14278 59200 14334 60000
rect 14738 59200 14794 60000
rect 15290 59200 15346 60000
rect 15750 59200 15806 60000
rect 16210 59200 16266 60000
rect 16670 59200 16726 60000
rect 17130 59200 17186 60000
rect 17590 59200 17646 60000
rect 18050 59200 18106 60000
rect 18510 59200 18566 60000
rect 19062 59200 19118 60000
rect 19522 59200 19578 60000
rect 19982 59200 20038 60000
rect 20442 59200 20498 60000
rect 20902 59200 20958 60000
rect 21362 59200 21418 60000
rect 21822 59200 21878 60000
rect 22282 59200 22338 60000
rect 22834 59200 22890 60000
rect 23294 59200 23350 60000
rect 23754 59200 23810 60000
rect 24214 59200 24270 60000
rect 24674 59200 24730 60000
rect 25134 59200 25190 60000
rect 25594 59200 25650 60000
rect 26146 59200 26202 60000
rect 26606 59200 26662 60000
rect 27066 59200 27122 60000
rect 27526 59200 27582 60000
rect 27986 59200 28042 60000
rect 28446 59200 28502 60000
rect 28906 59200 28962 60000
rect 29366 59200 29422 60000
rect 29918 59200 29974 60000
rect 30378 59200 30434 60000
rect 30838 59200 30894 60000
rect 31298 59200 31354 60000
rect 31758 59200 31814 60000
rect 32218 59200 32274 60000
rect 32678 59200 32734 60000
rect 33138 59200 33194 60000
rect 33690 59200 33746 60000
rect 34150 59200 34206 60000
rect 34610 59200 34666 60000
rect 35070 59200 35126 60000
rect 35530 59200 35586 60000
rect 35990 59200 36046 60000
rect 36450 59200 36506 60000
rect 36910 59200 36966 60000
rect 37462 59200 37518 60000
rect 37922 59200 37978 60000
rect 38382 59200 38438 60000
rect 38842 59200 38898 60000
rect 39302 59200 39358 60000
rect 39762 59200 39818 60000
rect 40222 59200 40278 60000
rect 40682 59200 40738 60000
rect 41234 59200 41290 60000
rect 41694 59200 41750 60000
rect 42154 59200 42210 60000
rect 42614 59200 42670 60000
rect 43074 59200 43130 60000
rect 43534 59200 43590 60000
rect 43994 59200 44050 60000
rect 44454 59200 44510 60000
rect 45006 59200 45062 60000
rect 45466 59200 45522 60000
rect 45926 59200 45982 60000
rect 46386 59200 46442 60000
rect 46846 59200 46902 60000
rect 47306 59200 47362 60000
rect 47766 59200 47822 60000
rect 48226 59200 48282 60000
rect 48778 59200 48834 60000
rect 49238 59200 49294 60000
rect 49698 59200 49754 60000
rect 50158 59200 50214 60000
rect 50618 59200 50674 60000
rect 51078 59200 51134 60000
rect 51538 59200 51594 60000
rect 52090 59200 52146 60000
rect 52550 59200 52606 60000
rect 53010 59200 53066 60000
rect 53470 59200 53526 60000
rect 53930 59200 53986 60000
rect 54390 59200 54446 60000
rect 54850 59200 54906 60000
rect 55310 59200 55366 60000
rect 55862 59200 55918 60000
rect 56322 59200 56378 60000
rect 56782 59200 56838 60000
rect 57242 59200 57298 60000
rect 57702 59200 57758 60000
rect 58162 59200 58218 60000
rect 58622 59200 58678 60000
rect 59082 59200 59138 60000
rect 59634 59200 59690 60000
rect 60094 59200 60150 60000
rect 60554 59200 60610 60000
rect 61014 59200 61070 60000
rect 61474 59200 61530 60000
rect 61934 59200 61990 60000
rect 62394 59200 62450 60000
rect 62854 59200 62910 60000
rect 63406 59200 63462 60000
rect 63866 59200 63922 60000
rect 64326 59200 64382 60000
rect 64786 59200 64842 60000
rect 65246 59200 65302 60000
rect 65706 59200 65762 60000
rect 66166 59200 66222 60000
rect 66626 59200 66682 60000
rect 67178 59200 67234 60000
rect 67638 59200 67694 60000
rect 68098 59200 68154 60000
rect 68558 59200 68614 60000
rect 69018 59200 69074 60000
rect 69478 59200 69534 60000
rect 69938 59200 69994 60000
rect 70398 59200 70454 60000
rect 70950 59200 71006 60000
rect 71410 59200 71466 60000
rect 71870 59200 71926 60000
rect 72330 59200 72386 60000
rect 72790 59200 72846 60000
rect 73250 59200 73306 60000
rect 73710 59200 73766 60000
rect 74170 59200 74226 60000
rect 74722 59200 74778 60000
rect 75182 59200 75238 60000
rect 75642 59200 75698 60000
rect 76102 59200 76158 60000
rect 76562 59200 76618 60000
rect 77022 59200 77078 60000
rect 77482 59200 77538 60000
rect 78034 59200 78090 60000
rect 78494 59200 78550 60000
rect 78954 59200 79010 60000
rect 79414 59200 79470 60000
rect 79874 59200 79930 60000
rect 80334 59200 80390 60000
rect 80794 59200 80850 60000
rect 81254 59200 81310 60000
rect 81806 59200 81862 60000
rect 82266 59200 82322 60000
rect 82726 59200 82782 60000
rect 83186 59200 83242 60000
rect 83646 59200 83702 60000
rect 84106 59200 84162 60000
rect 84566 59200 84622 60000
rect 85026 59200 85082 60000
rect 85578 59200 85634 60000
rect 86038 59200 86094 60000
rect 86498 59200 86554 60000
rect 86958 59200 87014 60000
rect 87418 59200 87474 60000
rect 87878 59200 87934 60000
rect 88338 59200 88394 60000
rect 88798 59200 88854 60000
rect 89350 59200 89406 60000
rect 89810 59200 89866 60000
rect 90270 59200 90326 60000
rect 90730 59200 90786 60000
rect 91190 59200 91246 60000
rect 91650 59200 91706 60000
rect 92110 59200 92166 60000
rect 92570 59200 92626 60000
rect 93122 59200 93178 60000
rect 93582 59200 93638 60000
rect 94042 59200 94098 60000
rect 94502 59200 94558 60000
rect 94962 59200 95018 60000
rect 95422 59200 95478 60000
rect 95882 59200 95938 60000
rect 96342 59200 96398 60000
rect 96894 59200 96950 60000
rect 97354 59200 97410 60000
rect 97814 59200 97870 60000
rect 98274 59200 98330 60000
rect 98734 59200 98790 60000
rect 99194 59200 99250 60000
rect 99654 59200 99710 60000
<< obsm2 >>
rect 314 59144 606 59673
rect 774 59144 1066 59673
rect 1234 59144 1526 59673
rect 1694 59144 1986 59673
rect 2154 59144 2446 59673
rect 2614 59144 2906 59673
rect 3074 59144 3366 59673
rect 3534 59144 3918 59673
rect 4086 59144 4378 59673
rect 4546 59144 4838 59673
rect 5006 59144 5298 59673
rect 5466 59144 5758 59673
rect 5926 59144 6218 59673
rect 6386 59144 6678 59673
rect 6846 59144 7138 59673
rect 7306 59144 7690 59673
rect 7858 59144 8150 59673
rect 8318 59144 8610 59673
rect 8778 59144 9070 59673
rect 9238 59144 9530 59673
rect 9698 59144 9990 59673
rect 10158 59144 10450 59673
rect 10618 59144 10910 59673
rect 11078 59144 11462 59673
rect 11630 59144 11922 59673
rect 12090 59144 12382 59673
rect 12550 59144 12842 59673
rect 13010 59144 13302 59673
rect 13470 59144 13762 59673
rect 13930 59144 14222 59673
rect 14390 59144 14682 59673
rect 14850 59144 15234 59673
rect 15402 59144 15694 59673
rect 15862 59144 16154 59673
rect 16322 59144 16614 59673
rect 16782 59144 17074 59673
rect 17242 59144 17534 59673
rect 17702 59144 17994 59673
rect 18162 59144 18454 59673
rect 18622 59144 19006 59673
rect 19174 59144 19466 59673
rect 19634 59144 19926 59673
rect 20094 59144 20386 59673
rect 20554 59144 20846 59673
rect 21014 59144 21306 59673
rect 21474 59144 21766 59673
rect 21934 59144 22226 59673
rect 22394 59144 22778 59673
rect 22946 59144 23238 59673
rect 23406 59144 23698 59673
rect 23866 59144 24158 59673
rect 24326 59144 24618 59673
rect 24786 59144 25078 59673
rect 25246 59144 25538 59673
rect 25706 59144 26090 59673
rect 26258 59144 26550 59673
rect 26718 59144 27010 59673
rect 27178 59144 27470 59673
rect 27638 59144 27930 59673
rect 28098 59144 28390 59673
rect 28558 59144 28850 59673
rect 29018 59144 29310 59673
rect 29478 59144 29862 59673
rect 30030 59144 30322 59673
rect 30490 59144 30782 59673
rect 30950 59144 31242 59673
rect 31410 59144 31702 59673
rect 31870 59144 32162 59673
rect 32330 59144 32622 59673
rect 32790 59144 33082 59673
rect 33250 59144 33634 59673
rect 33802 59144 34094 59673
rect 34262 59144 34554 59673
rect 34722 59144 35014 59673
rect 35182 59144 35474 59673
rect 35642 59144 35934 59673
rect 36102 59144 36394 59673
rect 36562 59144 36854 59673
rect 37022 59144 37406 59673
rect 37574 59144 37866 59673
rect 38034 59144 38326 59673
rect 38494 59144 38786 59673
rect 38954 59144 39246 59673
rect 39414 59144 39706 59673
rect 39874 59144 40166 59673
rect 40334 59144 40626 59673
rect 40794 59144 41178 59673
rect 41346 59144 41638 59673
rect 41806 59144 42098 59673
rect 42266 59144 42558 59673
rect 42726 59144 43018 59673
rect 43186 59144 43478 59673
rect 43646 59144 43938 59673
rect 44106 59144 44398 59673
rect 44566 59144 44950 59673
rect 45118 59144 45410 59673
rect 45578 59144 45870 59673
rect 46038 59144 46330 59673
rect 46498 59144 46790 59673
rect 46958 59144 47250 59673
rect 47418 59144 47710 59673
rect 47878 59144 48170 59673
rect 48338 59144 48722 59673
rect 48890 59144 49182 59673
rect 49350 59144 49642 59673
rect 49810 59144 50102 59673
rect 50270 59144 50562 59673
rect 50730 59144 51022 59673
rect 51190 59144 51482 59673
rect 51650 59144 52034 59673
rect 52202 59144 52494 59673
rect 52662 59144 52954 59673
rect 53122 59144 53414 59673
rect 53582 59144 53874 59673
rect 54042 59144 54334 59673
rect 54502 59144 54794 59673
rect 54962 59144 55254 59673
rect 55422 59144 55806 59673
rect 55974 59144 56266 59673
rect 56434 59144 56726 59673
rect 56894 59144 57186 59673
rect 57354 59144 57646 59673
rect 57814 59144 58106 59673
rect 58274 59144 58566 59673
rect 58734 59144 59026 59673
rect 59194 59144 59578 59673
rect 59746 59144 60038 59673
rect 60206 59144 60498 59673
rect 60666 59144 60958 59673
rect 61126 59144 61418 59673
rect 61586 59144 61878 59673
rect 62046 59144 62338 59673
rect 62506 59144 62798 59673
rect 62966 59144 63350 59673
rect 63518 59144 63810 59673
rect 63978 59144 64270 59673
rect 64438 59144 64730 59673
rect 64898 59144 65190 59673
rect 65358 59144 65650 59673
rect 65818 59144 66110 59673
rect 66278 59144 66570 59673
rect 66738 59144 67122 59673
rect 67290 59144 67582 59673
rect 67750 59144 68042 59673
rect 68210 59144 68502 59673
rect 68670 59144 68962 59673
rect 69130 59144 69422 59673
rect 69590 59144 69882 59673
rect 70050 59144 70342 59673
rect 70510 59144 70894 59673
rect 71062 59144 71354 59673
rect 71522 59144 71814 59673
rect 71982 59144 72274 59673
rect 72442 59144 72734 59673
rect 72902 59144 73194 59673
rect 73362 59144 73654 59673
rect 73822 59144 74114 59673
rect 74282 59144 74666 59673
rect 74834 59144 75126 59673
rect 75294 59144 75586 59673
rect 75754 59144 76046 59673
rect 76214 59144 76506 59673
rect 76674 59144 76966 59673
rect 77134 59144 77426 59673
rect 77594 59144 77978 59673
rect 78146 59144 78438 59673
rect 78606 59144 78898 59673
rect 79066 59144 79358 59673
rect 79526 59144 79818 59673
rect 79986 59144 80278 59673
rect 80446 59144 80738 59673
rect 80906 59144 81198 59673
rect 81366 59144 81750 59673
rect 81918 59144 82210 59673
rect 82378 59144 82670 59673
rect 82838 59144 83130 59673
rect 83298 59144 83590 59673
rect 83758 59144 84050 59673
rect 84218 59144 84510 59673
rect 84678 59144 84970 59673
rect 85138 59144 85522 59673
rect 85690 59144 85982 59673
rect 86150 59144 86442 59673
rect 86610 59144 86902 59673
rect 87070 59144 87362 59673
rect 87530 59144 87822 59673
rect 87990 59144 88282 59673
rect 88450 59144 88742 59673
rect 88910 59144 89294 59673
rect 89462 59144 89754 59673
rect 89922 59144 90214 59673
rect 90382 59144 90674 59673
rect 90842 59144 91134 59673
rect 91302 59144 91594 59673
rect 91762 59144 92054 59673
rect 92222 59144 92514 59673
rect 92682 59144 93066 59673
rect 93234 59144 93526 59673
rect 93694 59144 93986 59673
rect 94154 59144 94446 59673
rect 94614 59144 94906 59673
rect 95074 59144 95366 59673
rect 95534 59144 95826 59673
rect 95994 59144 96286 59673
rect 96454 59144 96838 59673
rect 97006 59144 97298 59673
rect 97466 59144 97758 59673
rect 97926 59144 98218 59673
rect 98386 59144 98678 59673
rect 98846 59144 99138 59673
rect 99306 59144 99598 59673
rect 204 303 99708 59144
<< metal3 >>
rect 0 59576 800 59696
rect 0 59032 800 59152
rect 0 58488 800 58608
rect 0 57944 800 58064
rect 0 57400 800 57520
rect 0 56856 800 56976
rect 0 56312 800 56432
rect 0 55768 800 55888
rect 0 55224 800 55344
rect 0 54680 800 54800
rect 0 54136 800 54256
rect 0 53592 800 53712
rect 0 52912 800 53032
rect 0 52368 800 52488
rect 0 51824 800 51944
rect 0 51280 800 51400
rect 0 50736 800 50856
rect 0 50192 800 50312
rect 0 49648 800 49768
rect 0 49104 800 49224
rect 0 48560 800 48680
rect 0 48016 800 48136
rect 0 47472 800 47592
rect 0 46928 800 47048
rect 0 46248 800 46368
rect 0 45704 800 45824
rect 0 45160 800 45280
rect 0 44616 800 44736
rect 0 44072 800 44192
rect 0 43528 800 43648
rect 0 42984 800 43104
rect 0 42440 800 42560
rect 0 41896 800 42016
rect 0 41352 800 41472
rect 0 40808 800 40928
rect 0 40264 800 40384
rect 0 39584 800 39704
rect 0 39040 800 39160
rect 0 38496 800 38616
rect 0 37952 800 38072
rect 0 37408 800 37528
rect 0 36864 800 36984
rect 0 36320 800 36440
rect 0 35776 800 35896
rect 0 35232 800 35352
rect 0 34688 800 34808
rect 0 34144 800 34264
rect 0 33600 800 33720
rect 0 32920 800 33040
rect 0 32376 800 32496
rect 0 31832 800 31952
rect 0 31288 800 31408
rect 0 30744 800 30864
rect 0 30200 800 30320
rect 0 29656 800 29776
rect 0 29112 800 29232
rect 0 28568 800 28688
rect 0 28024 800 28144
rect 0 27480 800 27600
rect 0 26936 800 27056
rect 0 26256 800 26376
rect 0 25712 800 25832
rect 0 25168 800 25288
rect 0 24624 800 24744
rect 0 24080 800 24200
rect 0 23536 800 23656
rect 0 22992 800 23112
rect 0 22448 800 22568
rect 0 21904 800 22024
rect 0 21360 800 21480
rect 0 20816 800 20936
rect 0 20272 800 20392
rect 0 19592 800 19712
rect 0 19048 800 19168
rect 0 18504 800 18624
rect 0 17960 800 18080
rect 0 17416 800 17536
rect 0 16872 800 16992
rect 0 16328 800 16448
rect 0 15784 800 15904
rect 0 15240 800 15360
rect 0 14696 800 14816
rect 0 14152 800 14272
rect 0 13608 800 13728
rect 0 12928 800 13048
rect 0 12384 800 12504
rect 0 11840 800 11960
rect 0 11296 800 11416
rect 0 10752 800 10872
rect 0 10208 800 10328
rect 0 9664 800 9784
rect 0 9120 800 9240
rect 0 8576 800 8696
rect 0 8032 800 8152
rect 0 7488 800 7608
rect 0 6944 800 7064
rect 0 6264 800 6384
rect 0 5720 800 5840
rect 0 5176 800 5296
rect 0 4632 800 4752
rect 0 4088 800 4208
rect 0 3544 800 3664
rect 0 3000 800 3120
rect 0 2456 800 2576
rect 0 1912 800 2032
rect 0 1368 800 1488
rect 0 824 800 944
rect 0 280 800 400
<< obsm3 >>
rect 880 59496 97967 59669
rect 800 59232 97967 59496
rect 880 58952 97967 59232
rect 800 58688 97967 58952
rect 880 58408 97967 58688
rect 800 58144 97967 58408
rect 880 57864 97967 58144
rect 800 57600 97967 57864
rect 880 57320 97967 57600
rect 800 57056 97967 57320
rect 880 56776 97967 57056
rect 800 56512 97967 56776
rect 880 56232 97967 56512
rect 800 55968 97967 56232
rect 880 55688 97967 55968
rect 800 55424 97967 55688
rect 880 55144 97967 55424
rect 800 54880 97967 55144
rect 880 54600 97967 54880
rect 800 54336 97967 54600
rect 880 54056 97967 54336
rect 800 53792 97967 54056
rect 880 53512 97967 53792
rect 800 53112 97967 53512
rect 880 52832 97967 53112
rect 800 52568 97967 52832
rect 880 52288 97967 52568
rect 800 52024 97967 52288
rect 880 51744 97967 52024
rect 800 51480 97967 51744
rect 880 51200 97967 51480
rect 800 50936 97967 51200
rect 880 50656 97967 50936
rect 800 50392 97967 50656
rect 880 50112 97967 50392
rect 800 49848 97967 50112
rect 880 49568 97967 49848
rect 800 49304 97967 49568
rect 880 49024 97967 49304
rect 800 48760 97967 49024
rect 880 48480 97967 48760
rect 800 48216 97967 48480
rect 880 47936 97967 48216
rect 800 47672 97967 47936
rect 880 47392 97967 47672
rect 800 47128 97967 47392
rect 880 46848 97967 47128
rect 800 46448 97967 46848
rect 880 46168 97967 46448
rect 800 45904 97967 46168
rect 880 45624 97967 45904
rect 800 45360 97967 45624
rect 880 45080 97967 45360
rect 800 44816 97967 45080
rect 880 44536 97967 44816
rect 800 44272 97967 44536
rect 880 43992 97967 44272
rect 800 43728 97967 43992
rect 880 43448 97967 43728
rect 800 43184 97967 43448
rect 880 42904 97967 43184
rect 800 42640 97967 42904
rect 880 42360 97967 42640
rect 800 42096 97967 42360
rect 880 41816 97967 42096
rect 800 41552 97967 41816
rect 880 41272 97967 41552
rect 800 41008 97967 41272
rect 880 40728 97967 41008
rect 800 40464 97967 40728
rect 880 40184 97967 40464
rect 800 39784 97967 40184
rect 880 39504 97967 39784
rect 800 39240 97967 39504
rect 880 38960 97967 39240
rect 800 38696 97967 38960
rect 880 38416 97967 38696
rect 800 38152 97967 38416
rect 880 37872 97967 38152
rect 800 37608 97967 37872
rect 880 37328 97967 37608
rect 800 37064 97967 37328
rect 880 36784 97967 37064
rect 800 36520 97967 36784
rect 880 36240 97967 36520
rect 800 35976 97967 36240
rect 880 35696 97967 35976
rect 800 35432 97967 35696
rect 880 35152 97967 35432
rect 800 34888 97967 35152
rect 880 34608 97967 34888
rect 800 34344 97967 34608
rect 880 34064 97967 34344
rect 800 33800 97967 34064
rect 880 33520 97967 33800
rect 800 33120 97967 33520
rect 880 32840 97967 33120
rect 800 32576 97967 32840
rect 880 32296 97967 32576
rect 800 32032 97967 32296
rect 880 31752 97967 32032
rect 800 31488 97967 31752
rect 880 31208 97967 31488
rect 800 30944 97967 31208
rect 880 30664 97967 30944
rect 800 30400 97967 30664
rect 880 30120 97967 30400
rect 800 29856 97967 30120
rect 880 29576 97967 29856
rect 800 29312 97967 29576
rect 880 29032 97967 29312
rect 800 28768 97967 29032
rect 880 28488 97967 28768
rect 800 28224 97967 28488
rect 880 27944 97967 28224
rect 800 27680 97967 27944
rect 880 27400 97967 27680
rect 800 27136 97967 27400
rect 880 26856 97967 27136
rect 800 26456 97967 26856
rect 880 26176 97967 26456
rect 800 25912 97967 26176
rect 880 25632 97967 25912
rect 800 25368 97967 25632
rect 880 25088 97967 25368
rect 800 24824 97967 25088
rect 880 24544 97967 24824
rect 800 24280 97967 24544
rect 880 24000 97967 24280
rect 800 23736 97967 24000
rect 880 23456 97967 23736
rect 800 23192 97967 23456
rect 880 22912 97967 23192
rect 800 22648 97967 22912
rect 880 22368 97967 22648
rect 800 22104 97967 22368
rect 880 21824 97967 22104
rect 800 21560 97967 21824
rect 880 21280 97967 21560
rect 800 21016 97967 21280
rect 880 20736 97967 21016
rect 800 20472 97967 20736
rect 880 20192 97967 20472
rect 800 19792 97967 20192
rect 880 19512 97967 19792
rect 800 19248 97967 19512
rect 880 18968 97967 19248
rect 800 18704 97967 18968
rect 880 18424 97967 18704
rect 800 18160 97967 18424
rect 880 17880 97967 18160
rect 800 17616 97967 17880
rect 880 17336 97967 17616
rect 800 17072 97967 17336
rect 880 16792 97967 17072
rect 800 16528 97967 16792
rect 880 16248 97967 16528
rect 800 15984 97967 16248
rect 880 15704 97967 15984
rect 800 15440 97967 15704
rect 880 15160 97967 15440
rect 800 14896 97967 15160
rect 880 14616 97967 14896
rect 800 14352 97967 14616
rect 880 14072 97967 14352
rect 800 13808 97967 14072
rect 880 13528 97967 13808
rect 800 13128 97967 13528
rect 880 12848 97967 13128
rect 800 12584 97967 12848
rect 880 12304 97967 12584
rect 800 12040 97967 12304
rect 880 11760 97967 12040
rect 800 11496 97967 11760
rect 880 11216 97967 11496
rect 800 10952 97967 11216
rect 880 10672 97967 10952
rect 800 10408 97967 10672
rect 880 10128 97967 10408
rect 800 9864 97967 10128
rect 880 9584 97967 9864
rect 800 9320 97967 9584
rect 880 9040 97967 9320
rect 800 8776 97967 9040
rect 880 8496 97967 8776
rect 800 8232 97967 8496
rect 880 7952 97967 8232
rect 800 7688 97967 7952
rect 880 7408 97967 7688
rect 800 7144 97967 7408
rect 880 6864 97967 7144
rect 800 6464 97967 6864
rect 880 6184 97967 6464
rect 800 5920 97967 6184
rect 880 5640 97967 5920
rect 800 5376 97967 5640
rect 880 5096 97967 5376
rect 800 4832 97967 5096
rect 880 4552 97967 4832
rect 800 4288 97967 4552
rect 880 4008 97967 4288
rect 800 3744 97967 4008
rect 880 3464 97967 3744
rect 800 3200 97967 3464
rect 880 2920 97967 3200
rect 800 2656 97967 2920
rect 880 2376 97967 2656
rect 800 2112 97967 2376
rect 880 1832 97967 2112
rect 800 1568 97967 1832
rect 880 1288 97967 1568
rect 800 1024 97967 1288
rect 880 744 97967 1024
rect 800 480 97967 744
rect 880 307 97967 480
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
rect 65648 2128 65968 57712
rect 81008 2128 81328 57712
rect 96368 2128 96688 57712
<< obsm4 >>
rect 1531 57792 77773 58309
rect 1531 3163 4128 57792
rect 4608 3163 19488 57792
rect 19968 3163 34848 57792
rect 35328 3163 50208 57792
rect 50688 3163 65568 57792
rect 66048 3163 77773 57792
<< labels >>
rlabel metal3 s 0 280 800 400 6 CLK
port 1 nsew signal input
rlabel metal3 s 0 824 800 944 6 RST_N
port 2 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 cpu_ack_o
port 3 nsew signal output
rlabel metal3 s 0 4632 800 4752 6 cpu_adr_i[0]
port 4 nsew signal input
rlabel metal3 s 0 23536 800 23656 6 cpu_adr_i[10]
port 5 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 cpu_adr_i[11]
port 6 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 cpu_adr_i[12]
port 7 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 cpu_adr_i[13]
port 8 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 cpu_adr_i[14]
port 9 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 cpu_adr_i[15]
port 10 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 cpu_adr_i[16]
port 11 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 cpu_adr_i[17]
port 12 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 cpu_adr_i[18]
port 13 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 cpu_adr_i[19]
port 14 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 cpu_adr_i[1]
port 15 nsew signal input
rlabel metal3 s 0 40264 800 40384 6 cpu_adr_i[20]
port 16 nsew signal input
rlabel metal3 s 0 41896 800 42016 6 cpu_adr_i[21]
port 17 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 cpu_adr_i[22]
port 18 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 cpu_adr_i[23]
port 19 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 cpu_adr_i[24]
port 20 nsew signal input
rlabel metal3 s 0 48560 800 48680 6 cpu_adr_i[25]
port 21 nsew signal input
rlabel metal3 s 0 50192 800 50312 6 cpu_adr_i[26]
port 22 nsew signal input
rlabel metal3 s 0 51824 800 51944 6 cpu_adr_i[27]
port 23 nsew signal input
rlabel metal3 s 0 53592 800 53712 6 cpu_adr_i[28]
port 24 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 cpu_adr_i[29]
port 25 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 cpu_adr_i[2]
port 26 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 cpu_adr_i[30]
port 27 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 cpu_adr_i[31]
port 28 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 cpu_adr_i[3]
port 29 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 cpu_adr_i[4]
port 30 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 cpu_adr_i[5]
port 31 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 cpu_adr_i[6]
port 32 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 cpu_adr_i[7]
port 33 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 cpu_adr_i[8]
port 34 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 cpu_adr_i[9]
port 35 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 cpu_cyc_i
port 36 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 cpu_dat_i[0]
port 37 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 cpu_dat_i[10]
port 38 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 cpu_dat_i[11]
port 39 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 cpu_dat_i[12]
port 40 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 cpu_dat_i[13]
port 41 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 cpu_dat_i[14]
port 42 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 cpu_dat_i[15]
port 43 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 cpu_dat_i[16]
port 44 nsew signal input
rlabel metal3 s 0 35776 800 35896 6 cpu_dat_i[17]
port 45 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 cpu_dat_i[18]
port 46 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 cpu_dat_i[19]
port 47 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 cpu_dat_i[1]
port 48 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 cpu_dat_i[20]
port 49 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 cpu_dat_i[21]
port 50 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 cpu_dat_i[22]
port 51 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 cpu_dat_i[23]
port 52 nsew signal input
rlabel metal3 s 0 47472 800 47592 6 cpu_dat_i[24]
port 53 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 cpu_dat_i[25]
port 54 nsew signal input
rlabel metal3 s 0 50736 800 50856 6 cpu_dat_i[26]
port 55 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 cpu_dat_i[27]
port 56 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 cpu_dat_i[28]
port 57 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 cpu_dat_i[29]
port 58 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 cpu_dat_i[2]
port 59 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 cpu_dat_i[30]
port 60 nsew signal input
rlabel metal3 s 0 59032 800 59152 6 cpu_dat_i[31]
port 61 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 cpu_dat_i[3]
port 62 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 cpu_dat_i[4]
port 63 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 cpu_dat_i[5]
port 64 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 cpu_dat_i[6]
port 65 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 cpu_dat_i[7]
port 66 nsew signal input
rlabel metal3 s 0 20816 800 20936 6 cpu_dat_i[8]
port 67 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 cpu_dat_i[9]
port 68 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 cpu_dat_o[0]
port 69 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 cpu_dat_o[10]
port 70 nsew signal output
rlabel metal3 s 0 26256 800 26376 6 cpu_dat_o[11]
port 71 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 cpu_dat_o[12]
port 72 nsew signal output
rlabel metal3 s 0 29656 800 29776 6 cpu_dat_o[13]
port 73 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 cpu_dat_o[14]
port 74 nsew signal output
rlabel metal3 s 0 32920 800 33040 6 cpu_dat_o[15]
port 75 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 cpu_dat_o[16]
port 76 nsew signal output
rlabel metal3 s 0 36320 800 36440 6 cpu_dat_o[17]
port 77 nsew signal output
rlabel metal3 s 0 37952 800 38072 6 cpu_dat_o[18]
port 78 nsew signal output
rlabel metal3 s 0 39584 800 39704 6 cpu_dat_o[19]
port 79 nsew signal output
rlabel metal3 s 0 8032 800 8152 6 cpu_dat_o[1]
port 80 nsew signal output
rlabel metal3 s 0 41352 800 41472 6 cpu_dat_o[20]
port 81 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 cpu_dat_o[21]
port 82 nsew signal output
rlabel metal3 s 0 44616 800 44736 6 cpu_dat_o[22]
port 83 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 cpu_dat_o[23]
port 84 nsew signal output
rlabel metal3 s 0 48016 800 48136 6 cpu_dat_o[24]
port 85 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 cpu_dat_o[25]
port 86 nsew signal output
rlabel metal3 s 0 51280 800 51400 6 cpu_dat_o[26]
port 87 nsew signal output
rlabel metal3 s 0 52912 800 53032 6 cpu_dat_o[27]
port 88 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 cpu_dat_o[28]
port 89 nsew signal output
rlabel metal3 s 0 56312 800 56432 6 cpu_dat_o[29]
port 90 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 cpu_dat_o[2]
port 91 nsew signal output
rlabel metal3 s 0 57944 800 58064 6 cpu_dat_o[30]
port 92 nsew signal output
rlabel metal3 s 0 59576 800 59696 6 cpu_dat_o[31]
port 93 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 cpu_dat_o[3]
port 94 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 cpu_dat_o[4]
port 95 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 cpu_dat_o[5]
port 96 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 cpu_dat_o[6]
port 97 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 cpu_dat_o[7]
port 98 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 cpu_dat_o[8]
port 99 nsew signal output
rlabel metal3 s 0 22992 800 23112 6 cpu_dat_o[9]
port 100 nsew signal output
rlabel metal3 s 0 2456 800 2576 6 cpu_err_o
port 101 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 cpu_rty_o
port 102 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 cpu_sel_i[0]
port 103 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 cpu_sel_i[1]
port 104 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 cpu_sel_i[2]
port 105 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 cpu_sel_i[3]
port 106 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 cpu_stb_i
port 107 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 cpu_we_i
port 108 nsew signal input
rlabel metal2 s 50158 59200 50214 60000 6 gpio_ack_i
port 109 nsew signal input
rlabel metal2 s 53010 59200 53066 60000 6 gpio_adr_o[0]
port 110 nsew signal output
rlabel metal2 s 69018 59200 69074 60000 6 gpio_adr_o[10]
port 111 nsew signal output
rlabel metal2 s 70398 59200 70454 60000 6 gpio_adr_o[11]
port 112 nsew signal output
rlabel metal2 s 71870 59200 71926 60000 6 gpio_adr_o[12]
port 113 nsew signal output
rlabel metal2 s 73250 59200 73306 60000 6 gpio_adr_o[13]
port 114 nsew signal output
rlabel metal2 s 74722 59200 74778 60000 6 gpio_adr_o[14]
port 115 nsew signal output
rlabel metal2 s 76102 59200 76158 60000 6 gpio_adr_o[15]
port 116 nsew signal output
rlabel metal2 s 77482 59200 77538 60000 6 gpio_adr_o[16]
port 117 nsew signal output
rlabel metal2 s 78954 59200 79010 60000 6 gpio_adr_o[17]
port 118 nsew signal output
rlabel metal2 s 80334 59200 80390 60000 6 gpio_adr_o[18]
port 119 nsew signal output
rlabel metal2 s 81806 59200 81862 60000 6 gpio_adr_o[19]
port 120 nsew signal output
rlabel metal2 s 54850 59200 54906 60000 6 gpio_adr_o[1]
port 121 nsew signal output
rlabel metal2 s 83186 59200 83242 60000 6 gpio_adr_o[20]
port 122 nsew signal output
rlabel metal2 s 84566 59200 84622 60000 6 gpio_adr_o[21]
port 123 nsew signal output
rlabel metal2 s 86038 59200 86094 60000 6 gpio_adr_o[22]
port 124 nsew signal output
rlabel metal2 s 87418 59200 87474 60000 6 gpio_adr_o[23]
port 125 nsew signal output
rlabel metal2 s 88798 59200 88854 60000 6 gpio_adr_o[24]
port 126 nsew signal output
rlabel metal2 s 90270 59200 90326 60000 6 gpio_adr_o[25]
port 127 nsew signal output
rlabel metal2 s 91650 59200 91706 60000 6 gpio_adr_o[26]
port 128 nsew signal output
rlabel metal2 s 93122 59200 93178 60000 6 gpio_adr_o[27]
port 129 nsew signal output
rlabel metal2 s 94502 59200 94558 60000 6 gpio_adr_o[28]
port 130 nsew signal output
rlabel metal2 s 95882 59200 95938 60000 6 gpio_adr_o[29]
port 131 nsew signal output
rlabel metal2 s 56782 59200 56838 60000 6 gpio_adr_o[2]
port 132 nsew signal output
rlabel metal2 s 97354 59200 97410 60000 6 gpio_adr_o[30]
port 133 nsew signal output
rlabel metal2 s 98734 59200 98790 60000 6 gpio_adr_o[31]
port 134 nsew signal output
rlabel metal2 s 58622 59200 58678 60000 6 gpio_adr_o[3]
port 135 nsew signal output
rlabel metal2 s 60554 59200 60610 60000 6 gpio_adr_o[4]
port 136 nsew signal output
rlabel metal2 s 61934 59200 61990 60000 6 gpio_adr_o[5]
port 137 nsew signal output
rlabel metal2 s 63406 59200 63462 60000 6 gpio_adr_o[6]
port 138 nsew signal output
rlabel metal2 s 64786 59200 64842 60000 6 gpio_adr_o[7]
port 139 nsew signal output
rlabel metal2 s 66166 59200 66222 60000 6 gpio_adr_o[8]
port 140 nsew signal output
rlabel metal2 s 67638 59200 67694 60000 6 gpio_adr_o[9]
port 141 nsew signal output
rlabel metal2 s 50618 59200 50674 60000 6 gpio_cyc_o
port 142 nsew signal output
rlabel metal2 s 53470 59200 53526 60000 6 gpio_dat_i[0]
port 143 nsew signal input
rlabel metal2 s 69478 59200 69534 60000 6 gpio_dat_i[10]
port 144 nsew signal input
rlabel metal2 s 70950 59200 71006 60000 6 gpio_dat_i[11]
port 145 nsew signal input
rlabel metal2 s 72330 59200 72386 60000 6 gpio_dat_i[12]
port 146 nsew signal input
rlabel metal2 s 73710 59200 73766 60000 6 gpio_dat_i[13]
port 147 nsew signal input
rlabel metal2 s 75182 59200 75238 60000 6 gpio_dat_i[14]
port 148 nsew signal input
rlabel metal2 s 76562 59200 76618 60000 6 gpio_dat_i[15]
port 149 nsew signal input
rlabel metal2 s 78034 59200 78090 60000 6 gpio_dat_i[16]
port 150 nsew signal input
rlabel metal2 s 79414 59200 79470 60000 6 gpio_dat_i[17]
port 151 nsew signal input
rlabel metal2 s 80794 59200 80850 60000 6 gpio_dat_i[18]
port 152 nsew signal input
rlabel metal2 s 82266 59200 82322 60000 6 gpio_dat_i[19]
port 153 nsew signal input
rlabel metal2 s 55310 59200 55366 60000 6 gpio_dat_i[1]
port 154 nsew signal input
rlabel metal2 s 83646 59200 83702 60000 6 gpio_dat_i[20]
port 155 nsew signal input
rlabel metal2 s 85026 59200 85082 60000 6 gpio_dat_i[21]
port 156 nsew signal input
rlabel metal2 s 86498 59200 86554 60000 6 gpio_dat_i[22]
port 157 nsew signal input
rlabel metal2 s 87878 59200 87934 60000 6 gpio_dat_i[23]
port 158 nsew signal input
rlabel metal2 s 89350 59200 89406 60000 6 gpio_dat_i[24]
port 159 nsew signal input
rlabel metal2 s 90730 59200 90786 60000 6 gpio_dat_i[25]
port 160 nsew signal input
rlabel metal2 s 92110 59200 92166 60000 6 gpio_dat_i[26]
port 161 nsew signal input
rlabel metal2 s 93582 59200 93638 60000 6 gpio_dat_i[27]
port 162 nsew signal input
rlabel metal2 s 94962 59200 95018 60000 6 gpio_dat_i[28]
port 163 nsew signal input
rlabel metal2 s 96342 59200 96398 60000 6 gpio_dat_i[29]
port 164 nsew signal input
rlabel metal2 s 57242 59200 57298 60000 6 gpio_dat_i[2]
port 165 nsew signal input
rlabel metal2 s 97814 59200 97870 60000 6 gpio_dat_i[30]
port 166 nsew signal input
rlabel metal2 s 99194 59200 99250 60000 6 gpio_dat_i[31]
port 167 nsew signal input
rlabel metal2 s 59082 59200 59138 60000 6 gpio_dat_i[3]
port 168 nsew signal input
rlabel metal2 s 61014 59200 61070 60000 6 gpio_dat_i[4]
port 169 nsew signal input
rlabel metal2 s 62394 59200 62450 60000 6 gpio_dat_i[5]
port 170 nsew signal input
rlabel metal2 s 63866 59200 63922 60000 6 gpio_dat_i[6]
port 171 nsew signal input
rlabel metal2 s 65246 59200 65302 60000 6 gpio_dat_i[7]
port 172 nsew signal input
rlabel metal2 s 66626 59200 66682 60000 6 gpio_dat_i[8]
port 173 nsew signal input
rlabel metal2 s 68098 59200 68154 60000 6 gpio_dat_i[9]
port 174 nsew signal input
rlabel metal2 s 53930 59200 53986 60000 6 gpio_dat_o[0]
port 175 nsew signal output
rlabel metal2 s 69938 59200 69994 60000 6 gpio_dat_o[10]
port 176 nsew signal output
rlabel metal2 s 71410 59200 71466 60000 6 gpio_dat_o[11]
port 177 nsew signal output
rlabel metal2 s 72790 59200 72846 60000 6 gpio_dat_o[12]
port 178 nsew signal output
rlabel metal2 s 74170 59200 74226 60000 6 gpio_dat_o[13]
port 179 nsew signal output
rlabel metal2 s 75642 59200 75698 60000 6 gpio_dat_o[14]
port 180 nsew signal output
rlabel metal2 s 77022 59200 77078 60000 6 gpio_dat_o[15]
port 181 nsew signal output
rlabel metal2 s 78494 59200 78550 60000 6 gpio_dat_o[16]
port 182 nsew signal output
rlabel metal2 s 79874 59200 79930 60000 6 gpio_dat_o[17]
port 183 nsew signal output
rlabel metal2 s 81254 59200 81310 60000 6 gpio_dat_o[18]
port 184 nsew signal output
rlabel metal2 s 82726 59200 82782 60000 6 gpio_dat_o[19]
port 185 nsew signal output
rlabel metal2 s 55862 59200 55918 60000 6 gpio_dat_o[1]
port 186 nsew signal output
rlabel metal2 s 84106 59200 84162 60000 6 gpio_dat_o[20]
port 187 nsew signal output
rlabel metal2 s 85578 59200 85634 60000 6 gpio_dat_o[21]
port 188 nsew signal output
rlabel metal2 s 86958 59200 87014 60000 6 gpio_dat_o[22]
port 189 nsew signal output
rlabel metal2 s 88338 59200 88394 60000 6 gpio_dat_o[23]
port 190 nsew signal output
rlabel metal2 s 89810 59200 89866 60000 6 gpio_dat_o[24]
port 191 nsew signal output
rlabel metal2 s 91190 59200 91246 60000 6 gpio_dat_o[25]
port 192 nsew signal output
rlabel metal2 s 92570 59200 92626 60000 6 gpio_dat_o[26]
port 193 nsew signal output
rlabel metal2 s 94042 59200 94098 60000 6 gpio_dat_o[27]
port 194 nsew signal output
rlabel metal2 s 95422 59200 95478 60000 6 gpio_dat_o[28]
port 195 nsew signal output
rlabel metal2 s 96894 59200 96950 60000 6 gpio_dat_o[29]
port 196 nsew signal output
rlabel metal2 s 57702 59200 57758 60000 6 gpio_dat_o[2]
port 197 nsew signal output
rlabel metal2 s 98274 59200 98330 60000 6 gpio_dat_o[30]
port 198 nsew signal output
rlabel metal2 s 99654 59200 99710 60000 6 gpio_dat_o[31]
port 199 nsew signal output
rlabel metal2 s 59634 59200 59690 60000 6 gpio_dat_o[3]
port 200 nsew signal output
rlabel metal2 s 61474 59200 61530 60000 6 gpio_dat_o[4]
port 201 nsew signal output
rlabel metal2 s 62854 59200 62910 60000 6 gpio_dat_o[5]
port 202 nsew signal output
rlabel metal2 s 64326 59200 64382 60000 6 gpio_dat_o[6]
port 203 nsew signal output
rlabel metal2 s 65706 59200 65762 60000 6 gpio_dat_o[7]
port 204 nsew signal output
rlabel metal2 s 67178 59200 67234 60000 6 gpio_dat_o[8]
port 205 nsew signal output
rlabel metal2 s 68558 59200 68614 60000 6 gpio_dat_o[9]
port 206 nsew signal output
rlabel metal2 s 51078 59200 51134 60000 6 gpio_err_i
port 207 nsew signal input
rlabel metal2 s 51538 59200 51594 60000 6 gpio_rty_i
port 208 nsew signal input
rlabel metal2 s 54390 59200 54446 60000 6 gpio_sel_o[0]
port 209 nsew signal output
rlabel metal2 s 56322 59200 56378 60000 6 gpio_sel_o[1]
port 210 nsew signal output
rlabel metal2 s 58162 59200 58218 60000 6 gpio_sel_o[2]
port 211 nsew signal output
rlabel metal2 s 60094 59200 60150 60000 6 gpio_sel_o[3]
port 212 nsew signal output
rlabel metal2 s 52090 59200 52146 60000 6 gpio_stb_o
port 213 nsew signal output
rlabel metal2 s 52550 59200 52606 60000 6 gpio_we_o
port 214 nsew signal output
rlabel metal2 s 202 59200 258 60000 6 spi_ack_i
port 215 nsew signal input
rlabel metal2 s 2962 59200 3018 60000 6 spi_adr_o[0]
port 216 nsew signal output
rlabel metal2 s 19062 59200 19118 60000 6 spi_adr_o[10]
port 217 nsew signal output
rlabel metal2 s 20442 59200 20498 60000 6 spi_adr_o[11]
port 218 nsew signal output
rlabel metal2 s 21822 59200 21878 60000 6 spi_adr_o[12]
port 219 nsew signal output
rlabel metal2 s 23294 59200 23350 60000 6 spi_adr_o[13]
port 220 nsew signal output
rlabel metal2 s 24674 59200 24730 60000 6 spi_adr_o[14]
port 221 nsew signal output
rlabel metal2 s 26146 59200 26202 60000 6 spi_adr_o[15]
port 222 nsew signal output
rlabel metal2 s 27526 59200 27582 60000 6 spi_adr_o[16]
port 223 nsew signal output
rlabel metal2 s 28906 59200 28962 60000 6 spi_adr_o[17]
port 224 nsew signal output
rlabel metal2 s 30378 59200 30434 60000 6 spi_adr_o[18]
port 225 nsew signal output
rlabel metal2 s 31758 59200 31814 60000 6 spi_adr_o[19]
port 226 nsew signal output
rlabel metal2 s 4894 59200 4950 60000 6 spi_adr_o[1]
port 227 nsew signal output
rlabel metal2 s 33138 59200 33194 60000 6 spi_adr_o[20]
port 228 nsew signal output
rlabel metal2 s 34610 59200 34666 60000 6 spi_adr_o[21]
port 229 nsew signal output
rlabel metal2 s 35990 59200 36046 60000 6 spi_adr_o[22]
port 230 nsew signal output
rlabel metal2 s 37462 59200 37518 60000 6 spi_adr_o[23]
port 231 nsew signal output
rlabel metal2 s 38842 59200 38898 60000 6 spi_adr_o[24]
port 232 nsew signal output
rlabel metal2 s 40222 59200 40278 60000 6 spi_adr_o[25]
port 233 nsew signal output
rlabel metal2 s 41694 59200 41750 60000 6 spi_adr_o[26]
port 234 nsew signal output
rlabel metal2 s 43074 59200 43130 60000 6 spi_adr_o[27]
port 235 nsew signal output
rlabel metal2 s 44454 59200 44510 60000 6 spi_adr_o[28]
port 236 nsew signal output
rlabel metal2 s 45926 59200 45982 60000 6 spi_adr_o[29]
port 237 nsew signal output
rlabel metal2 s 6734 59200 6790 60000 6 spi_adr_o[2]
port 238 nsew signal output
rlabel metal2 s 47306 59200 47362 60000 6 spi_adr_o[30]
port 239 nsew signal output
rlabel metal2 s 48778 59200 48834 60000 6 spi_adr_o[31]
port 240 nsew signal output
rlabel metal2 s 8666 59200 8722 60000 6 spi_adr_o[3]
port 241 nsew signal output
rlabel metal2 s 10506 59200 10562 60000 6 spi_adr_o[4]
port 242 nsew signal output
rlabel metal2 s 11978 59200 12034 60000 6 spi_adr_o[5]
port 243 nsew signal output
rlabel metal2 s 13358 59200 13414 60000 6 spi_adr_o[6]
port 244 nsew signal output
rlabel metal2 s 14738 59200 14794 60000 6 spi_adr_o[7]
port 245 nsew signal output
rlabel metal2 s 16210 59200 16266 60000 6 spi_adr_o[8]
port 246 nsew signal output
rlabel metal2 s 17590 59200 17646 60000 6 spi_adr_o[9]
port 247 nsew signal output
rlabel metal2 s 662 59200 718 60000 6 spi_cyc_o
port 248 nsew signal output
rlabel metal2 s 3422 59200 3478 60000 6 spi_dat_i[0]
port 249 nsew signal input
rlabel metal2 s 19522 59200 19578 60000 6 spi_dat_i[10]
port 250 nsew signal input
rlabel metal2 s 20902 59200 20958 60000 6 spi_dat_i[11]
port 251 nsew signal input
rlabel metal2 s 22282 59200 22338 60000 6 spi_dat_i[12]
port 252 nsew signal input
rlabel metal2 s 23754 59200 23810 60000 6 spi_dat_i[13]
port 253 nsew signal input
rlabel metal2 s 25134 59200 25190 60000 6 spi_dat_i[14]
port 254 nsew signal input
rlabel metal2 s 26606 59200 26662 60000 6 spi_dat_i[15]
port 255 nsew signal input
rlabel metal2 s 27986 59200 28042 60000 6 spi_dat_i[16]
port 256 nsew signal input
rlabel metal2 s 29366 59200 29422 60000 6 spi_dat_i[17]
port 257 nsew signal input
rlabel metal2 s 30838 59200 30894 60000 6 spi_dat_i[18]
port 258 nsew signal input
rlabel metal2 s 32218 59200 32274 60000 6 spi_dat_i[19]
port 259 nsew signal input
rlabel metal2 s 5354 59200 5410 60000 6 spi_dat_i[1]
port 260 nsew signal input
rlabel metal2 s 33690 59200 33746 60000 6 spi_dat_i[20]
port 261 nsew signal input
rlabel metal2 s 35070 59200 35126 60000 6 spi_dat_i[21]
port 262 nsew signal input
rlabel metal2 s 36450 59200 36506 60000 6 spi_dat_i[22]
port 263 nsew signal input
rlabel metal2 s 37922 59200 37978 60000 6 spi_dat_i[23]
port 264 nsew signal input
rlabel metal2 s 39302 59200 39358 60000 6 spi_dat_i[24]
port 265 nsew signal input
rlabel metal2 s 40682 59200 40738 60000 6 spi_dat_i[25]
port 266 nsew signal input
rlabel metal2 s 42154 59200 42210 60000 6 spi_dat_i[26]
port 267 nsew signal input
rlabel metal2 s 43534 59200 43590 60000 6 spi_dat_i[27]
port 268 nsew signal input
rlabel metal2 s 45006 59200 45062 60000 6 spi_dat_i[28]
port 269 nsew signal input
rlabel metal2 s 46386 59200 46442 60000 6 spi_dat_i[29]
port 270 nsew signal input
rlabel metal2 s 7194 59200 7250 60000 6 spi_dat_i[2]
port 271 nsew signal input
rlabel metal2 s 47766 59200 47822 60000 6 spi_dat_i[30]
port 272 nsew signal input
rlabel metal2 s 49238 59200 49294 60000 6 spi_dat_i[31]
port 273 nsew signal input
rlabel metal2 s 9126 59200 9182 60000 6 spi_dat_i[3]
port 274 nsew signal input
rlabel metal2 s 10966 59200 11022 60000 6 spi_dat_i[4]
port 275 nsew signal input
rlabel metal2 s 12438 59200 12494 60000 6 spi_dat_i[5]
port 276 nsew signal input
rlabel metal2 s 13818 59200 13874 60000 6 spi_dat_i[6]
port 277 nsew signal input
rlabel metal2 s 15290 59200 15346 60000 6 spi_dat_i[7]
port 278 nsew signal input
rlabel metal2 s 16670 59200 16726 60000 6 spi_dat_i[8]
port 279 nsew signal input
rlabel metal2 s 18050 59200 18106 60000 6 spi_dat_i[9]
port 280 nsew signal input
rlabel metal2 s 3974 59200 4030 60000 6 spi_dat_o[0]
port 281 nsew signal output
rlabel metal2 s 19982 59200 20038 60000 6 spi_dat_o[10]
port 282 nsew signal output
rlabel metal2 s 21362 59200 21418 60000 6 spi_dat_o[11]
port 283 nsew signal output
rlabel metal2 s 22834 59200 22890 60000 6 spi_dat_o[12]
port 284 nsew signal output
rlabel metal2 s 24214 59200 24270 60000 6 spi_dat_o[13]
port 285 nsew signal output
rlabel metal2 s 25594 59200 25650 60000 6 spi_dat_o[14]
port 286 nsew signal output
rlabel metal2 s 27066 59200 27122 60000 6 spi_dat_o[15]
port 287 nsew signal output
rlabel metal2 s 28446 59200 28502 60000 6 spi_dat_o[16]
port 288 nsew signal output
rlabel metal2 s 29918 59200 29974 60000 6 spi_dat_o[17]
port 289 nsew signal output
rlabel metal2 s 31298 59200 31354 60000 6 spi_dat_o[18]
port 290 nsew signal output
rlabel metal2 s 32678 59200 32734 60000 6 spi_dat_o[19]
port 291 nsew signal output
rlabel metal2 s 5814 59200 5870 60000 6 spi_dat_o[1]
port 292 nsew signal output
rlabel metal2 s 34150 59200 34206 60000 6 spi_dat_o[20]
port 293 nsew signal output
rlabel metal2 s 35530 59200 35586 60000 6 spi_dat_o[21]
port 294 nsew signal output
rlabel metal2 s 36910 59200 36966 60000 6 spi_dat_o[22]
port 295 nsew signal output
rlabel metal2 s 38382 59200 38438 60000 6 spi_dat_o[23]
port 296 nsew signal output
rlabel metal2 s 39762 59200 39818 60000 6 spi_dat_o[24]
port 297 nsew signal output
rlabel metal2 s 41234 59200 41290 60000 6 spi_dat_o[25]
port 298 nsew signal output
rlabel metal2 s 42614 59200 42670 60000 6 spi_dat_o[26]
port 299 nsew signal output
rlabel metal2 s 43994 59200 44050 60000 6 spi_dat_o[27]
port 300 nsew signal output
rlabel metal2 s 45466 59200 45522 60000 6 spi_dat_o[28]
port 301 nsew signal output
rlabel metal2 s 46846 59200 46902 60000 6 spi_dat_o[29]
port 302 nsew signal output
rlabel metal2 s 7746 59200 7802 60000 6 spi_dat_o[2]
port 303 nsew signal output
rlabel metal2 s 48226 59200 48282 60000 6 spi_dat_o[30]
port 304 nsew signal output
rlabel metal2 s 49698 59200 49754 60000 6 spi_dat_o[31]
port 305 nsew signal output
rlabel metal2 s 9586 59200 9642 60000 6 spi_dat_o[3]
port 306 nsew signal output
rlabel metal2 s 11518 59200 11574 60000 6 spi_dat_o[4]
port 307 nsew signal output
rlabel metal2 s 12898 59200 12954 60000 6 spi_dat_o[5]
port 308 nsew signal output
rlabel metal2 s 14278 59200 14334 60000 6 spi_dat_o[6]
port 309 nsew signal output
rlabel metal2 s 15750 59200 15806 60000 6 spi_dat_o[7]
port 310 nsew signal output
rlabel metal2 s 17130 59200 17186 60000 6 spi_dat_o[8]
port 311 nsew signal output
rlabel metal2 s 18510 59200 18566 60000 6 spi_dat_o[9]
port 312 nsew signal output
rlabel metal2 s 1122 59200 1178 60000 6 spi_err_i
port 313 nsew signal input
rlabel metal2 s 1582 59200 1638 60000 6 spi_rty_i
port 314 nsew signal input
rlabel metal2 s 4434 59200 4490 60000 6 spi_sel_o[0]
port 315 nsew signal output
rlabel metal2 s 6274 59200 6330 60000 6 spi_sel_o[1]
port 316 nsew signal output
rlabel metal2 s 8206 59200 8262 60000 6 spi_sel_o[2]
port 317 nsew signal output
rlabel metal2 s 10046 59200 10102 60000 6 spi_sel_o[3]
port 318 nsew signal output
rlabel metal2 s 2042 59200 2098 60000 6 spi_stb_o
port 319 nsew signal output
rlabel metal2 s 2502 59200 2558 60000 6 spi_we_o
port 320 nsew signal output
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 321 nsew power input
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 321 nsew power input
rlabel metal4 s 65648 2128 65968 57712 6 vccd1
port 321 nsew power input
rlabel metal4 s 96368 2128 96688 57712 6 vccd1
port 321 nsew power input
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 322 nsew ground input
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 322 nsew ground input
rlabel metal4 s 81008 2128 81328 57712 6 vssd1
port 322 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 100000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 13328732
string GDS_FILE /home/q3k/sky130/qf105/openlane/mkQF100Fabric/runs/mkQF100Fabric/results/finishing/mkQF100Fabric.magic.gds
string GDS_START 831944
<< end >>

