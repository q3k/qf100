magic
tech sky130A
magscale 1 2
timestamp 1647787412
<< viali >>
rect 12265 47209 12299 47243
rect 20269 47209 20303 47243
rect 28273 47209 28307 47243
rect 4261 47005 4295 47039
rect 12081 47005 12115 47039
rect 20085 47005 20119 47039
rect 28089 47005 28123 47039
rect 36185 47005 36219 47039
rect 4629 46937 4663 46971
rect 36277 46869 36311 46903
rect 12449 46665 12483 46699
rect 12633 46529 12667 46563
rect 16129 46529 16163 46563
rect 15945 46325 15979 46359
rect 22017 34561 22051 34595
rect 21833 34357 21867 34391
rect 19441 33949 19475 33983
rect 20545 33949 20579 33983
rect 22477 33949 22511 33983
rect 22661 33949 22695 33983
rect 22845 33949 22879 33983
rect 23489 33949 23523 33983
rect 20790 33881 20824 33915
rect 19257 33813 19291 33847
rect 21925 33813 21959 33847
rect 23305 33813 23339 33847
rect 17693 33609 17727 33643
rect 20269 33609 20303 33643
rect 21281 33609 21315 33643
rect 18582 33541 18616 33575
rect 22652 33541 22686 33575
rect 17877 33473 17911 33507
rect 20453 33473 20487 33507
rect 20913 33473 20947 33507
rect 21097 33473 21131 33507
rect 24409 33473 24443 33507
rect 18337 33405 18371 33439
rect 22385 33405 22419 33439
rect 19717 33269 19751 33303
rect 23765 33269 23799 33303
rect 24225 33269 24259 33303
rect 17877 33065 17911 33099
rect 18705 33065 18739 33099
rect 23305 33065 23339 33099
rect 24777 33065 24811 33099
rect 17509 32929 17543 32963
rect 18337 32929 18371 32963
rect 22937 32929 22971 32963
rect 24409 32929 24443 32963
rect 17049 32861 17083 32895
rect 17693 32861 17727 32895
rect 18521 32861 18555 32895
rect 19257 32861 19291 32895
rect 19524 32861 19558 32895
rect 21097 32861 21131 32895
rect 21364 32861 21398 32895
rect 23121 32861 23155 32895
rect 24593 32861 24627 32895
rect 16865 32725 16899 32759
rect 20637 32725 20671 32759
rect 22477 32725 22511 32759
rect 19717 32521 19751 32555
rect 21281 32521 21315 32555
rect 22661 32521 22695 32555
rect 17202 32453 17236 32487
rect 20913 32453 20947 32487
rect 22385 32453 22419 32487
rect 23664 32453 23698 32487
rect 16957 32385 16991 32419
rect 19165 32385 19199 32419
rect 19349 32385 19383 32419
rect 19441 32385 19475 32419
rect 19533 32385 19567 32419
rect 20729 32385 20763 32419
rect 21005 32385 21039 32419
rect 21097 32385 21131 32419
rect 22109 32385 22143 32419
rect 22293 32385 22327 32419
rect 22477 32385 22511 32419
rect 23397 32385 23431 32419
rect 25421 32385 25455 32419
rect 18337 32181 18371 32215
rect 24777 32181 24811 32215
rect 25237 32181 25271 32215
rect 17693 31977 17727 32011
rect 19809 31977 19843 32011
rect 21465 31977 21499 32011
rect 21925 31977 21959 32011
rect 23673 31977 23707 32011
rect 18705 31909 18739 31943
rect 22477 31841 22511 31875
rect 24409 31841 24443 31875
rect 17417 31773 17451 31807
rect 17509 31773 17543 31807
rect 18153 31773 18187 31807
rect 18521 31773 18555 31807
rect 19257 31773 19291 31807
rect 19441 31773 19475 31807
rect 19625 31773 19659 31807
rect 20913 31773 20947 31807
rect 21189 31773 21223 31807
rect 21281 31773 21315 31807
rect 23121 31773 23155 31807
rect 23305 31773 23339 31807
rect 23489 31773 23523 31807
rect 24676 31773 24710 31807
rect 18337 31705 18371 31739
rect 18429 31705 18463 31739
rect 19533 31705 19567 31739
rect 21097 31705 21131 31739
rect 23397 31705 23431 31739
rect 22293 31637 22327 31671
rect 22385 31637 22419 31671
rect 25789 31637 25823 31671
rect 18981 31433 19015 31467
rect 20269 31433 20303 31467
rect 21833 31433 21867 31467
rect 23029 31433 23063 31467
rect 25605 31433 25639 31467
rect 18245 31365 18279 31399
rect 20729 31365 20763 31399
rect 23397 31365 23431 31399
rect 24409 31365 24443 31399
rect 24501 31365 24535 31399
rect 16865 31297 16899 31331
rect 17969 31297 18003 31331
rect 18153 31297 18187 31331
rect 18337 31297 18371 31331
rect 19349 31297 19383 31331
rect 19441 31297 19475 31331
rect 20637 31297 20671 31331
rect 22201 31297 22235 31331
rect 22293 31297 22327 31331
rect 24225 31297 24259 31331
rect 24593 31297 24627 31331
rect 25421 31297 25455 31331
rect 26249 31297 26283 31331
rect 19625 31229 19659 31263
rect 20913 31229 20947 31263
rect 22385 31229 22419 31263
rect 23489 31229 23523 31263
rect 23581 31229 23615 31263
rect 25237 31229 25271 31263
rect 24777 31161 24811 31195
rect 16681 31093 16715 31127
rect 18521 31093 18555 31127
rect 26065 31093 26099 31127
rect 24409 30889 24443 30923
rect 18705 30821 18739 30855
rect 16773 30753 16807 30787
rect 21281 30753 21315 30787
rect 21557 30753 21591 30787
rect 23305 30753 23339 30787
rect 25053 30753 25087 30787
rect 16957 30685 16991 30719
rect 18153 30685 18187 30719
rect 18429 30685 18463 30719
rect 18521 30685 18555 30719
rect 19257 30685 19291 30719
rect 19533 30685 19567 30719
rect 23029 30685 23063 30719
rect 24593 30685 24627 30719
rect 18337 30617 18371 30651
rect 25320 30617 25354 30651
rect 17141 30549 17175 30583
rect 26433 30549 26467 30583
rect 20269 30345 20303 30379
rect 23305 30345 23339 30379
rect 24041 30345 24075 30379
rect 26341 30345 26375 30379
rect 16129 30277 16163 30311
rect 20177 30277 20211 30311
rect 25237 30277 25271 30311
rect 15945 30209 15979 30243
rect 16937 30209 16971 30243
rect 18797 30209 18831 30243
rect 21833 30209 21867 30243
rect 22017 30209 22051 30243
rect 23213 30209 23247 30243
rect 24225 30209 24259 30243
rect 24961 30209 24995 30243
rect 25145 30209 25179 30243
rect 25329 30209 25363 30243
rect 26157 30209 26191 30243
rect 27169 30209 27203 30243
rect 15761 30141 15795 30175
rect 16681 30141 16715 30175
rect 18521 30141 18555 30175
rect 20453 30141 20487 30175
rect 21925 30141 21959 30175
rect 23397 30141 23431 30175
rect 25973 30141 26007 30175
rect 26985 30141 27019 30175
rect 19809 30073 19843 30107
rect 22845 30073 22879 30107
rect 25513 30073 25547 30107
rect 18061 30005 18095 30039
rect 27353 30005 27387 30039
rect 14749 29801 14783 29835
rect 19257 29801 19291 29835
rect 20545 29801 20579 29835
rect 21925 29801 21959 29835
rect 22109 29801 22143 29835
rect 22753 29801 22787 29835
rect 23397 29801 23431 29835
rect 24685 29801 24719 29835
rect 15393 29733 15427 29767
rect 16405 29665 16439 29699
rect 19901 29665 19935 29699
rect 21097 29665 21131 29699
rect 25237 29665 25271 29699
rect 26433 29665 26467 29699
rect 14933 29597 14967 29631
rect 15669 29597 15703 29631
rect 16672 29597 16706 29631
rect 19625 29597 19659 29631
rect 20913 29597 20947 29631
rect 23397 29597 23431 29631
rect 23581 29597 23615 29631
rect 28457 29597 28491 29631
rect 15393 29529 15427 29563
rect 21741 29529 21775 29563
rect 22569 29529 22603 29563
rect 25053 29529 25087 29563
rect 26700 29529 26734 29563
rect 15577 29461 15611 29495
rect 17785 29461 17819 29495
rect 19717 29461 19751 29495
rect 21005 29461 21039 29495
rect 21941 29461 21975 29495
rect 22769 29461 22803 29495
rect 22937 29461 22971 29495
rect 25145 29461 25179 29495
rect 27813 29461 27847 29495
rect 28273 29461 28307 29495
rect 16773 29257 16807 29291
rect 18613 29257 18647 29291
rect 19073 29257 19107 29291
rect 19901 29257 19935 29291
rect 21189 29257 21223 29291
rect 22861 29257 22895 29291
rect 23029 29257 23063 29291
rect 23673 29257 23707 29291
rect 25605 29257 25639 29291
rect 27537 29257 27571 29291
rect 21833 29189 21867 29223
rect 22049 29189 22083 29223
rect 22661 29189 22695 29223
rect 27169 29189 27203 29223
rect 13093 29121 13127 29155
rect 13277 29121 13311 29155
rect 14197 29121 14231 29155
rect 14464 29121 14498 29155
rect 16957 29121 16991 29155
rect 18981 29121 19015 29155
rect 20085 29121 20119 29155
rect 21097 29121 21131 29155
rect 21281 29121 21315 29155
rect 23857 29121 23891 29155
rect 25973 29121 26007 29155
rect 26985 29121 27019 29155
rect 27261 29121 27295 29155
rect 27353 29121 27387 29155
rect 19257 29053 19291 29087
rect 24317 29053 24351 29087
rect 24593 29053 24627 29087
rect 26065 29053 26099 29087
rect 26249 29053 26283 29087
rect 15577 28985 15611 29019
rect 22201 28985 22235 29019
rect 13093 28917 13127 28951
rect 22017 28917 22051 28951
rect 22845 28917 22879 28951
rect 16681 28713 16715 28747
rect 21005 28713 21039 28747
rect 22109 28713 22143 28747
rect 23581 28713 23615 28747
rect 28549 28713 28583 28747
rect 12173 28577 12207 28611
rect 16773 28577 16807 28611
rect 24685 28577 24719 28611
rect 26525 28577 26559 28611
rect 8953 28509 8987 28543
rect 11069 28509 11103 28543
rect 11158 28509 11192 28543
rect 11253 28509 11287 28543
rect 11437 28509 11471 28543
rect 12440 28509 12474 28543
rect 14657 28509 14691 28543
rect 16497 28509 16531 28543
rect 16589 28509 16623 28543
rect 19625 28509 19659 28543
rect 19809 28509 19843 28543
rect 20729 28509 20763 28543
rect 20821 28509 20855 28543
rect 21833 28509 21867 28543
rect 22937 28509 22971 28543
rect 23581 28509 23615 28543
rect 23765 28509 23799 28543
rect 24961 28509 24995 28543
rect 27169 28509 27203 28543
rect 9198 28441 9232 28475
rect 14924 28441 14958 28475
rect 20453 28441 20487 28475
rect 21557 28441 21591 28475
rect 22569 28441 22603 28475
rect 23121 28441 23155 28475
rect 27436 28441 27470 28475
rect 10333 28373 10367 28407
rect 10793 28373 10827 28407
rect 13553 28373 13587 28407
rect 16037 28373 16071 28407
rect 19717 28373 19751 28407
rect 20637 28373 20671 28407
rect 21741 28373 21775 28407
rect 21925 28373 21959 28407
rect 22753 28373 22787 28407
rect 22845 28373 22879 28407
rect 25973 28373 26007 28407
rect 26341 28373 26375 28407
rect 26433 28373 26467 28407
rect 13093 28169 13127 28203
rect 15117 28169 15151 28203
rect 17325 28169 17359 28203
rect 20637 28169 20671 28203
rect 27813 28169 27847 28203
rect 9496 28101 9530 28135
rect 13553 28101 13587 28135
rect 26065 28101 26099 28135
rect 8585 28033 8619 28067
rect 8769 28033 8803 28067
rect 11980 28033 12014 28067
rect 13737 28033 13771 28067
rect 14473 28033 14507 28067
rect 14657 28033 14691 28067
rect 15301 28033 15335 28067
rect 15393 28033 15427 28067
rect 15577 28033 15611 28067
rect 15669 28033 15703 28067
rect 16681 28033 16715 28067
rect 16865 28033 16899 28067
rect 17509 28033 17543 28067
rect 18613 28033 18647 28067
rect 18797 28033 18831 28067
rect 19349 28033 19383 28067
rect 20177 28033 20211 28067
rect 20453 28033 20487 28067
rect 21281 28033 21315 28067
rect 22109 28033 22143 28067
rect 23765 28033 23799 28067
rect 23857 28033 23891 28067
rect 24593 28033 24627 28067
rect 25881 28033 25915 28067
rect 26157 28033 26191 28067
rect 26249 28033 26283 28067
rect 26985 28033 27019 28067
rect 27169 28033 27203 28067
rect 27353 28033 27387 28067
rect 27997 28033 28031 28067
rect 9229 27965 9263 27999
rect 11713 27965 11747 27999
rect 14565 27965 14599 27999
rect 17785 27965 17819 27999
rect 19533 27965 19567 27999
rect 20269 27965 20303 27999
rect 21833 27965 21867 27999
rect 23949 27965 23983 27999
rect 24869 27965 24903 27999
rect 18613 27897 18647 27931
rect 26433 27897 26467 27931
rect 8585 27829 8619 27863
rect 10609 27829 10643 27863
rect 13921 27829 13955 27863
rect 16773 27829 16807 27863
rect 17693 27829 17727 27863
rect 20177 27829 20211 27863
rect 21097 27829 21131 27863
rect 23397 27829 23431 27863
rect 8401 27625 8435 27659
rect 15853 27625 15887 27659
rect 20545 27625 20579 27659
rect 22937 27625 22971 27659
rect 23305 27625 23339 27659
rect 9689 27557 9723 27591
rect 14197 27557 14231 27591
rect 21005 27557 21039 27591
rect 21925 27557 21959 27591
rect 22477 27557 22511 27591
rect 8217 27489 8251 27523
rect 9321 27489 9355 27523
rect 12725 27489 12759 27523
rect 14381 27489 14415 27523
rect 15761 27489 15795 27523
rect 18705 27489 18739 27523
rect 19533 27489 19567 27523
rect 19809 27489 19843 27523
rect 23029 27489 23063 27523
rect 26709 27489 26743 27523
rect 8033 27421 8067 27455
rect 8401 27421 8435 27455
rect 8953 27421 8987 27455
rect 9137 27421 9171 27455
rect 9229 27421 9263 27455
rect 9505 27421 9539 27455
rect 10701 27421 10735 27455
rect 10957 27421 10991 27455
rect 13001 27421 13035 27455
rect 14105 27421 14139 27455
rect 14841 27421 14875 27455
rect 15485 27421 15519 27455
rect 16497 27421 16531 27455
rect 18337 27421 18371 27455
rect 18521 27421 18555 27455
rect 19441 27421 19475 27455
rect 20729 27421 20763 27455
rect 20821 27421 20855 27455
rect 22201 27421 22235 27455
rect 22293 27421 22327 27455
rect 22937 27421 22971 27455
rect 24409 27421 24443 27455
rect 24593 27421 24627 27455
rect 24777 27421 24811 27455
rect 25697 27421 25731 27455
rect 25973 27421 26007 27455
rect 26065 27421 26099 27455
rect 26893 27421 26927 27455
rect 27721 27421 27755 27455
rect 16742 27353 16776 27387
rect 20545 27353 20579 27387
rect 22109 27353 22143 27387
rect 24685 27353 24719 27387
rect 25881 27353 25915 27387
rect 8125 27285 8159 27319
rect 12081 27285 12115 27319
rect 14381 27285 14415 27319
rect 14933 27285 14967 27319
rect 16037 27285 16071 27319
rect 17877 27285 17911 27319
rect 24961 27285 24995 27319
rect 26249 27285 26283 27319
rect 27077 27285 27111 27319
rect 27537 27285 27571 27319
rect 8033 27081 8067 27115
rect 9137 27081 9171 27115
rect 9873 27081 9907 27115
rect 10977 27081 11011 27115
rect 13461 27081 13495 27115
rect 13645 27081 13679 27115
rect 14657 27081 14691 27115
rect 16037 27081 16071 27115
rect 17509 27081 17543 27115
rect 20085 27081 20119 27115
rect 20545 27081 20579 27115
rect 25513 27081 25547 27115
rect 25881 27081 25915 27115
rect 25973 27081 26007 27115
rect 28365 27081 28399 27115
rect 16865 27013 16899 27047
rect 19901 27013 19935 27047
rect 22845 27013 22879 27047
rect 27261 27013 27295 27047
rect 7757 26945 7791 26979
rect 8861 26945 8895 26979
rect 9597 26945 9631 26979
rect 11529 26945 11563 26979
rect 12449 26945 12483 26979
rect 13586 26945 13620 26979
rect 14105 26945 14139 26979
rect 14841 26945 14875 26979
rect 14933 26945 14967 26979
rect 15117 26945 15151 26979
rect 15301 26945 15335 26979
rect 15945 26945 15979 26979
rect 16129 26945 16163 26979
rect 17877 26945 17911 26979
rect 18889 26945 18923 26979
rect 19717 26945 19751 26979
rect 20729 26945 20763 26979
rect 21925 26945 21959 26979
rect 23673 26945 23707 26979
rect 23940 26945 23974 26979
rect 26985 26945 27019 26979
rect 27169 26945 27203 26979
rect 27353 26945 27387 26979
rect 28181 26945 28215 26979
rect 8033 26877 8067 26911
rect 8493 26877 8527 26911
rect 8953 26877 8987 26911
rect 9873 26877 9907 26911
rect 10333 26877 10367 26911
rect 10701 26877 10735 26911
rect 10793 26877 10827 26911
rect 12173 26877 12207 26911
rect 15025 26877 15059 26911
rect 17969 26877 18003 26911
rect 18153 26877 18187 26911
rect 18797 26877 18831 26911
rect 22017 26877 22051 26911
rect 26065 26877 26099 26911
rect 27997 26877 28031 26911
rect 9689 26809 9723 26843
rect 14013 26809 14047 26843
rect 17049 26809 17083 26843
rect 19257 26809 19291 26843
rect 27537 26809 27571 26843
rect 7849 26741 7883 26775
rect 11621 26741 11655 26775
rect 22109 26741 22143 26775
rect 22293 26741 22327 26775
rect 22937 26741 22971 26775
rect 25053 26741 25087 26775
rect 8033 26537 8067 26571
rect 8401 26537 8435 26571
rect 8953 26537 8987 26571
rect 9413 26537 9447 26571
rect 11161 26537 11195 26571
rect 12081 26537 12115 26571
rect 14841 26537 14875 26571
rect 17049 26537 17083 26571
rect 18153 26537 18187 26571
rect 19349 26537 19383 26571
rect 20177 26537 20211 26571
rect 20821 26537 20855 26571
rect 21189 26537 21223 26571
rect 22661 26537 22695 26571
rect 25513 26537 25547 26571
rect 9965 26469 9999 26503
rect 14381 26469 14415 26503
rect 23305 26469 23339 26503
rect 28273 26469 28307 26503
rect 10425 26401 10459 26435
rect 10609 26401 10643 26435
rect 13461 26401 13495 26435
rect 15485 26401 15519 26435
rect 17509 26401 17543 26435
rect 22201 26401 22235 26435
rect 26065 26401 26099 26435
rect 26893 26401 26927 26435
rect 8033 26333 8067 26367
rect 8217 26333 8251 26367
rect 8953 26333 8987 26367
rect 9137 26333 9171 26367
rect 9229 26333 9263 26367
rect 10333 26333 10367 26367
rect 11345 26333 11379 26367
rect 11529 26333 11563 26367
rect 11621 26333 11655 26367
rect 12265 26333 12299 26367
rect 12541 26333 12575 26367
rect 12725 26333 12759 26367
rect 13277 26333 13311 26367
rect 15025 26333 15059 26367
rect 15117 26333 15151 26367
rect 15393 26333 15427 26367
rect 16221 26333 16255 26367
rect 16313 26333 16347 26367
rect 16405 26333 16439 26367
rect 16589 26333 16623 26367
rect 17233 26333 17267 26367
rect 17417 26333 17451 26367
rect 19257 26333 19291 26367
rect 19441 26333 19475 26367
rect 20361 26333 20395 26367
rect 20821 26333 20855 26367
rect 20913 26333 20947 26367
rect 21925 26333 21959 26367
rect 22109 26333 22143 26367
rect 22661 26333 22695 26367
rect 22845 26333 22879 26367
rect 23489 26333 23523 26367
rect 24409 26333 24443 26367
rect 24593 26333 24627 26367
rect 25973 26333 26007 26367
rect 14197 26265 14231 26299
rect 17969 26265 18003 26299
rect 24777 26265 24811 26299
rect 27138 26265 27172 26299
rect 15945 26197 15979 26231
rect 18169 26197 18203 26231
rect 18337 26197 18371 26231
rect 25881 26197 25915 26231
rect 9229 25993 9263 26027
rect 12173 25993 12207 26027
rect 12725 25993 12759 26027
rect 16037 25993 16071 26027
rect 17969 25993 18003 26027
rect 19993 25993 20027 26027
rect 23581 25993 23615 26027
rect 25513 25993 25547 26027
rect 9597 25925 9631 25959
rect 10977 25925 11011 25959
rect 14372 25925 14406 25959
rect 25421 25925 25455 25959
rect 27436 25925 27470 25959
rect 7113 25857 7147 25891
rect 7297 25857 7331 25891
rect 7757 25857 7791 25891
rect 7941 25857 7975 25891
rect 8125 25857 8159 25891
rect 8309 25857 8343 25891
rect 10793 25857 10827 25891
rect 12081 25857 12115 25891
rect 12909 25857 12943 25891
rect 14105 25857 14139 25891
rect 15945 25857 15979 25891
rect 17049 25857 17083 25891
rect 17877 25857 17911 25891
rect 18061 25857 18095 25891
rect 18889 25857 18923 25891
rect 19809 25857 19843 25891
rect 19993 25857 20027 25891
rect 20453 25857 20487 25891
rect 22017 25857 22051 25891
rect 22109 25857 22143 25891
rect 22293 25857 22327 25891
rect 22385 25857 22419 25891
rect 22845 25857 22879 25891
rect 23029 25857 23063 25891
rect 23489 25857 23523 25891
rect 23685 25857 23719 25891
rect 24317 25857 24351 25891
rect 26249 25857 26283 25891
rect 27169 25857 27203 25891
rect 7205 25789 7239 25823
rect 8033 25789 8067 25823
rect 9689 25789 9723 25823
rect 9873 25789 9907 25823
rect 13001 25789 13035 25823
rect 13093 25789 13127 25823
rect 13185 25789 13219 25823
rect 16957 25789 16991 25823
rect 18797 25789 18831 25823
rect 20729 25789 20763 25823
rect 22937 25789 22971 25823
rect 15485 25721 15519 25755
rect 17417 25721 17451 25755
rect 26065 25721 26099 25755
rect 8493 25653 8527 25687
rect 19165 25653 19199 25687
rect 21833 25653 21867 25687
rect 24133 25653 24167 25687
rect 28549 25653 28583 25687
rect 9597 25449 9631 25483
rect 10149 25449 10183 25483
rect 10701 25449 10735 25483
rect 11897 25449 11931 25483
rect 12541 25449 12575 25483
rect 14381 25449 14415 25483
rect 15117 25449 15151 25483
rect 17417 25449 17451 25483
rect 17601 25449 17635 25483
rect 19441 25449 19475 25483
rect 20453 25449 20487 25483
rect 21189 25449 21223 25483
rect 22477 25449 22511 25483
rect 26893 25449 26927 25483
rect 8401 25381 8435 25415
rect 11161 25381 11195 25415
rect 20637 25381 20671 25415
rect 26157 25381 26191 25415
rect 9413 25313 9447 25347
rect 10793 25313 10827 25347
rect 24777 25313 24811 25347
rect 7021 25245 7055 25279
rect 7288 25245 7322 25279
rect 9321 25245 9355 25279
rect 10057 25245 10091 25279
rect 10977 25245 11011 25279
rect 11713 25245 11747 25279
rect 11805 25245 11839 25279
rect 12725 25245 12759 25279
rect 13001 25245 13035 25279
rect 14381 25245 14415 25279
rect 14657 25245 14691 25279
rect 15301 25245 15335 25279
rect 15393 25245 15427 25279
rect 16681 25245 16715 25279
rect 21373 25245 21407 25279
rect 21465 25245 21499 25279
rect 21649 25245 21683 25279
rect 21741 25245 21775 25279
rect 22753 25245 22787 25279
rect 22845 25245 22879 25279
rect 22937 25245 22971 25279
rect 23121 25245 23155 25279
rect 23857 25245 23891 25279
rect 24409 25245 24443 25279
rect 24593 25245 24627 25279
rect 25789 25245 25823 25279
rect 27077 25245 27111 25279
rect 10701 25177 10735 25211
rect 15669 25177 15703 25211
rect 15761 25177 15795 25211
rect 17233 25177 17267 25211
rect 19257 25177 19291 25211
rect 19473 25177 19507 25211
rect 20085 25177 20119 25211
rect 20462 25177 20496 25211
rect 25973 25177 26007 25211
rect 8953 25109 8987 25143
rect 12081 25109 12115 25143
rect 12909 25109 12943 25143
rect 14565 25109 14599 25143
rect 16681 25109 16715 25143
rect 17443 25109 17477 25143
rect 19625 25109 19659 25143
rect 23673 25109 23707 25143
rect 8125 24905 8159 24939
rect 8769 24905 8803 24939
rect 9137 24905 9171 24939
rect 25513 24905 25547 24939
rect 10333 24837 10367 24871
rect 10425 24837 10459 24871
rect 23918 24837 23952 24871
rect 25881 24837 25915 24871
rect 8033 24769 8067 24803
rect 8217 24769 8251 24803
rect 10149 24769 10183 24803
rect 10517 24769 10551 24803
rect 11529 24769 11563 24803
rect 11713 24769 11747 24803
rect 13093 24769 13127 24803
rect 13369 24769 13403 24803
rect 13553 24769 13587 24803
rect 14197 24769 14231 24803
rect 15577 24769 15611 24803
rect 15669 24769 15703 24803
rect 16681 24769 16715 24803
rect 16957 24769 16991 24803
rect 17049 24769 17083 24803
rect 18061 24769 18095 24803
rect 18797 24769 18831 24803
rect 18981 24769 19015 24803
rect 20913 24769 20947 24803
rect 21189 24769 21223 24803
rect 22477 24769 22511 24803
rect 22569 24769 22603 24803
rect 22661 24769 22695 24803
rect 22845 24769 22879 24803
rect 27804 24769 27838 24803
rect 9229 24701 9263 24735
rect 9413 24701 9447 24735
rect 14013 24701 14047 24735
rect 15301 24701 15335 24735
rect 15485 24701 15519 24735
rect 15761 24701 15795 24735
rect 19809 24701 19843 24735
rect 21281 24701 21315 24735
rect 22201 24701 22235 24735
rect 23673 24701 23707 24735
rect 25973 24701 26007 24735
rect 26157 24701 26191 24735
rect 27537 24701 27571 24735
rect 14381 24633 14415 24667
rect 18245 24633 18279 24667
rect 10701 24565 10735 24599
rect 11897 24565 11931 24599
rect 12909 24565 12943 24599
rect 25053 24565 25087 24599
rect 28917 24565 28951 24599
rect 9597 24361 9631 24395
rect 10793 24361 10827 24395
rect 12909 24361 12943 24395
rect 14289 24361 14323 24395
rect 15301 24361 15335 24395
rect 16957 24361 16991 24395
rect 19717 24361 19751 24395
rect 19901 24361 19935 24395
rect 21465 24361 21499 24395
rect 22109 24361 22143 24395
rect 23121 24361 23155 24395
rect 26065 24361 26099 24395
rect 26525 24361 26559 24395
rect 28457 24361 28491 24395
rect 15117 24293 15151 24327
rect 21649 24293 21683 24327
rect 11529 24225 11563 24259
rect 11621 24225 11655 24259
rect 13093 24225 13127 24259
rect 17509 24225 17543 24259
rect 17785 24225 17819 24259
rect 23581 24225 23615 24259
rect 23765 24225 23799 24259
rect 24685 24225 24719 24259
rect 26985 24225 27019 24259
rect 27169 24225 27203 24259
rect 27997 24225 28031 24259
rect 9505 24157 9539 24191
rect 10517 24157 10551 24191
rect 10609 24157 10643 24191
rect 10885 24157 10919 24191
rect 11713 24157 11747 24191
rect 12265 24157 12299 24191
rect 12909 24157 12943 24191
rect 13185 24157 13219 24191
rect 15761 24157 15795 24191
rect 15945 24157 15979 24191
rect 16129 24157 16163 24191
rect 16773 24157 16807 24191
rect 20361 24157 20395 24191
rect 22293 24157 22327 24191
rect 22385 24157 22419 24191
rect 22569 24157 22603 24191
rect 22661 24157 22695 24191
rect 28641 24157 28675 24191
rect 10333 24089 10367 24123
rect 14197 24089 14231 24123
rect 14841 24089 14875 24123
rect 16037 24089 16071 24123
rect 19533 24089 19567 24123
rect 19749 24089 19783 24123
rect 21281 24089 21315 24123
rect 24952 24089 24986 24123
rect 27813 24089 27847 24123
rect 11345 24021 11379 24055
rect 12357 24021 12391 24055
rect 13369 24021 13403 24055
rect 16313 24021 16347 24055
rect 20545 24021 20579 24055
rect 21481 24021 21515 24055
rect 23489 24021 23523 24055
rect 26893 24021 26927 24055
rect 14841 23817 14875 23851
rect 17049 23817 17083 23851
rect 19625 23817 19659 23851
rect 21189 23817 21223 23851
rect 21833 23817 21867 23851
rect 23949 23817 23983 23851
rect 25697 23817 25731 23851
rect 26985 23817 27019 23851
rect 28549 23817 28583 23851
rect 11621 23749 11655 23783
rect 13461 23749 13495 23783
rect 15945 23749 15979 23783
rect 18490 23749 18524 23783
rect 23673 23749 23707 23783
rect 26157 23749 26191 23783
rect 27445 23749 27479 23783
rect 7297 23681 7331 23715
rect 7564 23681 7598 23715
rect 9965 23681 9999 23715
rect 10609 23681 10643 23715
rect 10701 23681 10735 23715
rect 10885 23681 10919 23715
rect 10977 23681 11011 23715
rect 11529 23681 11563 23715
rect 11713 23681 11747 23715
rect 12449 23681 12483 23715
rect 12541 23681 12575 23715
rect 12633 23681 12667 23715
rect 12793 23681 12827 23715
rect 13277 23681 13311 23715
rect 13553 23681 13587 23715
rect 13650 23703 13684 23737
rect 14197 23681 14231 23715
rect 14381 23681 14415 23715
rect 15301 23681 15335 23715
rect 18245 23681 18279 23715
rect 21097 23681 21131 23715
rect 22201 23681 22235 23715
rect 23397 23681 23431 23715
rect 23581 23681 23615 23715
rect 23765 23681 23799 23715
rect 24593 23681 24627 23715
rect 26065 23681 26099 23715
rect 27353 23681 27387 23715
rect 28365 23681 28399 23715
rect 29193 23681 29227 23715
rect 29837 23681 29871 23715
rect 9781 23613 9815 23647
rect 13369 23613 13403 23647
rect 15025 23613 15059 23647
rect 15117 23613 15151 23647
rect 15209 23613 15243 23647
rect 16865 23613 16899 23647
rect 17233 23613 17267 23647
rect 22293 23613 22327 23647
rect 22385 23613 22419 23647
rect 24409 23613 24443 23647
rect 26341 23613 26375 23647
rect 27537 23613 27571 23647
rect 28181 23613 28215 23647
rect 9597 23545 9631 23579
rect 16129 23545 16163 23579
rect 8677 23477 8711 23511
rect 9781 23477 9815 23511
rect 9873 23477 9907 23511
rect 10425 23477 10459 23511
rect 12173 23477 12207 23511
rect 14197 23477 14231 23511
rect 17233 23477 17267 23511
rect 24777 23477 24811 23511
rect 29009 23477 29043 23511
rect 29653 23477 29687 23511
rect 8309 23273 8343 23307
rect 8953 23273 8987 23307
rect 11345 23273 11379 23307
rect 13001 23273 13035 23307
rect 14105 23273 14139 23307
rect 14749 23273 14783 23307
rect 17509 23273 17543 23307
rect 18245 23273 18279 23307
rect 22477 23273 22511 23307
rect 24961 23273 24995 23307
rect 27353 23273 27387 23307
rect 28641 23273 28675 23307
rect 10057 23205 10091 23239
rect 13185 23205 13219 23239
rect 23673 23205 23707 23239
rect 12541 23137 12575 23171
rect 14933 23137 14967 23171
rect 15025 23137 15059 23171
rect 16129 23137 16163 23171
rect 23121 23137 23155 23171
rect 29561 23137 29595 23171
rect 9229 23069 9263 23103
rect 9321 23069 9355 23103
rect 9413 23069 9447 23103
rect 9597 23069 9631 23103
rect 10057 23069 10091 23103
rect 10241 23069 10275 23103
rect 10333 23069 10367 23103
rect 11621 23069 11655 23103
rect 11713 23069 11747 23103
rect 11805 23069 11839 23103
rect 11989 23069 12023 23103
rect 12633 23069 12667 23103
rect 13001 23069 13035 23103
rect 14105 23069 14139 23103
rect 14289 23069 14323 23103
rect 15393 23069 15427 23103
rect 16396 23069 16430 23103
rect 17969 23069 18003 23103
rect 18061 23069 18095 23103
rect 18337 23069 18371 23103
rect 20637 23069 20671 23103
rect 23857 23069 23891 23103
rect 24409 23069 24443 23103
rect 24777 23069 24811 23103
rect 25605 23069 25639 23103
rect 26157 23069 26191 23103
rect 26801 23069 26835 23103
rect 27169 23069 27203 23103
rect 28273 23069 28307 23103
rect 28457 23069 28491 23103
rect 29817 23069 29851 23103
rect 8217 23001 8251 23035
rect 20882 23001 20916 23035
rect 24593 23001 24627 23035
rect 24685 23001 24719 23035
rect 26985 23001 27019 23035
rect 27077 23001 27111 23035
rect 15117 22933 15151 22967
rect 15301 22933 15335 22967
rect 18153 22933 18187 22967
rect 22017 22933 22051 22967
rect 22845 22933 22879 22967
rect 22937 22933 22971 22967
rect 25421 22933 25455 22967
rect 26249 22933 26283 22967
rect 30941 22933 30975 22967
rect 7113 22729 7147 22763
rect 10241 22729 10275 22763
rect 10885 22729 10919 22763
rect 11713 22729 11747 22763
rect 12265 22729 12299 22763
rect 12725 22729 12759 22763
rect 13737 22729 13771 22763
rect 13921 22729 13955 22763
rect 14381 22729 14415 22763
rect 15577 22729 15611 22763
rect 16957 22729 16991 22763
rect 21833 22729 21867 22763
rect 25881 22729 25915 22763
rect 28089 22729 28123 22763
rect 9321 22661 9355 22695
rect 10793 22661 10827 22695
rect 13645 22661 13679 22695
rect 23581 22661 23615 22695
rect 24768 22661 24802 22695
rect 27813 22661 27847 22695
rect 28816 22661 28850 22695
rect 6929 22593 6963 22627
rect 7113 22593 7147 22627
rect 7573 22593 7607 22627
rect 8217 22593 8251 22627
rect 8401 22593 8435 22627
rect 9137 22593 9171 22627
rect 9413 22593 9447 22627
rect 9873 22593 9907 22627
rect 11621 22593 11655 22627
rect 12541 22593 12575 22627
rect 12633 22593 12667 22627
rect 13553 22593 13587 22627
rect 14657 22593 14691 22627
rect 14841 22593 14875 22627
rect 15485 22593 15519 22627
rect 16773 22593 16807 22627
rect 16957 22593 16991 22627
rect 17601 22593 17635 22627
rect 18521 22593 18555 22627
rect 19349 22593 19383 22627
rect 22201 22593 22235 22627
rect 22293 22593 22327 22627
rect 23397 22593 23431 22627
rect 23673 22593 23707 22627
rect 23765 22593 23799 22627
rect 27537 22593 27571 22627
rect 27721 22593 27755 22627
rect 27905 22593 27939 22627
rect 9965 22525 9999 22559
rect 13001 22525 13035 22559
rect 13921 22525 13955 22559
rect 14566 22525 14600 22559
rect 14749 22525 14783 22559
rect 17877 22525 17911 22559
rect 18337 22525 18371 22559
rect 20085 22525 20119 22559
rect 20361 22525 20395 22559
rect 22477 22525 22511 22559
rect 24501 22525 24535 22559
rect 28549 22525 28583 22559
rect 7665 22457 7699 22491
rect 8309 22389 8343 22423
rect 8585 22389 8619 22423
rect 9413 22389 9447 22423
rect 9873 22389 9907 22423
rect 12909 22389 12943 22423
rect 17417 22389 17451 22423
rect 17785 22389 17819 22423
rect 18705 22389 18739 22423
rect 19533 22389 19567 22423
rect 23949 22389 23983 22423
rect 29929 22389 29963 22423
rect 7665 22185 7699 22219
rect 12265 22185 12299 22219
rect 15301 22185 15335 22219
rect 15485 22185 15519 22219
rect 18613 22185 18647 22219
rect 13369 22117 13403 22151
rect 20637 22117 20671 22151
rect 7481 22049 7515 22083
rect 9413 22049 9447 22083
rect 9597 22049 9631 22083
rect 11713 22049 11747 22083
rect 13553 22049 13587 22083
rect 21557 22049 21591 22083
rect 24409 22049 24443 22083
rect 26249 22049 26283 22083
rect 26525 22049 26559 22083
rect 28549 22049 28583 22083
rect 29561 22049 29595 22083
rect 29929 22049 29963 22083
rect 7389 21981 7423 22015
rect 8217 21981 8251 22015
rect 8401 21981 8435 22015
rect 10642 21981 10676 22015
rect 11069 21981 11103 22015
rect 11161 21981 11195 22015
rect 11621 21981 11655 22015
rect 11805 21981 11839 22015
rect 12449 21981 12483 22015
rect 12541 21981 12575 22015
rect 12725 21981 12759 22015
rect 12817 21981 12851 22015
rect 13277 21981 13311 22015
rect 14105 21981 14139 22015
rect 14933 21981 14967 22015
rect 16405 21981 16439 22015
rect 16681 21981 16715 22015
rect 17233 21981 17267 22015
rect 17500 21981 17534 22015
rect 20821 21981 20855 22015
rect 22017 21981 22051 22015
rect 22110 21981 22144 22015
rect 22482 21981 22516 22015
rect 23121 21981 23155 22015
rect 23397 21981 23431 22015
rect 23489 21981 23523 22015
rect 24685 21981 24719 22015
rect 27537 21981 27571 22015
rect 27905 21981 27939 22015
rect 28733 21981 28767 22015
rect 29745 21981 29779 22015
rect 8309 21913 8343 21947
rect 9321 21913 9355 21947
rect 13553 21913 13587 21947
rect 21373 21913 21407 21947
rect 22293 21913 22327 21947
rect 22385 21913 22419 21947
rect 23305 21913 23339 21947
rect 27721 21913 27755 21947
rect 27813 21913 27847 21947
rect 8953 21845 8987 21879
rect 10517 21845 10551 21879
rect 10701 21845 10735 21879
rect 14197 21845 14231 21879
rect 15301 21845 15335 21879
rect 16681 21845 16715 21879
rect 22661 21845 22695 21879
rect 23673 21845 23707 21879
rect 28089 21845 28123 21879
rect 28917 21845 28951 21879
rect 10241 21641 10275 21675
rect 11713 21641 11747 21675
rect 14933 21641 14967 21675
rect 17049 21641 17083 21675
rect 17325 21641 17359 21675
rect 17877 21641 17911 21675
rect 23489 21641 23523 21675
rect 24317 21641 24351 21675
rect 26985 21641 27019 21675
rect 28181 21641 28215 21675
rect 14197 21573 14231 21607
rect 15945 21573 15979 21607
rect 17166 21573 17200 21607
rect 21097 21573 21131 21607
rect 22201 21573 22235 21607
rect 24869 21573 24903 21607
rect 26249 21573 26283 21607
rect 29070 21573 29104 21607
rect 7757 21505 7791 21539
rect 7941 21505 7975 21539
rect 8125 21505 8159 21539
rect 8309 21505 8343 21539
rect 9229 21505 9263 21539
rect 9321 21505 9355 21539
rect 9413 21505 9447 21539
rect 9597 21505 9631 21539
rect 10609 21505 10643 21539
rect 11710 21505 11744 21539
rect 13277 21505 13311 21539
rect 13369 21505 13403 21539
rect 13461 21505 13495 21539
rect 13645 21505 13679 21539
rect 14105 21505 14139 21539
rect 14749 21505 14783 21539
rect 16681 21505 16715 21539
rect 17785 21505 17819 21539
rect 19340 21505 19374 21539
rect 21833 21505 21867 21539
rect 21981 21505 22015 21539
rect 22109 21505 22143 21539
rect 22339 21505 22373 21539
rect 23305 21505 23339 21539
rect 23949 21505 23983 21539
rect 24133 21505 24167 21539
rect 25053 21505 25087 21539
rect 27353 21505 27387 21539
rect 27445 21505 27479 21539
rect 28365 21505 28399 21539
rect 8033 21437 8067 21471
rect 10701 21437 10735 21471
rect 10885 21437 10919 21471
rect 12173 21437 12207 21471
rect 15117 21437 15151 21471
rect 16957 21437 16991 21471
rect 19073 21437 19107 21471
rect 23121 21437 23155 21471
rect 27537 21437 27571 21471
rect 28825 21437 28859 21471
rect 11529 21369 11563 21403
rect 12081 21369 12115 21403
rect 16129 21369 16163 21403
rect 21281 21369 21315 21403
rect 8493 21301 8527 21335
rect 8953 21301 8987 21335
rect 13001 21301 13035 21335
rect 15117 21301 15151 21335
rect 20453 21301 20487 21335
rect 22477 21301 22511 21335
rect 26341 21301 26375 21335
rect 30205 21301 30239 21335
rect 8401 21097 8435 21131
rect 19257 21097 19291 21131
rect 21557 21097 21591 21131
rect 27077 21097 27111 21131
rect 28273 21097 28307 21131
rect 7757 20961 7791 20995
rect 9229 20961 9263 20995
rect 9505 20961 9539 20995
rect 10793 20961 10827 20995
rect 19625 20961 19659 20995
rect 25697 20961 25731 20995
rect 8125 20893 8159 20927
rect 8217 20893 8251 20927
rect 10517 20893 10551 20927
rect 12449 20893 12483 20927
rect 12817 20893 12851 20927
rect 12909 20893 12943 20927
rect 13369 20893 13403 20927
rect 14565 20893 14599 20927
rect 16865 20893 16899 20927
rect 19441 20893 19475 20927
rect 19717 20893 19751 20927
rect 20177 20893 20211 20927
rect 22017 20893 22051 20927
rect 22110 20893 22144 20927
rect 22385 20893 22419 20927
rect 22523 20893 22557 20927
rect 23213 20893 23247 20927
rect 23361 20893 23395 20927
rect 23489 20893 23523 20927
rect 23719 20893 23753 20927
rect 24409 20893 24443 20927
rect 24685 20893 24719 20927
rect 27721 20893 27755 20927
rect 27905 20893 27939 20927
rect 28089 20893 28123 20927
rect 28825 20893 28859 20927
rect 12541 20825 12575 20859
rect 12633 20825 12667 20859
rect 14832 20825 14866 20859
rect 17132 20825 17166 20859
rect 20444 20825 20478 20859
rect 22293 20825 22327 20859
rect 23581 20825 23615 20859
rect 25964 20825 25998 20859
rect 27997 20825 28031 20859
rect 12265 20757 12299 20791
rect 13461 20757 13495 20791
rect 15945 20757 15979 20791
rect 18245 20757 18279 20791
rect 22661 20757 22695 20791
rect 23857 20757 23891 20791
rect 28917 20757 28951 20791
rect 8033 20553 8067 20587
rect 9873 20553 9907 20587
rect 10701 20553 10735 20587
rect 12357 20553 12391 20587
rect 13093 20553 13127 20587
rect 15577 20553 15611 20587
rect 17141 20553 17175 20587
rect 25053 20553 25087 20587
rect 8760 20485 8794 20519
rect 11805 20485 11839 20519
rect 22100 20485 22134 20519
rect 25789 20485 25823 20519
rect 28181 20485 28215 20519
rect 6653 20417 6687 20451
rect 6920 20417 6954 20451
rect 8493 20417 8527 20451
rect 10609 20417 10643 20451
rect 10793 20417 10827 20451
rect 10885 20417 10919 20451
rect 12173 20417 12207 20451
rect 12265 20417 12299 20451
rect 13001 20417 13035 20451
rect 14453 20417 14487 20451
rect 17417 20417 17451 20451
rect 17509 20417 17543 20451
rect 17601 20417 17635 20451
rect 17785 20417 17819 20451
rect 18521 20417 18555 20451
rect 18797 20417 18831 20451
rect 19257 20417 19291 20451
rect 19513 20417 19547 20451
rect 21833 20417 21867 20451
rect 23673 20417 23707 20451
rect 23940 20417 23974 20451
rect 25513 20417 25547 20451
rect 25661 20417 25695 20451
rect 25878 20417 25912 20451
rect 25978 20417 26012 20451
rect 26985 20417 27019 20451
rect 27078 20417 27112 20451
rect 27261 20417 27295 20451
rect 27353 20417 27387 20451
rect 27450 20417 27484 20451
rect 14197 20349 14231 20383
rect 18337 20281 18371 20315
rect 23213 20281 23247 20315
rect 11989 20213 12023 20247
rect 12081 20213 12115 20247
rect 18705 20213 18739 20247
rect 20637 20213 20671 20247
rect 26157 20213 26191 20247
rect 27629 20213 27663 20247
rect 28273 20213 28307 20247
rect 9321 20009 9355 20043
rect 10149 20009 10183 20043
rect 12357 20009 12391 20043
rect 13001 20009 13035 20043
rect 13185 20009 13219 20043
rect 14749 20009 14783 20043
rect 17509 20009 17543 20043
rect 18705 20009 18739 20043
rect 19993 20009 20027 20043
rect 20821 20009 20855 20043
rect 22937 20009 22971 20043
rect 26157 20009 26191 20043
rect 26801 20009 26835 20043
rect 28825 20009 28859 20043
rect 11069 19941 11103 19975
rect 16221 19873 16255 19907
rect 18337 19873 18371 19907
rect 19533 19873 19567 19907
rect 21557 19873 21591 19907
rect 24777 19873 24811 19907
rect 9321 19805 9355 19839
rect 9505 19805 9539 19839
rect 10149 19805 10183 19839
rect 10793 19805 10827 19839
rect 10977 19805 11011 19839
rect 11253 19805 11287 19839
rect 11989 19805 12023 19839
rect 12081 19805 12115 19839
rect 12173 19805 12207 19839
rect 12817 19805 12851 19839
rect 13001 19805 13035 19839
rect 14105 19805 14139 19839
rect 15025 19805 15059 19839
rect 15117 19805 15151 19839
rect 15209 19805 15243 19839
rect 15393 19805 15427 19839
rect 15853 19805 15887 19839
rect 17141 19805 17175 19839
rect 17969 19805 18003 19839
rect 18153 19805 18187 19839
rect 18245 19805 18279 19839
rect 18521 19805 18555 19839
rect 19257 19805 19291 19839
rect 19441 19805 19475 19839
rect 19625 19805 19659 19839
rect 19809 19805 19843 19839
rect 20637 19805 20671 19839
rect 20913 19805 20947 19839
rect 21824 19805 21858 19839
rect 25044 19805 25078 19839
rect 27445 19805 27479 19839
rect 27712 19805 27746 19839
rect 16037 19737 16071 19771
rect 17325 19737 17359 19771
rect 26709 19737 26743 19771
rect 14197 19669 14231 19703
rect 20453 19669 20487 19703
rect 9413 19465 9447 19499
rect 12081 19465 12115 19499
rect 14289 19465 14323 19499
rect 26341 19465 26375 19499
rect 29009 19465 29043 19499
rect 12633 19397 12667 19431
rect 14933 19397 14967 19431
rect 16957 19397 16991 19431
rect 25973 19397 26007 19431
rect 10333 19329 10367 19363
rect 10425 19329 10459 19363
rect 10609 19329 10643 19363
rect 11529 19329 11563 19363
rect 11897 19329 11931 19363
rect 13461 19329 13495 19363
rect 14105 19329 14139 19363
rect 15761 19329 15795 19363
rect 15853 19329 15887 19363
rect 16129 19329 16163 19363
rect 16773 19329 16807 19363
rect 17877 19329 17911 19363
rect 19441 19329 19475 19363
rect 20545 19329 20579 19363
rect 20729 19329 20763 19363
rect 20821 19329 20855 19363
rect 21097 19329 21131 19363
rect 21925 19329 21959 19363
rect 22109 19329 22143 19363
rect 22201 19329 22235 19363
rect 22477 19329 22511 19363
rect 23949 19329 23983 19363
rect 25697 19329 25731 19363
rect 25790 19329 25824 19363
rect 26085 19329 26119 19363
rect 26203 19329 26237 19363
rect 27629 19329 27663 19363
rect 27885 19329 27919 19363
rect 9229 19261 9263 19295
rect 9597 19261 9631 19295
rect 10977 19261 11011 19295
rect 15577 19261 15611 19295
rect 17601 19261 17635 19295
rect 19165 19261 19199 19295
rect 20913 19261 20947 19295
rect 22293 19261 22327 19295
rect 23673 19261 23707 19295
rect 12817 19193 12851 19227
rect 9781 19125 9815 19159
rect 11621 19125 11655 19159
rect 13553 19125 13587 19159
rect 15025 19125 15059 19159
rect 16037 19125 16071 19159
rect 17141 19125 17175 19159
rect 21281 19125 21315 19159
rect 22661 19125 22695 19159
rect 11805 18921 11839 18955
rect 12265 18921 12299 18955
rect 17693 18921 17727 18955
rect 21097 18921 21131 18955
rect 27629 18921 27663 18955
rect 11989 18785 12023 18819
rect 16129 18785 16163 18819
rect 22477 18785 22511 18819
rect 10425 18717 10459 18751
rect 10701 18717 10735 18751
rect 11713 18717 11747 18751
rect 13093 18717 13127 18751
rect 13185 18717 13219 18751
rect 13277 18717 13311 18751
rect 13461 18717 13495 18751
rect 14565 18717 14599 18751
rect 14657 18717 14691 18751
rect 14770 18714 14804 18748
rect 14933 18717 14967 18751
rect 15761 18717 15795 18751
rect 16037 18717 16071 18751
rect 16865 18717 16899 18751
rect 16954 18714 16988 18748
rect 17049 18717 17083 18751
rect 17245 18717 17279 18751
rect 17923 18717 17957 18751
rect 18061 18717 18095 18751
rect 18153 18717 18187 18751
rect 18337 18717 18371 18751
rect 24501 18717 24535 18751
rect 26985 18717 27019 18751
rect 27133 18717 27167 18751
rect 27450 18717 27484 18751
rect 28273 18717 28307 18751
rect 28457 18717 28491 18751
rect 28549 18717 28583 18751
rect 19625 18649 19659 18683
rect 22722 18649 22756 18683
rect 24768 18649 24802 18683
rect 27261 18649 27295 18683
rect 27353 18649 27387 18683
rect 12817 18581 12851 18615
rect 14289 18581 14323 18615
rect 16589 18581 16623 18615
rect 23857 18581 23891 18615
rect 25881 18581 25915 18615
rect 28089 18581 28123 18615
rect 10057 18377 10091 18411
rect 10701 18377 10735 18411
rect 10609 18309 10643 18343
rect 17478 18309 17512 18343
rect 20076 18309 20110 18343
rect 26433 18309 26467 18343
rect 8677 18241 8711 18275
rect 8944 18241 8978 18275
rect 11529 18241 11563 18275
rect 13093 18241 13127 18275
rect 13185 18241 13219 18275
rect 13277 18241 13311 18275
rect 13461 18241 13495 18275
rect 14197 18241 14231 18275
rect 14289 18241 14323 18275
rect 14381 18241 14415 18275
rect 14565 18241 14599 18275
rect 15209 18241 15243 18275
rect 15761 18241 15795 18275
rect 19809 18241 19843 18275
rect 23121 18241 23155 18275
rect 23305 18241 23339 18275
rect 23673 18241 23707 18275
rect 24317 18241 24351 18275
rect 24501 18241 24535 18275
rect 24869 18241 24903 18275
rect 25701 18241 25735 18275
rect 25869 18241 25903 18275
rect 25973 18241 26007 18275
rect 26249 18241 26283 18275
rect 27252 18241 27286 18275
rect 28825 18241 28859 18275
rect 29009 18241 29043 18275
rect 12817 18173 12851 18207
rect 16037 18173 16071 18207
rect 17233 18173 17267 18207
rect 21833 18173 21867 18207
rect 22109 18173 22143 18207
rect 23397 18173 23431 18207
rect 23489 18173 23523 18207
rect 24593 18173 24627 18207
rect 24685 18173 24719 18207
rect 26065 18173 26099 18207
rect 26985 18173 27019 18207
rect 29285 18173 29319 18207
rect 15301 18105 15335 18139
rect 11713 18037 11747 18071
rect 13921 18037 13955 18071
rect 18613 18037 18647 18071
rect 21189 18037 21223 18071
rect 23857 18037 23891 18071
rect 25053 18037 25087 18071
rect 28365 18037 28399 18071
rect 29193 18037 29227 18071
rect 10333 17833 10367 17867
rect 19993 17833 20027 17867
rect 21833 17833 21867 17867
rect 22201 17833 22235 17867
rect 26433 17833 26467 17867
rect 8953 17697 8987 17731
rect 17417 17697 17451 17731
rect 18337 17697 18371 17731
rect 19625 17697 19659 17731
rect 20821 17697 20855 17731
rect 24685 17697 24719 17731
rect 24777 17697 24811 17731
rect 25973 17697 26007 17731
rect 27445 17697 27479 17731
rect 9220 17629 9254 17663
rect 11161 17629 11195 17663
rect 13185 17629 13219 17663
rect 13277 17629 13311 17663
rect 13369 17629 13403 17663
rect 13553 17629 13587 17663
rect 14105 17629 14139 17663
rect 14361 17629 14395 17663
rect 16221 17629 16255 17663
rect 16313 17629 16347 17663
rect 16497 17629 16531 17663
rect 16589 17629 16623 17663
rect 17233 17629 17267 17663
rect 17509 17629 17543 17663
rect 17969 17629 18003 17663
rect 18153 17629 18187 17663
rect 18248 17629 18282 17663
rect 18521 17629 18555 17663
rect 19257 17629 19291 17663
rect 19445 17629 19479 17663
rect 19533 17629 19567 17663
rect 19809 17629 19843 17663
rect 20545 17629 20579 17663
rect 22017 17629 22051 17663
rect 22293 17629 22327 17663
rect 22753 17629 22787 17663
rect 23029 17629 23063 17663
rect 24409 17629 24443 17663
rect 24593 17629 24627 17663
rect 24961 17629 24995 17663
rect 25697 17629 25731 17663
rect 25885 17629 25919 17663
rect 26065 17629 26099 17663
rect 26249 17629 26283 17663
rect 27712 17629 27746 17663
rect 11713 17561 11747 17595
rect 17049 17561 17083 17595
rect 10977 17493 11011 17527
rect 11805 17493 11839 17527
rect 12909 17493 12943 17527
rect 15485 17493 15519 17527
rect 16037 17493 16071 17527
rect 18705 17493 18739 17527
rect 25145 17493 25179 17527
rect 28825 17493 28859 17527
rect 10333 17289 10367 17323
rect 12725 17289 12759 17323
rect 15853 17289 15887 17323
rect 16037 17289 16071 17323
rect 20913 17289 20947 17323
rect 22063 17289 22097 17323
rect 25789 17289 25823 17323
rect 11989 17221 12023 17255
rect 28181 17221 28215 17255
rect 7849 17153 7883 17187
rect 8105 17153 8139 17187
rect 10517 17153 10551 17187
rect 11897 17153 11931 17187
rect 12081 17153 12115 17187
rect 12541 17153 12575 17187
rect 12725 17153 12759 17187
rect 14473 17153 14507 17187
rect 15761 17153 15795 17187
rect 16129 17143 16163 17177
rect 17509 17153 17543 17187
rect 17601 17153 17635 17187
rect 17693 17153 17727 17187
rect 17877 17153 17911 17187
rect 18889 17153 18923 17187
rect 20181 17163 20215 17197
rect 20361 17153 20395 17187
rect 20729 17153 20763 17187
rect 23305 17153 23339 17187
rect 23489 17153 23523 17187
rect 23949 17153 23983 17187
rect 24216 17153 24250 17187
rect 25973 17153 26007 17187
rect 26985 17153 27019 17187
rect 27169 17153 27203 17187
rect 27261 17153 27295 17187
rect 27537 17153 27571 17187
rect 28365 17153 28399 17187
rect 13185 17085 13219 17119
rect 13461 17085 13495 17119
rect 14749 17085 14783 17119
rect 15945 17085 15979 17119
rect 19165 17085 19199 17119
rect 20453 17085 20487 17119
rect 20545 17085 20579 17119
rect 21833 17085 21867 17119
rect 26249 17085 26283 17119
rect 27353 17085 27387 17119
rect 28641 17085 28675 17119
rect 28549 17017 28583 17051
rect 9229 16949 9263 16983
rect 17233 16949 17267 16983
rect 23305 16949 23339 16983
rect 25329 16949 25363 16983
rect 26157 16949 26191 16983
rect 27721 16949 27755 16983
rect 11989 16745 12023 16779
rect 15117 16745 15151 16779
rect 26893 16745 26927 16779
rect 9321 16677 9355 16711
rect 15945 16677 15979 16711
rect 10609 16609 10643 16643
rect 17325 16609 17359 16643
rect 19809 16609 19843 16643
rect 24869 16609 24903 16643
rect 26433 16609 26467 16643
rect 27629 16609 27663 16643
rect 8401 16541 8435 16575
rect 9137 16541 9171 16575
rect 10876 16541 10910 16575
rect 12633 16541 12667 16575
rect 13369 16541 13403 16575
rect 14105 16541 14139 16575
rect 14289 16541 14323 16575
rect 14933 16541 14967 16575
rect 15209 16541 15243 16575
rect 16037 16541 16071 16575
rect 17581 16541 17615 16575
rect 20065 16541 20099 16575
rect 21649 16541 21683 16575
rect 23489 16541 23523 16575
rect 25145 16541 25179 16575
rect 26157 16541 26191 16575
rect 26341 16541 26375 16575
rect 26525 16541 26559 16575
rect 26709 16541 26743 16575
rect 8953 16473 8987 16507
rect 13461 16473 13495 16507
rect 15669 16473 15703 16507
rect 16129 16473 16163 16507
rect 16681 16473 16715 16507
rect 16865 16473 16899 16507
rect 21916 16473 21950 16507
rect 27896 16473 27930 16507
rect 8217 16405 8251 16439
rect 12449 16405 12483 16439
rect 14289 16405 14323 16439
rect 14749 16405 14783 16439
rect 15761 16405 15795 16439
rect 18705 16405 18739 16439
rect 21189 16405 21223 16439
rect 23029 16405 23063 16439
rect 23581 16405 23615 16439
rect 29009 16405 29043 16439
rect 15853 16201 15887 16235
rect 17693 16201 17727 16235
rect 18521 16201 18555 16235
rect 28181 16201 28215 16235
rect 8116 16133 8150 16167
rect 11796 16133 11830 16167
rect 17325 16133 17359 16167
rect 18153 16133 18187 16167
rect 22652 16133 22686 16167
rect 7389 16065 7423 16099
rect 9689 16065 9723 16099
rect 9873 16065 9907 16099
rect 10793 16065 10827 16099
rect 10977 16065 11011 16099
rect 14933 16065 14967 16099
rect 15025 16065 15059 16099
rect 15117 16065 15151 16099
rect 15301 16065 15335 16099
rect 15761 16065 15795 16099
rect 16681 16065 16715 16099
rect 16865 16065 16899 16099
rect 17509 16065 17543 16099
rect 18337 16065 18371 16099
rect 19257 16065 19291 16099
rect 19441 16065 19475 16099
rect 19993 16065 20027 16099
rect 20269 16065 20303 16099
rect 24225 16065 24259 16099
rect 25789 16065 25823 16099
rect 26985 16065 27019 16099
rect 27169 16065 27203 16099
rect 27353 16065 27387 16099
rect 27537 16065 27571 16099
rect 28365 16065 28399 16099
rect 28641 16065 28675 16099
rect 7849 15997 7883 16031
rect 11529 15997 11563 16031
rect 13369 15997 13403 16031
rect 13645 15997 13679 16031
rect 19533 15997 19567 16031
rect 22385 15997 22419 16031
rect 24501 15997 24535 16031
rect 25513 15997 25547 16031
rect 27261 15997 27295 16031
rect 10057 15929 10091 15963
rect 10885 15929 10919 15963
rect 23765 15929 23799 15963
rect 7205 15861 7239 15895
rect 9229 15861 9263 15895
rect 12909 15861 12943 15895
rect 14657 15861 14691 15895
rect 16681 15861 16715 15895
rect 19073 15861 19107 15895
rect 27721 15861 27755 15895
rect 28549 15861 28583 15895
rect 8401 15657 8435 15691
rect 12633 15657 12667 15691
rect 12817 15657 12851 15691
rect 17509 15657 17543 15691
rect 17693 15657 17727 15691
rect 18337 15657 18371 15691
rect 21925 15657 21959 15691
rect 22569 15657 22603 15691
rect 22937 15657 22971 15691
rect 23581 15657 23615 15691
rect 16865 15589 16899 15623
rect 19625 15589 19659 15623
rect 21465 15589 21499 15623
rect 27813 15589 27847 15623
rect 28733 15589 28767 15623
rect 10333 15521 10367 15555
rect 23029 15521 23063 15555
rect 24777 15521 24811 15555
rect 26157 15521 26191 15555
rect 26433 15521 26467 15555
rect 27905 15521 27939 15555
rect 28825 15521 28859 15555
rect 7021 15453 7055 15487
rect 8953 15453 8987 15487
rect 13461 15453 13495 15487
rect 14637 15453 14671 15487
rect 14730 15450 14764 15484
rect 14841 15453 14875 15487
rect 15025 15453 15059 15487
rect 15485 15453 15519 15487
rect 20085 15453 20119 15487
rect 22109 15453 22143 15487
rect 22753 15453 22787 15487
rect 23489 15453 23523 15487
rect 24409 15453 24443 15487
rect 24581 15453 24615 15487
rect 24685 15453 24719 15487
rect 24961 15453 24995 15487
rect 27629 15453 27663 15487
rect 28549 15453 28583 15487
rect 7288 15385 7322 15419
rect 9137 15385 9171 15419
rect 10600 15385 10634 15419
rect 12449 15385 12483 15419
rect 15730 15385 15764 15419
rect 17325 15385 17359 15419
rect 18245 15385 18279 15419
rect 19441 15385 19475 15419
rect 20330 15385 20364 15419
rect 9321 15317 9355 15351
rect 11713 15317 11747 15351
rect 12649 15317 12683 15351
rect 13277 15317 13311 15351
rect 14381 15317 14415 15351
rect 17535 15317 17569 15351
rect 25145 15317 25179 15351
rect 27445 15317 27479 15351
rect 28365 15317 28399 15351
rect 7205 15113 7239 15147
rect 9229 15113 9263 15147
rect 10057 15113 10091 15147
rect 10793 15113 10827 15147
rect 11739 15113 11773 15147
rect 22201 15113 22235 15147
rect 25973 15113 26007 15147
rect 28365 15113 28399 15147
rect 9873 15045 9907 15079
rect 11529 15045 11563 15079
rect 12992 15045 13026 15079
rect 17509 15045 17543 15079
rect 27252 15045 27286 15079
rect 7389 14977 7423 15011
rect 8116 14977 8150 15011
rect 9689 14977 9723 15011
rect 10977 14977 11011 15011
rect 14565 14977 14599 15011
rect 14821 14977 14855 15011
rect 17141 14977 17175 15011
rect 17234 14977 17268 15011
rect 17417 14977 17451 15011
rect 17647 14977 17681 15011
rect 18337 14977 18371 15011
rect 18430 14977 18464 15011
rect 18613 14977 18647 15011
rect 18705 14977 18739 15011
rect 18802 14977 18836 15011
rect 19533 14977 19567 15011
rect 21005 14977 21039 15011
rect 22385 14977 22419 15011
rect 22661 14977 22695 15011
rect 23489 14977 23523 15011
rect 24133 14977 24167 15011
rect 24860 14977 24894 15011
rect 26985 14977 27019 15011
rect 7849 14909 7883 14943
rect 12725 14909 12759 14943
rect 19809 14909 19843 14943
rect 22569 14909 22603 14943
rect 24593 14909 24627 14943
rect 11897 14841 11931 14875
rect 14105 14841 14139 14875
rect 15945 14841 15979 14875
rect 18981 14841 19015 14875
rect 11713 14773 11747 14807
rect 17785 14773 17819 14807
rect 20821 14773 20855 14807
rect 23305 14773 23339 14807
rect 23949 14773 23983 14807
rect 7573 14569 7607 14603
rect 8217 14569 8251 14603
rect 9321 14569 9355 14603
rect 12633 14569 12667 14603
rect 13553 14569 13587 14603
rect 17877 14569 17911 14603
rect 23489 14569 23523 14603
rect 24869 14569 24903 14603
rect 25237 14569 25271 14603
rect 28089 14569 28123 14603
rect 17233 14501 17267 14535
rect 21281 14501 21315 14535
rect 10425 14433 10459 14467
rect 14105 14433 14139 14467
rect 19257 14433 19291 14467
rect 22477 14433 22511 14467
rect 25329 14433 25363 14467
rect 26709 14433 26743 14467
rect 7757 14365 7791 14399
rect 8401 14365 8435 14399
rect 9965 14365 9999 14399
rect 12541 14365 12575 14399
rect 12725 14365 12759 14399
rect 13185 14365 13219 14399
rect 13369 14365 13403 14399
rect 14372 14365 14406 14399
rect 15945 14365 15979 14399
rect 16589 14365 16623 14399
rect 16682 14365 16716 14399
rect 16957 14365 16991 14399
rect 17095 14365 17129 14399
rect 18705 14365 18739 14399
rect 19524 14365 19558 14399
rect 21097 14365 21131 14399
rect 21833 14365 21867 14399
rect 22017 14365 22051 14399
rect 22661 14365 22695 14399
rect 23397 14365 23431 14399
rect 25053 14365 25087 14399
rect 26976 14365 27010 14399
rect 8953 14297 8987 14331
rect 9137 14297 9171 14331
rect 10692 14297 10726 14331
rect 16865 14297 16899 14331
rect 17693 14297 17727 14331
rect 17893 14297 17927 14331
rect 21925 14297 21959 14331
rect 9781 14229 9815 14263
rect 11805 14229 11839 14263
rect 15485 14229 15519 14263
rect 16037 14229 16071 14263
rect 18061 14229 18095 14263
rect 18521 14229 18555 14263
rect 20637 14229 20671 14263
rect 22845 14229 22879 14263
rect 9229 14025 9263 14059
rect 10333 14025 10367 14059
rect 14105 14025 14139 14059
rect 15577 14025 15611 14059
rect 17049 14025 17083 14059
rect 26249 14025 26283 14059
rect 11529 13957 11563 13991
rect 11745 13957 11779 13991
rect 13737 13957 13771 13991
rect 16681 13957 16715 13991
rect 16897 13957 16931 13991
rect 17509 13957 17543 13991
rect 17725 13957 17759 13991
rect 20361 13957 20395 13991
rect 21189 13957 21223 13991
rect 22100 13957 22134 13991
rect 25973 13957 26007 13991
rect 7849 13889 7883 13923
rect 8116 13889 8150 13923
rect 10241 13889 10275 13923
rect 12633 13889 12667 13923
rect 12817 13889 12851 13923
rect 13921 13889 13955 13923
rect 14830 13889 14864 13923
rect 15853 13889 15887 13923
rect 16037 13889 16071 13923
rect 18521 13889 18555 13923
rect 19165 13889 19199 13923
rect 19257 13889 19291 13923
rect 19533 13889 19567 13923
rect 20177 13889 20211 13923
rect 21005 13889 21039 13923
rect 21833 13889 21867 13923
rect 23673 13889 23707 13923
rect 23940 13889 23974 13923
rect 25605 13889 25639 13923
rect 25698 13889 25732 13923
rect 25881 13889 25915 13923
rect 26070 13889 26104 13923
rect 27169 13889 27203 13923
rect 14750 13821 14784 13855
rect 14924 13821 14958 13855
rect 15025 13821 15059 13855
rect 15761 13821 15795 13855
rect 15945 13821 15979 13855
rect 18981 13821 19015 13855
rect 19993 13821 20027 13855
rect 20821 13821 20855 13855
rect 14565 13753 14599 13787
rect 11713 13685 11747 13719
rect 11897 13685 11931 13719
rect 12633 13685 12667 13719
rect 16865 13685 16899 13719
rect 17693 13685 17727 13719
rect 17877 13685 17911 13719
rect 18337 13685 18371 13719
rect 19441 13685 19475 13719
rect 23213 13685 23247 13719
rect 25053 13685 25087 13719
rect 26985 13685 27019 13719
rect 11805 13481 11839 13515
rect 12449 13481 12483 13515
rect 14289 13481 14323 13515
rect 16221 13481 16255 13515
rect 16405 13481 16439 13515
rect 17049 13481 17083 13515
rect 18153 13481 18187 13515
rect 19441 13481 19475 13515
rect 19625 13481 19659 13515
rect 27629 13481 27663 13515
rect 12633 13413 12667 13447
rect 14473 13413 14507 13447
rect 10425 13345 10459 13379
rect 24869 13345 24903 13379
rect 8401 13277 8435 13311
rect 13185 13277 13219 13311
rect 14105 13277 14139 13311
rect 14289 13277 14323 13311
rect 15393 13277 15427 13311
rect 20637 13277 20671 13311
rect 20785 13277 20819 13311
rect 21143 13277 21177 13311
rect 21833 13277 21867 13311
rect 21926 13277 21960 13311
rect 22201 13277 22235 13311
rect 22339 13277 22373 13311
rect 23213 13277 23247 13311
rect 23306 13277 23340 13311
rect 23678 13277 23712 13311
rect 25136 13277 25170 13311
rect 26801 13277 26835 13311
rect 28365 13277 28399 13311
rect 9321 13209 9355 13243
rect 9505 13209 9539 13243
rect 10692 13209 10726 13243
rect 12265 13209 12299 13243
rect 12465 13209 12499 13243
rect 13553 13209 13587 13243
rect 16037 13209 16071 13243
rect 16865 13209 16899 13243
rect 17969 13209 18003 13243
rect 18169 13209 18203 13243
rect 19257 13209 19291 13243
rect 19473 13209 19507 13243
rect 20913 13209 20947 13243
rect 21005 13209 21039 13243
rect 22109 13209 22143 13243
rect 23489 13209 23523 13243
rect 23581 13209 23615 13243
rect 26985 13209 27019 13243
rect 27537 13209 27571 13243
rect 8217 13141 8251 13175
rect 9689 13141 9723 13175
rect 15485 13141 15519 13175
rect 16237 13141 16271 13175
rect 17065 13141 17099 13175
rect 17233 13141 17267 13175
rect 18337 13141 18371 13175
rect 21281 13141 21315 13175
rect 22477 13141 22511 13175
rect 23857 13141 23891 13175
rect 26249 13141 26283 13175
rect 28181 13141 28215 13175
rect 7849 12937 7883 12971
rect 9873 12937 9907 12971
rect 10517 12937 10551 12971
rect 11897 12937 11931 12971
rect 13093 12937 13127 12971
rect 15961 12937 15995 12971
rect 16129 12937 16163 12971
rect 21281 12937 21315 12971
rect 23489 12937 23523 12971
rect 24317 12937 24351 12971
rect 28365 12937 28399 12971
rect 28825 12937 28859 12971
rect 11529 12869 11563 12903
rect 11745 12869 11779 12903
rect 15761 12869 15795 12903
rect 18613 12869 18647 12903
rect 18705 12869 18739 12903
rect 23305 12869 23339 12903
rect 25697 12869 25731 12903
rect 27252 12869 27286 12903
rect 8033 12801 8067 12835
rect 8493 12801 8527 12835
rect 8760 12801 8794 12835
rect 10701 12801 10735 12835
rect 13001 12801 13035 12835
rect 14013 12801 14047 12835
rect 14289 12801 14323 12835
rect 16681 12801 16715 12835
rect 18337 12801 18371 12835
rect 18485 12801 18519 12835
rect 18843 12801 18877 12835
rect 19901 12801 19935 12835
rect 20168 12801 20202 12835
rect 22477 12801 22511 12835
rect 23121 12801 23155 12835
rect 23949 12801 23983 12835
rect 24133 12801 24167 12835
rect 25329 12801 25363 12835
rect 25477 12801 25511 12835
rect 25605 12801 25639 12835
rect 25794 12801 25828 12835
rect 26985 12801 27019 12835
rect 29009 12801 29043 12835
rect 16957 12733 16991 12767
rect 22293 12733 22327 12767
rect 11713 12597 11747 12631
rect 15945 12597 15979 12631
rect 18981 12597 19015 12631
rect 22661 12597 22695 12631
rect 25973 12597 26007 12631
rect 9137 12393 9171 12427
rect 11805 12393 11839 12427
rect 13461 12393 13495 12427
rect 14381 12393 14415 12427
rect 14749 12393 14783 12427
rect 15761 12393 15795 12427
rect 21281 12393 21315 12427
rect 21465 12393 21499 12427
rect 23765 12393 23799 12427
rect 25605 12393 25639 12427
rect 28549 12393 28583 12427
rect 7573 12325 7607 12359
rect 14243 12325 14277 12359
rect 22661 12325 22695 12359
rect 13369 12257 13403 12291
rect 14473 12257 14507 12291
rect 15669 12257 15703 12291
rect 16865 12257 16899 12291
rect 17141 12257 17175 12291
rect 19809 12257 19843 12291
rect 26985 12257 27019 12291
rect 7757 12189 7791 12223
rect 8401 12189 8435 12223
rect 9321 12189 9355 12223
rect 9965 12189 9999 12223
rect 10425 12189 10459 12223
rect 10692 12189 10726 12223
rect 12541 12189 12575 12223
rect 13277 12189 13311 12223
rect 15485 12189 15519 12223
rect 15853 12189 15887 12223
rect 18521 12189 18555 12223
rect 20085 12189 20119 12223
rect 22385 12189 22419 12223
rect 22477 12189 22511 12223
rect 22753 12189 22787 12223
rect 24777 12189 24811 12223
rect 26249 12189 26283 12223
rect 26709 12189 26743 12223
rect 27997 12189 28031 12223
rect 28365 12189 28399 12223
rect 12357 12121 12391 12155
rect 13553 12121 13587 12155
rect 14105 12121 14139 12155
rect 18705 12121 18739 12155
rect 21123 12121 21157 12155
rect 23673 12121 23707 12155
rect 24409 12121 24443 12155
rect 24593 12121 24627 12155
rect 25237 12121 25271 12155
rect 25421 12121 25455 12155
rect 28181 12121 28215 12155
rect 28273 12121 28307 12155
rect 8217 12053 8251 12087
rect 9781 12053 9815 12087
rect 21297 12053 21331 12087
rect 22201 12053 22235 12087
rect 26065 12053 26099 12087
rect 10793 11849 10827 11883
rect 11529 11849 11563 11883
rect 12449 11849 12483 11883
rect 15025 11849 15059 11883
rect 19257 11849 19291 11883
rect 23305 11849 23339 11883
rect 26433 11849 26467 11883
rect 28365 11849 28399 11883
rect 12173 11781 12207 11815
rect 12357 11781 12391 11815
rect 13829 11781 13863 11815
rect 16037 11781 16071 11815
rect 17049 11781 17083 11815
rect 22192 11781 22226 11815
rect 26065 11781 26099 11815
rect 27252 11781 27286 11815
rect 6377 11713 6411 11747
rect 6633 11713 6667 11747
rect 8576 11713 8610 11747
rect 10977 11713 11011 11747
rect 11713 11713 11747 11747
rect 12449 11713 12483 11747
rect 12909 11713 12943 11747
rect 13093 11713 13127 11747
rect 14013 11713 14047 11747
rect 14105 11713 14139 11747
rect 15209 11713 15243 11747
rect 15485 11713 15519 11747
rect 15945 11713 15979 11747
rect 16865 11713 16899 11747
rect 17141 11713 17175 11747
rect 17877 11713 17911 11747
rect 18144 11713 18178 11747
rect 19717 11713 19751 11747
rect 19901 11713 19935 11747
rect 20269 11713 20303 11747
rect 21281 11713 21315 11747
rect 21925 11713 21959 11747
rect 25329 11713 25363 11747
rect 26249 11713 26283 11747
rect 29009 11713 29043 11747
rect 8309 11645 8343 11679
rect 19993 11645 20027 11679
rect 20085 11645 20119 11679
rect 23949 11645 23983 11679
rect 24225 11645 24259 11679
rect 25513 11645 25547 11679
rect 26985 11645 27019 11679
rect 14289 11577 14323 11611
rect 15393 11577 15427 11611
rect 20453 11577 20487 11611
rect 21097 11577 21131 11611
rect 7757 11509 7791 11543
rect 9689 11509 9723 11543
rect 13277 11509 13311 11543
rect 13829 11509 13863 11543
rect 16681 11509 16715 11543
rect 28825 11509 28859 11543
rect 7205 11305 7239 11339
rect 8033 11305 8067 11339
rect 12909 11305 12943 11339
rect 14197 11305 14231 11339
rect 14933 11305 14967 11339
rect 15485 11305 15519 11339
rect 21189 11305 21223 11339
rect 22569 11305 22603 11339
rect 27077 11305 27111 11339
rect 10241 11237 10275 11271
rect 19441 11237 19475 11271
rect 28273 11237 28307 11271
rect 29561 11237 29595 11271
rect 5825 11169 5859 11203
rect 7665 11169 7699 11203
rect 12541 11169 12575 11203
rect 12909 11169 12943 11203
rect 16957 11169 16991 11203
rect 17417 11169 17451 11203
rect 4813 11101 4847 11135
rect 5549 11101 5583 11135
rect 5641 11101 5675 11135
rect 6929 11101 6963 11135
rect 7024 11095 7058 11129
rect 7849 11101 7883 11135
rect 8953 11101 8987 11135
rect 9137 11101 9171 11135
rect 10425 11101 10459 11135
rect 10977 11101 11011 11135
rect 11897 11101 11931 11135
rect 14105 11101 14139 11135
rect 14289 11101 14323 11135
rect 15669 11101 15703 11135
rect 15853 11101 15887 11135
rect 16129 11101 16163 11135
rect 16589 11101 16623 11135
rect 16865 11101 16899 11135
rect 17601 11101 17635 11135
rect 17785 11101 17819 11135
rect 19257 11101 19291 11135
rect 20085 11101 20119 11135
rect 20233 11101 20267 11135
rect 20591 11101 20625 11135
rect 21373 11101 21407 11135
rect 23213 11101 23247 11135
rect 23306 11101 23340 11135
rect 23581 11101 23615 11135
rect 23678 11101 23712 11135
rect 24409 11101 24443 11135
rect 24676 11101 24710 11135
rect 26709 11101 26743 11135
rect 27629 11101 27663 11135
rect 28457 11101 28491 11135
rect 29745 11101 29779 11135
rect 9321 11033 9355 11067
rect 11161 11033 11195 11067
rect 12081 11033 12115 11067
rect 14841 11033 14875 11067
rect 15761 11033 15795 11067
rect 15991 11033 16025 11067
rect 18337 11033 18371 11067
rect 18521 11033 18555 11067
rect 20361 11033 20395 11067
rect 20453 11033 20487 11067
rect 22201 11033 22235 11067
rect 22385 11033 22419 11067
rect 23489 11033 23523 11067
rect 26893 11033 26927 11067
rect 27813 11033 27847 11067
rect 4629 10965 4663 10999
rect 12725 10965 12759 10999
rect 20729 10965 20763 10999
rect 23857 10965 23891 10999
rect 25789 10965 25823 10999
rect 6469 10761 6503 10795
rect 7665 10761 7699 10795
rect 23397 10761 23431 10795
rect 17877 10693 17911 10727
rect 24225 10693 24259 10727
rect 25053 10693 25087 10727
rect 26249 10693 26283 10727
rect 4905 10625 4939 10659
rect 5641 10625 5675 10659
rect 6653 10625 6687 10659
rect 7113 10625 7147 10659
rect 7297 10625 7331 10659
rect 7389 10625 7423 10659
rect 7481 10625 7515 10659
rect 8401 10625 8435 10659
rect 9117 10625 9151 10659
rect 10793 10625 10827 10659
rect 12081 10625 12115 10659
rect 13441 10625 13475 10659
rect 15669 10625 15703 10659
rect 15853 10625 15887 10659
rect 17141 10625 17175 10659
rect 18521 10625 18555 10659
rect 19625 10625 19659 10659
rect 19892 10625 19926 10659
rect 22017 10625 22051 10659
rect 22284 10625 22318 10659
rect 24869 10625 24903 10659
rect 25141 10625 25175 10659
rect 25283 10625 25317 10659
rect 27445 10625 27479 10659
rect 28273 10625 28307 10659
rect 28917 10625 28951 10659
rect 29377 10625 29411 10659
rect 29561 10625 29595 10659
rect 30205 10625 30239 10659
rect 30849 10625 30883 10659
rect 5457 10557 5491 10591
rect 5825 10557 5859 10591
rect 8861 10557 8895 10591
rect 13185 10557 13219 10591
rect 18613 10557 18647 10591
rect 24409 10557 24443 10591
rect 27629 10557 27663 10591
rect 10977 10489 11011 10523
rect 14565 10489 14599 10523
rect 17325 10489 17359 10523
rect 21005 10489 21039 10523
rect 28733 10489 28767 10523
rect 30021 10489 30055 10523
rect 4721 10421 4755 10455
rect 8217 10421 8251 10455
rect 10241 10421 10275 10455
rect 12173 10421 12207 10455
rect 17969 10421 18003 10455
rect 25421 10421 25455 10455
rect 26341 10421 26375 10455
rect 28089 10421 28123 10455
rect 29377 10421 29411 10455
rect 30665 10421 30699 10455
rect 6377 10217 6411 10251
rect 7665 10217 7699 10251
rect 8125 10217 8159 10251
rect 12817 10217 12851 10251
rect 17233 10217 17267 10251
rect 20085 10217 20119 10251
rect 21005 10217 21039 10251
rect 23489 10217 23523 10251
rect 27169 10217 27203 10251
rect 9183 10149 9217 10183
rect 20269 10149 20303 10183
rect 22017 10149 22051 10183
rect 29561 10149 29595 10183
rect 12449 10081 12483 10115
rect 17877 10081 17911 10115
rect 18153 10081 18187 10115
rect 27629 10081 27663 10115
rect 3985 10013 4019 10047
rect 4252 10013 4286 10047
rect 5825 10013 5859 10047
rect 6009 10013 6043 10047
rect 6193 10013 6227 10047
rect 7113 10013 7147 10047
rect 7297 10013 7331 10047
rect 7481 10013 7515 10047
rect 8309 10013 8343 10047
rect 8953 10013 8987 10047
rect 10609 10013 10643 10047
rect 12633 10013 12667 10047
rect 13369 10013 13403 10047
rect 14473 10013 14507 10047
rect 14841 10013 14875 10047
rect 15853 10013 15887 10047
rect 19263 10013 19297 10047
rect 19441 10013 19475 10047
rect 22201 10013 22235 10047
rect 22845 10013 22879 10047
rect 23397 10013 23431 10047
rect 24961 10013 24995 10047
rect 25145 10013 25179 10047
rect 25789 10013 25823 10047
rect 27896 10013 27930 10047
rect 29745 10013 29779 10047
rect 30389 10013 30423 10047
rect 31217 10013 31251 10047
rect 6101 9945 6135 9979
rect 7389 9945 7423 9979
rect 10854 9945 10888 9979
rect 13553 9945 13587 9979
rect 14657 9945 14691 9979
rect 14749 9945 14783 9979
rect 16120 9945 16154 9979
rect 19901 9945 19935 9979
rect 20821 9945 20855 9979
rect 21037 9945 21071 9979
rect 26056 9945 26090 9979
rect 5365 9877 5399 9911
rect 11989 9877 12023 9911
rect 15025 9877 15059 9911
rect 19349 9877 19383 9911
rect 20111 9877 20145 9911
rect 21189 9877 21223 9911
rect 22661 9877 22695 9911
rect 25329 9877 25363 9911
rect 29009 9877 29043 9911
rect 30205 9877 30239 9911
rect 31033 9877 31067 9911
rect 7757 9673 7791 9707
rect 25513 9673 25547 9707
rect 26985 9673 27019 9707
rect 10977 9605 11011 9639
rect 11805 9605 11839 9639
rect 12909 9605 12943 9639
rect 14289 9605 14323 9639
rect 18061 9605 18095 9639
rect 23397 9605 23431 9639
rect 23581 9605 23615 9639
rect 25145 9605 25179 9639
rect 25237 9605 25271 9639
rect 28181 9605 28215 9639
rect 3893 9537 3927 9571
rect 4160 9537 4194 9571
rect 6377 9537 6411 9571
rect 6644 9537 6678 9571
rect 9025 9537 9059 9571
rect 10609 9537 10643 9571
rect 10793 9537 10827 9571
rect 11621 9537 11655 9571
rect 11897 9537 11931 9571
rect 11989 9537 12023 9571
rect 12725 9537 12759 9571
rect 14105 9537 14139 9571
rect 15301 9537 15335 9571
rect 17877 9537 17911 9571
rect 18153 9537 18187 9571
rect 18705 9537 18739 9571
rect 20269 9537 20303 9571
rect 20361 9537 20395 9571
rect 20637 9537 20671 9571
rect 21281 9537 21315 9571
rect 22477 9537 22511 9571
rect 22569 9537 22603 9571
rect 22845 9537 22879 9571
rect 24225 9537 24259 9571
rect 24961 9537 24995 9571
rect 25329 9537 25363 9571
rect 26157 9537 26191 9571
rect 27169 9537 27203 9571
rect 27905 9537 27939 9571
rect 28089 9537 28123 9571
rect 28365 9537 28399 9571
rect 28641 9537 28675 9571
rect 29285 9537 29319 9571
rect 29929 9537 29963 9571
rect 30573 9537 30607 9571
rect 31217 9537 31251 9571
rect 8769 9469 8803 9503
rect 13921 9469 13955 9503
rect 15577 9469 15611 9503
rect 16681 9469 16715 9503
rect 18981 9469 19015 9503
rect 24041 9469 24075 9503
rect 24409 9469 24443 9503
rect 12173 9401 12207 9435
rect 17049 9401 17083 9435
rect 21097 9401 21131 9435
rect 22293 9401 22327 9435
rect 29101 9401 29135 9435
rect 30389 9401 30423 9435
rect 5273 9333 5307 9367
rect 10149 9333 10183 9367
rect 17141 9333 17175 9367
rect 17877 9333 17911 9367
rect 18981 9333 19015 9367
rect 19257 9333 19291 9367
rect 20085 9333 20119 9367
rect 20545 9333 20579 9367
rect 22753 9333 22787 9367
rect 25973 9333 26007 9367
rect 29745 9333 29779 9367
rect 31033 9333 31067 9367
rect 6929 9129 6963 9163
rect 8033 9129 8067 9163
rect 18705 9129 18739 9163
rect 21189 9129 21223 9163
rect 23489 9129 23523 9163
rect 29837 9129 29871 9163
rect 25789 9061 25823 9095
rect 31033 9061 31067 9095
rect 9229 8993 9263 9027
rect 16681 8993 16715 9027
rect 24409 8993 24443 9027
rect 3249 8925 3283 8959
rect 4537 8925 4571 8959
rect 5181 8925 5215 8959
rect 5365 8925 5399 8959
rect 5549 8925 5583 8959
rect 5825 8925 5859 8959
rect 5917 8925 5951 8959
rect 6377 8925 6411 8959
rect 6653 8925 6687 8959
rect 6745 8925 6779 8959
rect 7481 8925 7515 8959
rect 7849 8925 7883 8959
rect 8953 8925 8987 8959
rect 10333 8925 10367 8959
rect 12173 8925 12207 8959
rect 14105 8925 14139 8959
rect 15117 8925 15151 8959
rect 15393 8925 15427 8959
rect 16497 8925 16531 8959
rect 16773 8925 16807 8959
rect 17325 8925 17359 8959
rect 19809 8925 19843 8959
rect 22109 8925 22143 8959
rect 24676 8925 24710 8959
rect 26249 8925 26283 8959
rect 26617 8925 26651 8959
rect 27813 8925 27847 8959
rect 28089 8925 28123 8959
rect 28365 8925 28399 8959
rect 28641 8925 28675 8959
rect 29653 8925 29687 8959
rect 30573 8925 30607 8959
rect 31217 8925 31251 8959
rect 31861 8925 31895 8959
rect 6561 8857 6595 8891
rect 7665 8857 7699 8891
rect 7757 8857 7791 8891
rect 10578 8857 10612 8891
rect 12440 8857 12474 8891
rect 16865 8857 16899 8891
rect 17592 8857 17626 8891
rect 20076 8857 20110 8891
rect 22376 8857 22410 8891
rect 26433 8857 26467 8891
rect 26525 8857 26559 8891
rect 28181 8857 28215 8891
rect 3065 8789 3099 8823
rect 4353 8789 4387 8823
rect 11713 8789 11747 8823
rect 13553 8789 13587 8823
rect 14289 8789 14323 8823
rect 14933 8789 14967 8823
rect 15301 8789 15335 8823
rect 26801 8789 26835 8823
rect 30389 8789 30423 8823
rect 31677 8789 31711 8823
rect 3709 8585 3743 8619
rect 4353 8585 4387 8619
rect 5641 8585 5675 8619
rect 9505 8585 9539 8619
rect 10333 8585 10367 8619
rect 11897 8585 11931 8619
rect 13921 8585 13955 8619
rect 19257 8585 19291 8619
rect 24501 8585 24535 8619
rect 26341 8585 26375 8619
rect 28733 8585 28767 8619
rect 29193 8585 29227 8619
rect 31125 8585 31159 8619
rect 32965 8585 32999 8619
rect 9137 8517 9171 8551
rect 11713 8517 11747 8551
rect 14841 8517 14875 8551
rect 19901 8517 19935 8551
rect 20269 8517 20303 8551
rect 24133 8517 24167 8551
rect 24225 8517 24259 8551
rect 27620 8517 27654 8551
rect 29929 8517 29963 8551
rect 1593 8449 1627 8483
rect 3893 8449 3927 8483
rect 4537 8449 4571 8483
rect 4997 8449 5031 8483
rect 5181 8449 5215 8483
rect 5825 8449 5859 8483
rect 6653 8449 6687 8483
rect 7113 8449 7147 8483
rect 7389 8449 7423 8483
rect 8309 8449 8343 8483
rect 9321 8449 9355 8483
rect 9965 8449 9999 8483
rect 10149 8449 10183 8483
rect 10793 8449 10827 8483
rect 10977 8449 11011 8483
rect 11529 8449 11563 8483
rect 12725 8449 12759 8483
rect 12909 8449 12943 8483
rect 13553 8449 13587 8483
rect 13737 8449 13771 8483
rect 15669 8449 15703 8483
rect 15853 8449 15887 8483
rect 17141 8449 17175 8483
rect 17233 8449 17267 8483
rect 17877 8449 17911 8483
rect 18144 8449 18178 8483
rect 20085 8449 20119 8483
rect 20913 8449 20947 8483
rect 22100 8449 22134 8483
rect 23949 8449 23983 8483
rect 24317 8449 24351 8483
rect 24961 8449 24995 8483
rect 25228 8449 25262 8483
rect 27353 8449 27387 8483
rect 29377 8449 29411 8483
rect 29837 8449 29871 8483
rect 30021 8449 30055 8483
rect 30665 8449 30699 8483
rect 31309 8449 31343 8483
rect 32505 8449 32539 8483
rect 33149 8449 33183 8483
rect 33968 8449 34002 8483
rect 5089 8381 5123 8415
rect 7297 8381 7331 8415
rect 17417 8381 17451 8415
rect 21833 8381 21867 8415
rect 33701 8381 33735 8415
rect 7573 8313 7607 8347
rect 8125 8313 8159 8347
rect 10885 8313 10919 8347
rect 15025 8313 15059 8347
rect 15853 8313 15887 8347
rect 20729 8313 20763 8347
rect 30481 8313 30515 8347
rect 32321 8313 32355 8347
rect 1409 8245 1443 8279
rect 6469 8245 6503 8279
rect 7113 8245 7147 8279
rect 13093 8245 13127 8279
rect 23213 8245 23247 8279
rect 35081 8245 35115 8279
rect 9965 8041 9999 8075
rect 10425 8041 10459 8075
rect 10977 8041 11011 8075
rect 11437 8041 11471 8075
rect 13001 8041 13035 8075
rect 16129 8041 16163 8075
rect 16589 8041 16623 8075
rect 17509 8041 17543 8075
rect 18061 8041 18095 8075
rect 19809 8041 19843 8075
rect 21925 8041 21959 8075
rect 22293 8041 22327 8075
rect 23213 8041 23247 8075
rect 31493 8041 31527 8075
rect 34713 8041 34747 8075
rect 2697 7973 2731 8007
rect 9413 7973 9447 8007
rect 25421 7973 25455 8007
rect 30205 7973 30239 8007
rect 2329 7905 2363 7939
rect 8953 7905 8987 7939
rect 11989 7905 12023 7939
rect 12449 7905 12483 7939
rect 13461 7905 13495 7939
rect 14473 7905 14507 7939
rect 14749 7905 14783 7939
rect 22385 7905 22419 7939
rect 26985 7905 27019 7939
rect 1685 7837 1719 7871
rect 1777 7837 1811 7871
rect 1961 7837 1995 7871
rect 3249 7837 3283 7871
rect 4261 7837 4295 7871
rect 5457 7837 5491 7871
rect 6101 7837 6135 7871
rect 7021 7837 7055 7871
rect 7481 7837 7515 7871
rect 7757 7837 7791 7871
rect 9137 7837 9171 7871
rect 9229 7837 9263 7871
rect 9505 7837 9539 7871
rect 10149 7837 10183 7871
rect 10241 7837 10275 7871
rect 10517 7837 10551 7871
rect 11161 7837 11195 7871
rect 11253 7837 11287 7871
rect 11529 7837 11563 7871
rect 12173 7837 12207 7871
rect 12265 7837 12299 7871
rect 12541 7837 12575 7871
rect 13185 7837 13219 7871
rect 13277 7837 13311 7871
rect 13553 7837 13587 7871
rect 16589 7837 16623 7871
rect 16865 7837 16899 7871
rect 17417 7837 17451 7871
rect 18061 7837 18095 7871
rect 18245 7837 18279 7871
rect 18337 7837 18371 7871
rect 20453 7837 20487 7871
rect 21097 7837 21131 7871
rect 22109 7837 22143 7871
rect 22937 7837 22971 7871
rect 23029 7837 23063 7871
rect 23857 7837 23891 7871
rect 24593 7837 24627 7871
rect 25145 7837 25179 7871
rect 25237 7837 25271 7871
rect 26065 7837 26099 7871
rect 26801 7837 26835 7871
rect 27077 7837 27111 7871
rect 27261 7837 27295 7871
rect 27537 7837 27571 7871
rect 29009 7837 29043 7871
rect 29561 7837 29595 7871
rect 29745 7837 29779 7871
rect 30389 7837 30423 7871
rect 31033 7837 31067 7871
rect 31677 7837 31711 7871
rect 32321 7837 32355 7871
rect 34897 7837 34931 7871
rect 35173 7837 35207 7871
rect 35817 7837 35851 7871
rect 36093 7837 36127 7871
rect 4445 7769 4479 7803
rect 15761 7769 15795 7803
rect 15945 7769 15979 7803
rect 16773 7769 16807 7803
rect 19441 7769 19475 7803
rect 19625 7769 19659 7803
rect 28181 7769 28215 7803
rect 28365 7769 28399 7803
rect 32588 7769 32622 7803
rect 4629 7701 4663 7735
rect 5273 7701 5307 7735
rect 5917 7701 5951 7735
rect 6837 7701 6871 7735
rect 20269 7701 20303 7735
rect 20913 7701 20947 7735
rect 23673 7701 23707 7735
rect 24409 7701 24443 7735
rect 25881 7701 25915 7735
rect 28825 7701 28859 7735
rect 29653 7701 29687 7735
rect 30849 7701 30883 7735
rect 33701 7701 33735 7735
rect 35081 7701 35115 7735
rect 35633 7701 35667 7735
rect 36001 7701 36035 7735
rect 1409 7497 1443 7531
rect 2329 7497 2363 7531
rect 2973 7497 3007 7531
rect 5457 7497 5491 7531
rect 15485 7497 15519 7531
rect 22385 7497 22419 7531
rect 25789 7497 25823 7531
rect 28365 7497 28399 7531
rect 29423 7497 29457 7531
rect 30681 7497 30715 7531
rect 30849 7497 30883 7531
rect 32873 7497 32907 7531
rect 33241 7497 33275 7531
rect 35173 7497 35207 7531
rect 8484 7429 8518 7463
rect 12142 7429 12176 7463
rect 18337 7429 18371 7463
rect 21097 7429 21131 7463
rect 22201 7429 22235 7463
rect 27252 7429 27286 7463
rect 30481 7429 30515 7463
rect 34060 7429 34094 7463
rect 1593 7361 1627 7395
rect 2513 7361 2547 7395
rect 3157 7361 3191 7395
rect 3884 7361 3918 7395
rect 5641 7361 5675 7395
rect 6377 7361 6411 7395
rect 6633 7361 6667 7395
rect 8217 7361 8251 7395
rect 10333 7361 10367 7395
rect 11897 7361 11931 7395
rect 15669 7361 15703 7395
rect 15761 7361 15795 7395
rect 16037 7361 16071 7395
rect 16957 7361 16991 7395
rect 18245 7361 18279 7395
rect 19533 7361 19567 7395
rect 20913 7361 20947 7395
rect 22017 7361 22051 7395
rect 23029 7361 23063 7395
rect 23673 7361 23707 7395
rect 24317 7361 24351 7395
rect 24409 7361 24443 7395
rect 24685 7361 24719 7395
rect 25329 7361 25363 7395
rect 25973 7361 26007 7395
rect 26985 7361 27019 7395
rect 29193 7361 29227 7395
rect 31493 7361 31527 7395
rect 32413 7361 32447 7395
rect 33057 7361 33091 7395
rect 33333 7361 33367 7395
rect 35817 7361 35851 7395
rect 36461 7361 36495 7395
rect 3617 7293 3651 7327
rect 10057 7293 10091 7327
rect 14197 7293 14231 7327
rect 14473 7293 14507 7327
rect 17233 7293 17267 7327
rect 19257 7293 19291 7327
rect 21281 7293 21315 7327
rect 33793 7293 33827 7327
rect 4997 7225 5031 7259
rect 15945 7225 15979 7259
rect 23489 7225 23523 7259
rect 25145 7225 25179 7259
rect 36277 7225 36311 7259
rect 7757 7157 7791 7191
rect 9597 7157 9631 7191
rect 13277 7157 13311 7191
rect 22845 7157 22879 7191
rect 24133 7157 24167 7191
rect 24593 7157 24627 7191
rect 30665 7157 30699 7191
rect 31309 7157 31343 7191
rect 32229 7157 32263 7191
rect 35633 7157 35667 7191
rect 1777 6953 1811 6987
rect 3065 6953 3099 6987
rect 9229 6953 9263 6987
rect 9413 6953 9447 6987
rect 11713 6953 11747 6987
rect 13001 6953 13035 6987
rect 16405 6953 16439 6987
rect 28733 6953 28767 6987
rect 33885 6953 33919 6987
rect 34897 6953 34931 6987
rect 5181 6885 5215 6919
rect 13185 6885 13219 6919
rect 18429 6885 18463 6919
rect 24869 6885 24903 6919
rect 32229 6885 32263 6919
rect 35633 6885 35667 6919
rect 3801 6817 3835 6851
rect 5641 6817 5675 6851
rect 6101 6817 6135 6851
rect 6929 6817 6963 6851
rect 9045 6817 9079 6851
rect 10333 6817 10367 6851
rect 1961 6749 1995 6783
rect 2605 6749 2639 6783
rect 3249 6749 3283 6783
rect 4068 6749 4102 6783
rect 5825 6749 5859 6783
rect 5917 6749 5951 6783
rect 6193 6749 6227 6783
rect 7205 6749 7239 6783
rect 8401 6749 8435 6783
rect 9229 6749 9263 6783
rect 12909 6749 12943 6783
rect 13001 6749 13035 6783
rect 14105 6749 14139 6783
rect 16129 6749 16163 6783
rect 16221 6749 16255 6783
rect 16497 6749 16531 6783
rect 17049 6749 17083 6783
rect 19257 6749 19291 6783
rect 19901 6749 19935 6783
rect 21833 6749 21867 6783
rect 22100 6749 22134 6783
rect 23857 6749 23891 6783
rect 24593 6749 24627 6783
rect 24685 6749 24719 6783
rect 24961 6749 24995 6783
rect 25605 6749 25639 6783
rect 26249 6749 26283 6783
rect 26893 6749 26927 6783
rect 28089 6749 28123 6783
rect 29745 6749 29779 6783
rect 31769 6749 31803 6783
rect 32413 6749 32447 6783
rect 33425 6749 33459 6783
rect 34069 6749 34103 6783
rect 35817 6749 35851 6783
rect 36461 6749 36495 6783
rect 8953 6681 8987 6715
rect 10600 6681 10634 6715
rect 12725 6681 12759 6715
rect 14372 6681 14406 6715
rect 17316 6681 17350 6715
rect 20168 6681 20202 6715
rect 28549 6681 28583 6715
rect 28754 6681 28788 6715
rect 30012 6681 30046 6715
rect 34713 6681 34747 6715
rect 2421 6613 2455 6647
rect 8217 6613 8251 6647
rect 15485 6613 15519 6647
rect 15945 6613 15979 6647
rect 19349 6613 19383 6647
rect 21281 6613 21315 6647
rect 23213 6613 23247 6647
rect 23673 6613 23707 6647
rect 24409 6613 24443 6647
rect 25421 6613 25455 6647
rect 26065 6613 26099 6647
rect 26709 6613 26743 6647
rect 27905 6613 27939 6647
rect 28917 6613 28951 6647
rect 31125 6613 31159 6647
rect 31585 6613 31619 6647
rect 33241 6613 33275 6647
rect 34913 6613 34947 6647
rect 35081 6613 35115 6647
rect 36277 6613 36311 6647
rect 1777 6409 1811 6443
rect 3065 6409 3099 6443
rect 3709 6409 3743 6443
rect 5825 6409 5859 6443
rect 9597 6409 9631 6443
rect 10609 6409 10643 6443
rect 12817 6409 12851 6443
rect 14289 6409 14323 6443
rect 36185 6409 36219 6443
rect 5457 6341 5491 6375
rect 6377 6341 6411 6375
rect 7665 6341 7699 6375
rect 8585 6341 8619 6375
rect 11529 6341 11563 6375
rect 13829 6341 13863 6375
rect 18420 6341 18454 6375
rect 34244 6341 34278 6375
rect 35817 6341 35851 6375
rect 36017 6341 36051 6375
rect 1961 6273 1995 6307
rect 2421 6273 2455 6307
rect 2697 6273 2731 6307
rect 3249 6273 3283 6307
rect 3893 6273 3927 6307
rect 4537 6273 4571 6307
rect 4629 6273 4663 6307
rect 4905 6273 4939 6307
rect 5641 6273 5675 6307
rect 6561 6273 6595 6307
rect 6653 6273 6687 6307
rect 6929 6273 6963 6307
rect 7481 6273 7515 6307
rect 8769 6273 8803 6307
rect 9781 6273 9815 6307
rect 9873 6273 9907 6307
rect 10149 6273 10183 6307
rect 10793 6273 10827 6307
rect 11805 6273 11839 6307
rect 13001 6273 13035 6307
rect 13093 6273 13127 6307
rect 13369 6273 13403 6307
rect 14105 6273 14139 6307
rect 14749 6273 14783 6307
rect 15016 6273 15050 6307
rect 20453 6273 20487 6307
rect 22293 6273 22327 6307
rect 22560 6273 22594 6307
rect 24133 6273 24167 6307
rect 24317 6273 24351 6307
rect 24961 6273 24995 6307
rect 25228 6273 25262 6307
rect 27445 6273 27479 6307
rect 27712 6273 27746 6307
rect 29285 6273 29319 6307
rect 29552 6273 29586 6307
rect 31309 6273 31343 6307
rect 32404 6273 32438 6307
rect 33977 6273 34011 6307
rect 37473 6273 37507 6307
rect 8953 6205 8987 6239
rect 11621 6205 11655 6239
rect 13921 6205 13955 6239
rect 16681 6205 16715 6239
rect 16957 6205 16991 6239
rect 18153 6205 18187 6239
rect 20729 6205 20763 6239
rect 32137 6205 32171 6239
rect 11989 6137 12023 6171
rect 13277 6137 13311 6171
rect 19533 6137 19567 6171
rect 23673 6137 23707 6171
rect 2237 6069 2271 6103
rect 4353 6069 4387 6103
rect 4813 6069 4847 6103
rect 6837 6069 6871 6103
rect 10057 6069 10091 6103
rect 11529 6069 11563 6103
rect 13829 6069 13863 6103
rect 16129 6069 16163 6103
rect 24501 6069 24535 6103
rect 26341 6069 26375 6103
rect 28825 6069 28859 6103
rect 30665 6069 30699 6103
rect 31125 6069 31159 6103
rect 33517 6069 33551 6103
rect 35357 6069 35391 6103
rect 36001 6069 36035 6103
rect 37289 6069 37323 6103
rect 1593 5865 1627 5899
rect 4537 5865 4571 5899
rect 8033 5865 8067 5899
rect 11989 5865 12023 5899
rect 15485 5865 15519 5899
rect 16589 5865 16623 5899
rect 19349 5865 19383 5899
rect 21005 5865 21039 5899
rect 23857 5865 23891 5899
rect 26617 5865 26651 5899
rect 33425 5865 33459 5899
rect 33609 5865 33643 5899
rect 34897 5865 34931 5899
rect 35081 5865 35115 5899
rect 3065 5797 3099 5831
rect 10609 5797 10643 5831
rect 12173 5797 12207 5831
rect 15669 5797 15703 5831
rect 17877 5797 17911 5831
rect 21465 5797 21499 5831
rect 22569 5797 22603 5831
rect 36277 5797 36311 5831
rect 11805 5729 11839 5763
rect 15301 5729 15335 5763
rect 17417 5729 17451 5763
rect 18613 5729 18647 5763
rect 19809 5729 19843 5763
rect 27537 5729 27571 5763
rect 31953 5729 31987 5763
rect 1777 5661 1811 5695
rect 2145 5661 2179 5695
rect 2605 5661 2639 5695
rect 3249 5637 3283 5671
rect 4169 5661 4203 5695
rect 5733 5661 5767 5695
rect 6561 5661 6595 5695
rect 7849 5661 7883 5695
rect 9229 5661 9263 5695
rect 11253 5661 11287 5695
rect 11713 5661 11747 5695
rect 11989 5661 12023 5695
rect 12909 5661 12943 5695
rect 13553 5661 13587 5695
rect 14289 5661 14323 5695
rect 14473 5661 14507 5695
rect 15485 5661 15519 5695
rect 17142 5661 17176 5695
rect 17234 5661 17268 5695
rect 17509 5661 17543 5695
rect 18337 5661 18371 5695
rect 18429 5661 18463 5695
rect 18705 5661 18739 5695
rect 19533 5661 19567 5695
rect 19625 5661 19659 5695
rect 19901 5661 19935 5695
rect 20545 5661 20579 5695
rect 21189 5661 21223 5695
rect 21281 5661 21315 5695
rect 21557 5661 21591 5695
rect 22293 5661 22327 5695
rect 22385 5661 22419 5695
rect 22661 5661 22695 5695
rect 23489 5661 23523 5695
rect 24409 5661 24443 5695
rect 25237 5661 25271 5695
rect 27813 5661 27847 5695
rect 29009 5661 29043 5695
rect 30113 5661 30147 5695
rect 32229 5661 32263 5695
rect 35725 5661 35759 5695
rect 36461 5661 36495 5695
rect 37105 5661 37139 5695
rect 37749 5661 37783 5695
rect 4353 5593 4387 5627
rect 6193 5593 6227 5627
rect 6377 5593 6411 5627
rect 7205 5593 7239 5627
rect 9496 5593 9530 5627
rect 14105 5593 14139 5627
rect 15209 5593 15243 5627
rect 16313 5593 16347 5627
rect 22109 5593 22143 5627
rect 23673 5593 23707 5627
rect 24593 5593 24627 5627
rect 24777 5593 24811 5627
rect 25504 5593 25538 5627
rect 30380 5593 30414 5627
rect 33241 5593 33275 5627
rect 33457 5593 33491 5627
rect 34713 5593 34747 5627
rect 2421 5525 2455 5559
rect 5549 5525 5583 5559
rect 7297 5525 7331 5559
rect 11069 5525 11103 5559
rect 12725 5525 12759 5559
rect 13369 5525 13403 5559
rect 16957 5525 16991 5559
rect 18153 5525 18187 5559
rect 20361 5525 20395 5559
rect 28825 5525 28859 5559
rect 31493 5525 31527 5559
rect 34913 5525 34947 5559
rect 35541 5525 35575 5559
rect 36921 5525 36955 5559
rect 37565 5525 37599 5559
rect 4997 5321 5031 5355
rect 5457 5321 5491 5355
rect 7849 5321 7883 5355
rect 9873 5321 9907 5355
rect 10885 5321 10919 5355
rect 12817 5321 12851 5355
rect 17417 5321 17451 5355
rect 18521 5321 18555 5355
rect 20729 5321 20763 5355
rect 24685 5321 24719 5355
rect 25145 5321 25179 5355
rect 30389 5321 30423 5355
rect 32781 5321 32815 5355
rect 34805 5321 34839 5355
rect 2237 5253 2271 5287
rect 3884 5253 3918 5287
rect 6377 5253 6411 5287
rect 10609 5253 10643 5287
rect 15209 5253 15243 5287
rect 17049 5253 17083 5287
rect 17233 5253 17267 5287
rect 18153 5253 18187 5287
rect 19616 5253 19650 5287
rect 23572 5253 23606 5287
rect 28825 5253 28859 5287
rect 29025 5253 29059 5287
rect 30757 5253 30791 5287
rect 34437 5253 34471 5287
rect 34653 5253 34687 5287
rect 1869 5185 1903 5219
rect 2513 5185 2547 5219
rect 3157 5185 3191 5219
rect 3617 5185 3651 5219
rect 5649 5185 5683 5219
rect 6561 5185 6595 5219
rect 7389 5185 7423 5219
rect 7665 5185 7699 5219
rect 8861 5185 8895 5219
rect 9597 5185 9631 5219
rect 9689 5185 9723 5219
rect 10333 5185 10367 5219
rect 10517 5185 10551 5219
rect 10725 5185 10759 5219
rect 11713 5185 11747 5219
rect 13001 5185 13035 5219
rect 13461 5185 13495 5219
rect 13645 5185 13679 5219
rect 15025 5185 15059 5219
rect 15853 5185 15887 5219
rect 18337 5185 18371 5219
rect 19349 5185 19383 5219
rect 21833 5185 21867 5219
rect 22569 5185 22603 5219
rect 25329 5185 25363 5219
rect 25421 5185 25455 5219
rect 25697 5185 25731 5219
rect 26341 5185 26375 5219
rect 27169 5185 27203 5219
rect 27813 5185 27847 5219
rect 29837 5185 29871 5219
rect 30573 5185 30607 5219
rect 30849 5185 30883 5219
rect 31493 5185 31527 5219
rect 32689 5185 32723 5219
rect 33517 5185 33551 5219
rect 35449 5185 35483 5219
rect 36093 5185 36127 5219
rect 36737 5185 36771 5219
rect 37841 5185 37875 5219
rect 7481 5117 7515 5151
rect 11529 5117 11563 5151
rect 14841 5117 14875 5151
rect 15669 5117 15703 5151
rect 23305 5117 23339 5151
rect 25605 5117 25639 5151
rect 1685 5049 1719 5083
rect 26985 5049 27019 5083
rect 29193 5049 29227 5083
rect 35265 5049 35299 5083
rect 2329 4981 2363 5015
rect 2973 4981 3007 5015
rect 6745 4981 6779 5015
rect 7665 4981 7699 5015
rect 8677 4981 8711 5015
rect 11897 4981 11931 5015
rect 13829 4981 13863 5015
rect 16037 4981 16071 5015
rect 22017 4981 22051 5015
rect 22753 4981 22787 5015
rect 26157 4981 26191 5015
rect 27629 4981 27663 5015
rect 29009 4981 29043 5015
rect 29653 4981 29687 5015
rect 31309 4981 31343 5015
rect 33333 4981 33367 5015
rect 34621 4981 34655 5015
rect 35909 4981 35943 5015
rect 36553 4981 36587 5015
rect 38025 4981 38059 5015
rect 4353 4777 4387 4811
rect 7665 4777 7699 4811
rect 8125 4777 8159 4811
rect 11805 4777 11839 4811
rect 14657 4777 14691 4811
rect 18613 4777 18647 4811
rect 22017 4777 22051 4811
rect 29745 4777 29779 4811
rect 31401 4777 31435 4811
rect 31585 4777 31619 4811
rect 32229 4777 32263 4811
rect 33057 4777 33091 4811
rect 33241 4777 33275 4811
rect 34897 4777 34931 4811
rect 35081 4777 35115 4811
rect 2421 4709 2455 4743
rect 3065 4709 3099 4743
rect 5273 4709 5307 4743
rect 7205 4709 7239 4743
rect 9781 4709 9815 4743
rect 23397 4709 23431 4743
rect 25329 4709 25363 4743
rect 29929 4709 29963 4743
rect 32413 4709 32447 4743
rect 8953 4641 8987 4675
rect 10425 4641 10459 4675
rect 15117 4641 15151 4675
rect 17233 4641 17267 4675
rect 18245 4641 18279 4675
rect 19533 4641 19567 4675
rect 19901 4641 19935 4675
rect 1961 4573 1995 4607
rect 2605 4573 2639 4607
rect 3249 4573 3283 4607
rect 3985 4573 4019 4607
rect 4813 4573 4847 4607
rect 4997 4573 5031 4607
rect 5089 4573 5123 4607
rect 5365 4573 5399 4607
rect 5825 4573 5859 4607
rect 6081 4573 6115 4607
rect 7849 4573 7883 4607
rect 7941 4573 7975 4607
rect 8217 4573 8251 4607
rect 9137 4573 9171 4607
rect 9321 4573 9355 4607
rect 9965 4573 9999 4607
rect 12449 4573 12483 4607
rect 12909 4573 12943 4607
rect 13093 4573 13127 4607
rect 14105 4573 14139 4607
rect 14381 4573 14415 4607
rect 14473 4573 14507 4607
rect 16957 4573 16991 4607
rect 18429 4573 18463 4607
rect 19717 4573 19751 4607
rect 20361 4573 20395 4607
rect 21649 4573 21683 4607
rect 21833 4573 21867 4607
rect 22477 4573 22511 4607
rect 23213 4573 23247 4607
rect 24409 4573 24443 4607
rect 25145 4573 25179 4607
rect 26249 4573 26283 4607
rect 26433 4573 26467 4607
rect 27813 4573 27847 4607
rect 28089 4573 28123 4607
rect 28733 4573 28767 4607
rect 29009 4573 29043 4607
rect 30573 4573 30607 4607
rect 33885 4573 33919 4607
rect 35725 4573 35759 4607
rect 36369 4573 36403 4607
rect 37013 4573 37047 4607
rect 37841 4573 37875 4607
rect 4169 4505 4203 4539
rect 10692 4505 10726 4539
rect 14289 4505 14323 4539
rect 15362 4505 15396 4539
rect 26617 4505 26651 4539
rect 29561 4505 29595 4539
rect 31217 4505 31251 4539
rect 31433 4505 31467 4539
rect 32045 4505 32079 4539
rect 32873 4505 32907 4539
rect 34713 4505 34747 4539
rect 1777 4437 1811 4471
rect 12265 4437 12299 4471
rect 13277 4437 13311 4471
rect 16497 4437 16531 4471
rect 20545 4437 20579 4471
rect 22661 4437 22695 4471
rect 24593 4437 24627 4471
rect 27629 4437 27663 4471
rect 27997 4437 28031 4471
rect 28549 4437 28583 4471
rect 28917 4437 28951 4471
rect 29761 4437 29795 4471
rect 30389 4437 30423 4471
rect 32245 4437 32279 4471
rect 33073 4437 33107 4471
rect 33701 4437 33735 4471
rect 34913 4437 34947 4471
rect 35541 4437 35575 4471
rect 36185 4437 36219 4471
rect 36829 4437 36863 4471
rect 38025 4437 38059 4471
rect 1961 4233 1995 4267
rect 3249 4233 3283 4267
rect 15025 4233 15059 4267
rect 16037 4233 16071 4267
rect 19809 4233 19843 4267
rect 23857 4233 23891 4267
rect 33517 4233 33551 4267
rect 35817 4233 35851 4267
rect 12050 4165 12084 4199
rect 15669 4165 15703 4199
rect 19441 4165 19475 4199
rect 36277 4165 36311 4199
rect 36477 4165 36511 4199
rect 2145 4097 2179 4131
rect 2789 4097 2823 4131
rect 3433 4097 3467 4131
rect 3893 4097 3927 4131
rect 4160 4097 4194 4131
rect 6561 4097 6595 4131
rect 6653 4097 6687 4131
rect 6929 4097 6963 4131
rect 7389 4097 7423 4131
rect 7656 4097 7690 4131
rect 9229 4097 9263 4131
rect 9496 4097 9530 4131
rect 11805 4097 11839 4131
rect 13645 4097 13679 4131
rect 13912 4097 13946 4131
rect 15485 4097 15519 4131
rect 15761 4097 15795 4131
rect 15853 4097 15887 4131
rect 17305 4097 17339 4131
rect 19257 4097 19291 4131
rect 19533 4097 19567 4131
rect 19625 4097 19659 4131
rect 20453 4097 20487 4131
rect 21281 4097 21315 4131
rect 21833 4097 21867 4131
rect 22100 4097 22134 4131
rect 23673 4097 23707 4131
rect 24685 4097 24719 4131
rect 24869 4097 24903 4131
rect 25513 4097 25547 4131
rect 26065 4097 26099 4131
rect 26157 4097 26191 4131
rect 26341 4097 26375 4131
rect 27252 4097 27286 4131
rect 28825 4097 28859 4131
rect 30297 4097 30331 4131
rect 30481 4097 30515 4131
rect 30573 4097 30607 4131
rect 31217 4097 31251 4131
rect 31401 4097 31435 4131
rect 31493 4097 31527 4131
rect 32404 4097 32438 4131
rect 34704 4097 34738 4131
rect 37841 4097 37875 4131
rect 17049 4029 17083 4063
rect 20269 4029 20303 4063
rect 24501 4029 24535 4063
rect 26985 4029 27019 4063
rect 29101 4029 29135 4063
rect 32137 4029 32171 4063
rect 34437 4029 34471 4063
rect 6377 3961 6411 3995
rect 6837 3961 6871 3995
rect 10609 3961 10643 3995
rect 20637 3961 20671 3995
rect 25329 3961 25363 3995
rect 36645 3961 36679 3995
rect 2605 3893 2639 3927
rect 5273 3893 5307 3927
rect 8769 3893 8803 3927
rect 13185 3893 13219 3927
rect 18429 3893 18463 3927
rect 21097 3893 21131 3927
rect 23213 3893 23247 3927
rect 28365 3893 28399 3927
rect 30113 3893 30147 3927
rect 31033 3893 31067 3927
rect 36461 3893 36495 3927
rect 38025 3893 38059 3927
rect 2421 3689 2455 3723
rect 3801 3689 3835 3723
rect 7113 3689 7147 3723
rect 8217 3689 8251 3723
rect 10977 3689 11011 3723
rect 11989 3689 12023 3723
rect 13553 3689 13587 3723
rect 16221 3689 16255 3723
rect 18705 3689 18739 3723
rect 25973 3689 26007 3723
rect 31125 3689 31159 3723
rect 31769 3689 31803 3723
rect 31953 3689 31987 3723
rect 32597 3689 32631 3723
rect 33425 3689 33459 3723
rect 33609 3689 33643 3723
rect 36737 3689 36771 3723
rect 36921 3689 36955 3723
rect 6653 3621 6687 3655
rect 25881 3621 25915 3655
rect 32781 3621 32815 3655
rect 7573 3553 7607 3587
rect 14841 3553 14875 3587
rect 17325 3553 17359 3587
rect 19257 3553 19291 3587
rect 21649 3553 21683 3587
rect 22477 3553 22511 3587
rect 24409 3553 24443 3587
rect 25513 3553 25547 3587
rect 27169 3553 27203 3587
rect 34713 3553 34747 3587
rect 1961 3485 1995 3519
rect 2605 3485 2639 3519
rect 3249 3485 3283 3519
rect 3985 3485 4019 3519
rect 4445 3485 4479 3519
rect 5273 3485 5307 3519
rect 7297 3485 7331 3519
rect 7389 3485 7423 3519
rect 7665 3485 7699 3519
rect 8401 3485 8435 3519
rect 9137 3485 9171 3519
rect 9413 3485 9447 3519
rect 10425 3485 10459 3519
rect 10701 3485 10735 3519
rect 10793 3485 10827 3519
rect 11457 3485 11491 3519
rect 11713 3485 11747 3519
rect 11805 3485 11839 3519
rect 13001 3485 13035 3519
rect 13277 3485 13311 3519
rect 13369 3485 13403 3519
rect 14381 3485 14415 3519
rect 16865 3485 16899 3519
rect 19441 3485 19475 3519
rect 20545 3485 20579 3519
rect 20913 3485 20947 3519
rect 21833 3485 21867 3519
rect 24593 3485 24627 3519
rect 24777 3485 24811 3519
rect 26433 3485 26467 3519
rect 29745 3485 29779 3519
rect 34980 3485 35014 3519
rect 37657 3485 37691 3519
rect 4629 3417 4663 3451
rect 5540 3417 5574 3451
rect 10609 3417 10643 3451
rect 11621 3417 11655 3451
rect 13185 3417 13219 3451
rect 15086 3417 15120 3451
rect 17570 3417 17604 3451
rect 19625 3417 19659 3451
rect 20729 3417 20763 3451
rect 20821 3417 20855 3451
rect 22744 3417 22778 3451
rect 27436 3417 27470 3451
rect 30012 3417 30046 3451
rect 31585 3417 31619 3451
rect 32413 3417 32447 3451
rect 33241 3417 33275 3451
rect 36553 3417 36587 3451
rect 1777 3349 1811 3383
rect 3065 3349 3099 3383
rect 4813 3349 4847 3383
rect 14197 3349 14231 3383
rect 16681 3349 16715 3383
rect 21097 3349 21131 3383
rect 22017 3349 22051 3383
rect 23857 3349 23891 3383
rect 26617 3349 26651 3383
rect 28549 3349 28583 3383
rect 31795 3349 31829 3383
rect 32623 3349 32657 3383
rect 33451 3349 33485 3383
rect 36093 3349 36127 3383
rect 36753 3349 36787 3383
rect 37841 3349 37875 3383
rect 1777 3145 1811 3179
rect 4353 3145 4387 3179
rect 5641 3145 5675 3179
rect 8033 3145 8067 3179
rect 15945 3145 15979 3179
rect 18521 3145 18555 3179
rect 19901 3145 19935 3179
rect 20729 3145 20763 3179
rect 24501 3145 24535 3179
rect 25789 3145 25823 3179
rect 27813 3145 27847 3179
rect 28667 3145 28701 3179
rect 29485 3145 29519 3179
rect 29653 3145 29687 3179
rect 31493 3145 31527 3179
rect 33993 3145 34027 3179
rect 34161 3145 34195 3179
rect 35557 3145 35591 3179
rect 35725 3145 35759 3179
rect 36553 3145 36587 3179
rect 10425 3077 10459 3111
rect 18245 3077 18279 3111
rect 22017 3077 22051 3111
rect 22109 3077 22143 3111
rect 27353 3077 27387 3111
rect 28457 3077 28491 3111
rect 29285 3077 29319 3111
rect 30380 3077 30414 3111
rect 33793 3077 33827 3111
rect 35357 3077 35391 3111
rect 36185 3077 36219 3111
rect 36385 3077 36419 3111
rect 1961 3009 1995 3043
rect 2605 3009 2639 3043
rect 3249 3009 3283 3043
rect 3893 3009 3927 3043
rect 4537 3009 4571 3043
rect 5181 3009 5215 3043
rect 5825 3009 5859 3043
rect 6653 3009 6687 3043
rect 6920 3009 6954 3043
rect 10149 3009 10183 3043
rect 10333 3009 10367 3043
rect 10517 3009 10551 3043
rect 11529 3009 11563 3043
rect 11796 3009 11830 3043
rect 13369 3009 13403 3043
rect 13553 3009 13587 3043
rect 13645 3009 13679 3043
rect 13737 3009 13771 3043
rect 16129 3009 16163 3043
rect 17969 3009 18003 3043
rect 18153 3009 18187 3043
rect 18337 3009 18371 3043
rect 19625 3009 19659 3043
rect 19717 3009 19751 3043
rect 20361 3009 20395 3043
rect 20545 3009 20579 3043
rect 21833 3009 21867 3043
rect 22201 3009 22235 3043
rect 23029 3009 23063 3043
rect 24317 3009 24351 3043
rect 26433 3009 26467 3043
rect 30113 3009 30147 3043
rect 32137 3009 32171 3043
rect 32873 3009 32907 3043
rect 34621 3009 34655 3043
rect 37289 3009 37323 3043
rect 8861 2941 8895 2975
rect 9137 2941 9171 2975
rect 14657 2941 14691 2975
rect 14933 2941 14967 2975
rect 16681 2941 16715 2975
rect 16957 2941 16991 2975
rect 22845 2941 22879 2975
rect 24133 2941 24167 2975
rect 25329 2941 25363 2975
rect 3065 2873 3099 2907
rect 22385 2873 22419 2907
rect 25697 2873 25731 2907
rect 27721 2873 27755 2907
rect 33057 2873 33091 2907
rect 34805 2873 34839 2907
rect 2421 2805 2455 2839
rect 3709 2805 3743 2839
rect 4997 2805 5031 2839
rect 10701 2805 10735 2839
rect 12909 2805 12943 2839
rect 13921 2805 13955 2839
rect 23213 2805 23247 2839
rect 26249 2805 26283 2839
rect 28641 2805 28675 2839
rect 28825 2805 28859 2839
rect 29469 2805 29503 2839
rect 32321 2805 32355 2839
rect 33977 2805 34011 2839
rect 35541 2805 35575 2839
rect 36369 2805 36403 2839
rect 37473 2805 37507 2839
rect 6745 2601 6779 2635
rect 7389 2601 7423 2635
rect 10333 2601 10367 2635
rect 10793 2601 10827 2635
rect 11897 2601 11931 2635
rect 15945 2601 15979 2635
rect 19441 2601 19475 2635
rect 21281 2601 21315 2635
rect 22753 2601 22787 2635
rect 26249 2601 26283 2635
rect 27721 2601 27755 2635
rect 28549 2601 28583 2635
rect 31217 2601 31251 2635
rect 17325 2533 17359 2567
rect 20177 2533 20211 2567
rect 23765 2533 23799 2567
rect 27169 2533 27203 2567
rect 30481 2533 30515 2567
rect 33793 2533 33827 2567
rect 35633 2533 35667 2567
rect 37473 2533 37507 2567
rect 3249 2465 3283 2499
rect 8401 2465 8435 2499
rect 9965 2465 9999 2499
rect 12633 2465 12667 2499
rect 14105 2465 14139 2499
rect 14381 2465 14415 2499
rect 20913 2465 20947 2499
rect 22385 2465 22419 2499
rect 25789 2465 25823 2499
rect 1409 2397 1443 2431
rect 2605 2397 2639 2431
rect 3801 2397 3835 2431
rect 4721 2397 4755 2431
rect 4997 2397 5031 2431
rect 6929 2397 6963 2431
rect 7573 2397 7607 2431
rect 8125 2397 8159 2431
rect 8217 2397 8251 2431
rect 8953 2397 8987 2431
rect 9321 2397 9355 2431
rect 10149 2397 10183 2431
rect 10977 2397 11011 2431
rect 12081 2397 12115 2431
rect 12817 2397 12851 2431
rect 15393 2397 15427 2431
rect 15577 2397 15611 2431
rect 15761 2397 15795 2431
rect 16773 2397 16807 2431
rect 16957 2397 16991 2431
rect 17187 2397 17221 2431
rect 17877 2397 17911 2431
rect 17969 2397 18003 2431
rect 19257 2397 19291 2431
rect 19993 2397 20027 2431
rect 21097 2397 21131 2431
rect 22569 2397 22603 2431
rect 23581 2397 23615 2431
rect 24409 2397 24443 2431
rect 25513 2397 25547 2431
rect 25605 2397 25639 2431
rect 26433 2397 26467 2431
rect 26985 2397 27019 2431
rect 27905 2397 27939 2431
rect 29561 2397 29595 2431
rect 30297 2397 30331 2431
rect 31033 2397 31067 2431
rect 32137 2397 32171 2431
rect 32873 2397 32907 2431
rect 33609 2397 33643 2431
rect 34713 2397 34747 2431
rect 35449 2397 35483 2431
rect 36185 2397 36219 2431
rect 37289 2397 37323 2431
rect 9137 2329 9171 2363
rect 9229 2329 9263 2363
rect 13001 2329 13035 2363
rect 15669 2329 15703 2363
rect 17049 2329 17083 2363
rect 28365 2329 28399 2363
rect 28581 2329 28615 2363
rect 1593 2261 1627 2295
rect 2421 2261 2455 2295
rect 3985 2261 4019 2295
rect 9505 2261 9539 2295
rect 18153 2261 18187 2295
rect 24593 2261 24627 2295
rect 28733 2261 28767 2295
rect 29745 2261 29779 2295
rect 32321 2261 32355 2295
rect 33057 2261 33091 2295
rect 34897 2261 34931 2295
rect 36369 2261 36403 2295
<< metal1 >>
rect 1104 47354 38824 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 38824 47354
rect 1104 47280 38824 47302
rect 12250 47240 12256 47252
rect 12211 47212 12256 47240
rect 12250 47200 12256 47212
rect 12308 47200 12314 47252
rect 20254 47240 20260 47252
rect 20215 47212 20260 47240
rect 20254 47200 20260 47212
rect 20312 47200 20318 47252
rect 28258 47240 28264 47252
rect 28219 47212 28264 47240
rect 28258 47200 28264 47212
rect 28316 47200 28322 47252
rect 4154 46996 4160 47048
rect 4212 47036 4218 47048
rect 4249 47039 4307 47045
rect 4249 47036 4261 47039
rect 4212 47008 4261 47036
rect 4212 46996 4218 47008
rect 4249 47005 4261 47008
rect 4295 47005 4307 47039
rect 4249 46999 4307 47005
rect 12069 47039 12127 47045
rect 12069 47005 12081 47039
rect 12115 47036 12127 47039
rect 12434 47036 12440 47048
rect 12115 47008 12440 47036
rect 12115 47005 12127 47008
rect 12069 46999 12127 47005
rect 12434 46996 12440 47008
rect 12492 46996 12498 47048
rect 20073 47039 20131 47045
rect 20073 47005 20085 47039
rect 20119 47036 20131 47039
rect 20346 47036 20352 47048
rect 20119 47008 20352 47036
rect 20119 47005 20131 47008
rect 20073 46999 20131 47005
rect 20346 46996 20352 47008
rect 20404 46996 20410 47048
rect 28074 47036 28080 47048
rect 28035 47008 28080 47036
rect 28074 46996 28080 47008
rect 28132 46996 28138 47048
rect 36170 47036 36176 47048
rect 36131 47008 36176 47036
rect 36170 46996 36176 47008
rect 36228 46996 36234 47048
rect 4614 46968 4620 46980
rect 4575 46940 4620 46968
rect 4614 46928 4620 46940
rect 4672 46928 4678 46980
rect 36262 46900 36268 46912
rect 36223 46872 36268 46900
rect 36262 46860 36268 46872
rect 36320 46860 36326 46912
rect 1104 46810 38824 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 38824 46810
rect 1104 46736 38824 46758
rect 12434 46696 12440 46708
rect 12395 46668 12440 46696
rect 12434 46656 12440 46668
rect 12492 46656 12498 46708
rect 12618 46560 12624 46572
rect 12579 46532 12624 46560
rect 12618 46520 12624 46532
rect 12676 46520 12682 46572
rect 15378 46520 15384 46572
rect 15436 46560 15442 46572
rect 16117 46563 16175 46569
rect 16117 46560 16129 46563
rect 15436 46532 16129 46560
rect 15436 46520 15442 46532
rect 16117 46529 16129 46532
rect 16163 46529 16175 46563
rect 16117 46523 16175 46529
rect 15933 46359 15991 46365
rect 15933 46325 15945 46359
rect 15979 46356 15991 46359
rect 28074 46356 28080 46368
rect 15979 46328 28080 46356
rect 15979 46325 15991 46328
rect 15933 46319 15991 46325
rect 28074 46316 28080 46328
rect 28132 46316 28138 46368
rect 1104 46266 38824 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 38824 46266
rect 1104 46192 38824 46214
rect 1104 45722 38824 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 38824 45722
rect 1104 45648 38824 45670
rect 1104 45178 38824 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 38824 45178
rect 1104 45104 38824 45126
rect 1104 44634 38824 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 38824 44634
rect 1104 44560 38824 44582
rect 1104 44090 38824 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 38824 44090
rect 1104 44016 38824 44038
rect 1104 43546 38824 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 38824 43546
rect 1104 43472 38824 43494
rect 1104 43002 38824 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 38824 43002
rect 1104 42928 38824 42950
rect 1104 42458 38824 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 38824 42458
rect 1104 42384 38824 42406
rect 1104 41914 38824 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 38824 41914
rect 1104 41840 38824 41862
rect 1104 41370 38824 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 38824 41370
rect 1104 41296 38824 41318
rect 1104 40826 38824 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 38824 40826
rect 1104 40752 38824 40774
rect 1104 40282 38824 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 38824 40282
rect 1104 40208 38824 40230
rect 1104 39738 38824 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 38824 39738
rect 1104 39664 38824 39686
rect 1104 39194 38824 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 38824 39194
rect 1104 39120 38824 39142
rect 1104 38650 38824 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 38824 38650
rect 1104 38576 38824 38598
rect 1104 38106 38824 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 38824 38106
rect 1104 38032 38824 38054
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 22002 34592 22008 34604
rect 21963 34564 22008 34592
rect 22002 34552 22008 34564
rect 22060 34552 22066 34604
rect 21818 34388 21824 34400
rect 21779 34360 21824 34388
rect 21818 34348 21824 34360
rect 21876 34348 21882 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 17954 33940 17960 33992
rect 18012 33980 18018 33992
rect 19429 33983 19487 33989
rect 19429 33980 19441 33983
rect 18012 33952 19441 33980
rect 18012 33940 18018 33952
rect 19429 33949 19441 33952
rect 19475 33949 19487 33983
rect 19429 33943 19487 33949
rect 20533 33983 20591 33989
rect 20533 33949 20545 33983
rect 20579 33980 20591 33983
rect 21174 33980 21180 33992
rect 20579 33952 21180 33980
rect 20579 33949 20591 33952
rect 20533 33943 20591 33949
rect 21174 33940 21180 33952
rect 21232 33940 21238 33992
rect 22462 33980 22468 33992
rect 22423 33952 22468 33980
rect 22462 33940 22468 33952
rect 22520 33940 22526 33992
rect 22646 33980 22652 33992
rect 22607 33952 22652 33980
rect 22646 33940 22652 33952
rect 22704 33940 22710 33992
rect 22833 33983 22891 33989
rect 22833 33949 22845 33983
rect 22879 33980 22891 33983
rect 23477 33983 23535 33989
rect 23477 33980 23489 33983
rect 22879 33952 23489 33980
rect 22879 33949 22891 33952
rect 22833 33943 22891 33949
rect 23477 33949 23489 33952
rect 23523 33949 23535 33983
rect 23477 33943 23535 33949
rect 20254 33872 20260 33924
rect 20312 33912 20318 33924
rect 20778 33915 20836 33921
rect 20778 33912 20790 33915
rect 20312 33884 20790 33912
rect 20312 33872 20318 33884
rect 20778 33881 20790 33884
rect 20824 33881 20836 33915
rect 20778 33875 20836 33881
rect 19245 33847 19303 33853
rect 19245 33813 19257 33847
rect 19291 33844 19303 33847
rect 19426 33844 19432 33856
rect 19291 33816 19432 33844
rect 19291 33813 19303 33816
rect 19245 33807 19303 33813
rect 19426 33804 19432 33816
rect 19484 33804 19490 33856
rect 21910 33844 21916 33856
rect 21871 33816 21916 33844
rect 21910 33804 21916 33816
rect 21968 33804 21974 33856
rect 23290 33844 23296 33856
rect 23251 33816 23296 33844
rect 23290 33804 23296 33816
rect 23348 33804 23354 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 17681 33643 17739 33649
rect 17681 33609 17693 33643
rect 17727 33609 17739 33643
rect 20254 33640 20260 33652
rect 20215 33612 20260 33640
rect 17681 33603 17739 33609
rect 17696 33572 17724 33603
rect 20254 33600 20260 33612
rect 20312 33600 20318 33652
rect 21269 33643 21327 33649
rect 21269 33609 21281 33643
rect 21315 33640 21327 33643
rect 22002 33640 22008 33652
rect 21315 33612 22008 33640
rect 21315 33609 21327 33612
rect 21269 33603 21327 33609
rect 22002 33600 22008 33612
rect 22060 33600 22066 33652
rect 18570 33575 18628 33581
rect 18570 33572 18582 33575
rect 17696 33544 18582 33572
rect 18570 33541 18582 33544
rect 18616 33541 18628 33575
rect 22462 33572 22468 33584
rect 18570 33535 18628 33541
rect 20916 33544 22468 33572
rect 17865 33507 17923 33513
rect 17865 33473 17877 33507
rect 17911 33504 17923 33507
rect 18414 33504 18420 33516
rect 17911 33476 18420 33504
rect 17911 33473 17923 33476
rect 17865 33467 17923 33473
rect 18414 33464 18420 33476
rect 18472 33464 18478 33516
rect 20441 33507 20499 33513
rect 20441 33473 20453 33507
rect 20487 33504 20499 33507
rect 20806 33504 20812 33516
rect 20487 33476 20812 33504
rect 20487 33473 20499 33476
rect 20441 33467 20499 33473
rect 20806 33464 20812 33476
rect 20864 33464 20870 33516
rect 20916 33513 20944 33544
rect 22462 33532 22468 33544
rect 22520 33532 22526 33584
rect 22640 33575 22698 33581
rect 22640 33541 22652 33575
rect 22686 33572 22698 33575
rect 23290 33572 23296 33584
rect 22686 33544 23296 33572
rect 22686 33541 22698 33544
rect 22640 33535 22698 33541
rect 23290 33532 23296 33544
rect 23348 33532 23354 33584
rect 20901 33507 20959 33513
rect 20901 33473 20913 33507
rect 20947 33473 20959 33507
rect 21082 33504 21088 33516
rect 21043 33476 21088 33504
rect 20901 33467 20959 33473
rect 21082 33464 21088 33476
rect 21140 33464 21146 33516
rect 24394 33504 24400 33516
rect 24355 33476 24400 33504
rect 24394 33464 24400 33476
rect 24452 33464 24458 33516
rect 16942 33396 16948 33448
rect 17000 33436 17006 33448
rect 18325 33439 18383 33445
rect 18325 33436 18337 33439
rect 17000 33408 18337 33436
rect 17000 33396 17006 33408
rect 18325 33405 18337 33408
rect 18371 33405 18383 33439
rect 18325 33399 18383 33405
rect 21174 33396 21180 33448
rect 21232 33436 21238 33448
rect 22373 33439 22431 33445
rect 22373 33436 22385 33439
rect 21232 33408 22385 33436
rect 21232 33396 21238 33408
rect 22373 33405 22385 33408
rect 22419 33405 22431 33439
rect 22373 33399 22431 33405
rect 19705 33303 19763 33309
rect 19705 33269 19717 33303
rect 19751 33300 19763 33303
rect 19978 33300 19984 33312
rect 19751 33272 19984 33300
rect 19751 33269 19763 33272
rect 19705 33263 19763 33269
rect 19978 33260 19984 33272
rect 20036 33260 20042 33312
rect 22370 33260 22376 33312
rect 22428 33300 22434 33312
rect 23753 33303 23811 33309
rect 23753 33300 23765 33303
rect 22428 33272 23765 33300
rect 22428 33260 22434 33272
rect 23753 33269 23765 33272
rect 23799 33269 23811 33303
rect 24210 33300 24216 33312
rect 24171 33272 24216 33300
rect 23753 33263 23811 33269
rect 24210 33260 24216 33272
rect 24268 33260 24274 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 17865 33099 17923 33105
rect 17865 33065 17877 33099
rect 17911 33096 17923 33099
rect 17954 33096 17960 33108
rect 17911 33068 17960 33096
rect 17911 33065 17923 33068
rect 17865 33059 17923 33065
rect 17954 33056 17960 33068
rect 18012 33056 18018 33108
rect 18414 33056 18420 33108
rect 18472 33096 18478 33108
rect 18693 33099 18751 33105
rect 18693 33096 18705 33099
rect 18472 33068 18705 33096
rect 18472 33056 18478 33068
rect 18693 33065 18705 33068
rect 18739 33065 18751 33099
rect 18693 33059 18751 33065
rect 20806 33056 20812 33108
rect 20864 33096 20870 33108
rect 23293 33099 23351 33105
rect 23293 33096 23305 33099
rect 20864 33068 23305 33096
rect 20864 33056 20870 33068
rect 23293 33065 23305 33068
rect 23339 33065 23351 33099
rect 23293 33059 23351 33065
rect 24394 33056 24400 33108
rect 24452 33096 24458 33108
rect 24765 33099 24823 33105
rect 24765 33096 24777 33099
rect 24452 33068 24777 33096
rect 24452 33056 24458 33068
rect 24765 33065 24777 33068
rect 24811 33065 24823 33099
rect 24765 33059 24823 33065
rect 17402 32920 17408 32972
rect 17460 32960 17466 32972
rect 17497 32963 17555 32969
rect 17497 32960 17509 32963
rect 17460 32932 17509 32960
rect 17460 32920 17466 32932
rect 17497 32929 17509 32932
rect 17543 32960 17555 32963
rect 18325 32963 18383 32969
rect 18325 32960 18337 32963
rect 17543 32932 18337 32960
rect 17543 32929 17555 32932
rect 17497 32923 17555 32929
rect 18325 32929 18337 32932
rect 18371 32929 18383 32963
rect 18325 32923 18383 32929
rect 22462 32920 22468 32972
rect 22520 32960 22526 32972
rect 22925 32963 22983 32969
rect 22925 32960 22937 32963
rect 22520 32932 22937 32960
rect 22520 32920 22526 32932
rect 22925 32929 22937 32932
rect 22971 32960 22983 32963
rect 24397 32963 24455 32969
rect 24397 32960 24409 32963
rect 22971 32932 24409 32960
rect 22971 32929 22983 32932
rect 22925 32923 22983 32929
rect 24397 32929 24409 32932
rect 24443 32960 24455 32963
rect 24762 32960 24768 32972
rect 24443 32932 24768 32960
rect 24443 32929 24455 32932
rect 24397 32923 24455 32929
rect 24762 32920 24768 32932
rect 24820 32920 24826 32972
rect 17034 32892 17040 32904
rect 16995 32864 17040 32892
rect 17034 32852 17040 32864
rect 17092 32852 17098 32904
rect 17678 32892 17684 32904
rect 17639 32864 17684 32892
rect 17678 32852 17684 32864
rect 17736 32852 17742 32904
rect 18506 32892 18512 32904
rect 18467 32864 18512 32892
rect 18506 32852 18512 32864
rect 18564 32852 18570 32904
rect 19245 32895 19303 32901
rect 19245 32861 19257 32895
rect 19291 32861 19303 32895
rect 19245 32855 19303 32861
rect 19512 32895 19570 32901
rect 19512 32861 19524 32895
rect 19558 32861 19570 32895
rect 19512 32855 19570 32861
rect 21085 32895 21143 32901
rect 21085 32861 21097 32895
rect 21131 32892 21143 32895
rect 21174 32892 21180 32904
rect 21131 32864 21180 32892
rect 21131 32861 21143 32864
rect 21085 32855 21143 32861
rect 16850 32756 16856 32768
rect 16811 32728 16856 32756
rect 16850 32716 16856 32728
rect 16908 32716 16914 32768
rect 19260 32756 19288 32855
rect 19426 32784 19432 32836
rect 19484 32824 19490 32836
rect 19536 32824 19564 32855
rect 21100 32824 21128 32855
rect 21174 32852 21180 32864
rect 21232 32852 21238 32904
rect 21352 32895 21410 32901
rect 21352 32861 21364 32895
rect 21398 32892 21410 32895
rect 21818 32892 21824 32904
rect 21398 32864 21824 32892
rect 21398 32861 21410 32864
rect 21352 32855 21410 32861
rect 21818 32852 21824 32864
rect 21876 32852 21882 32904
rect 23109 32895 23167 32901
rect 23109 32861 23121 32895
rect 23155 32861 23167 32895
rect 24578 32892 24584 32904
rect 24539 32864 24584 32892
rect 23109 32855 23167 32861
rect 19484 32796 19564 32824
rect 19628 32796 21128 32824
rect 19484 32784 19490 32796
rect 19628 32756 19656 32796
rect 21450 32784 21456 32836
rect 21508 32824 21514 32836
rect 23124 32824 23152 32855
rect 24578 32852 24584 32864
rect 24636 32852 24642 32904
rect 21508 32796 23152 32824
rect 21508 32784 21514 32796
rect 20622 32756 20628 32768
rect 19260 32728 19656 32756
rect 20583 32728 20628 32756
rect 20622 32716 20628 32728
rect 20680 32716 20686 32768
rect 20990 32716 20996 32768
rect 21048 32756 21054 32768
rect 22465 32759 22523 32765
rect 22465 32756 22477 32759
rect 21048 32728 22477 32756
rect 21048 32716 21054 32728
rect 22465 32725 22477 32728
rect 22511 32725 22523 32759
rect 22465 32719 22523 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 17678 32512 17684 32564
rect 17736 32552 17742 32564
rect 19705 32555 19763 32561
rect 19705 32552 19717 32555
rect 17736 32524 19717 32552
rect 17736 32512 17742 32524
rect 19705 32521 19717 32524
rect 19751 32521 19763 32555
rect 19705 32515 19763 32521
rect 21082 32512 21088 32564
rect 21140 32552 21146 32564
rect 21269 32555 21327 32561
rect 21269 32552 21281 32555
rect 21140 32524 21281 32552
rect 21140 32512 21146 32524
rect 21269 32521 21281 32524
rect 21315 32521 21327 32555
rect 22646 32552 22652 32564
rect 21269 32515 21327 32521
rect 22066 32524 22508 32552
rect 22607 32524 22652 32552
rect 16850 32444 16856 32496
rect 16908 32484 16914 32496
rect 17190 32487 17248 32493
rect 17190 32484 17202 32487
rect 16908 32456 17202 32484
rect 16908 32444 16914 32456
rect 17190 32453 17202 32456
rect 17236 32453 17248 32487
rect 17190 32447 17248 32453
rect 20530 32444 20536 32496
rect 20588 32484 20594 32496
rect 20901 32487 20959 32493
rect 20901 32484 20913 32487
rect 20588 32456 20913 32484
rect 20588 32444 20594 32456
rect 20901 32453 20913 32456
rect 20947 32453 20959 32487
rect 22066 32484 22094 32524
rect 22370 32484 22376 32496
rect 20901 32447 20959 32453
rect 21100 32456 22094 32484
rect 22331 32456 22376 32484
rect 16666 32376 16672 32428
rect 16724 32416 16730 32428
rect 16942 32416 16948 32428
rect 16724 32388 16948 32416
rect 16724 32376 16730 32388
rect 16942 32376 16948 32388
rect 17000 32376 17006 32428
rect 19153 32419 19211 32425
rect 19153 32385 19165 32419
rect 19199 32385 19211 32419
rect 19334 32416 19340 32428
rect 19295 32388 19340 32416
rect 19153 32379 19211 32385
rect 19168 32348 19196 32379
rect 19334 32376 19340 32388
rect 19392 32376 19398 32428
rect 19429 32419 19487 32425
rect 19429 32385 19441 32419
rect 19475 32385 19487 32419
rect 19429 32379 19487 32385
rect 19521 32419 19579 32425
rect 19521 32385 19533 32419
rect 19567 32416 19579 32419
rect 19610 32416 19616 32428
rect 19567 32388 19616 32416
rect 19567 32385 19579 32388
rect 19521 32379 19579 32385
rect 19242 32348 19248 32360
rect 19168 32320 19248 32348
rect 19242 32308 19248 32320
rect 19300 32308 19306 32360
rect 19444 32348 19472 32379
rect 19610 32376 19616 32388
rect 19668 32376 19674 32428
rect 20714 32416 20720 32428
rect 20675 32388 20720 32416
rect 20714 32376 20720 32388
rect 20772 32376 20778 32428
rect 20990 32416 20996 32428
rect 20951 32388 20996 32416
rect 20990 32376 20996 32388
rect 21048 32376 21054 32428
rect 21100 32425 21128 32456
rect 22370 32444 22376 32456
rect 22428 32444 22434 32496
rect 21085 32419 21143 32425
rect 21085 32385 21097 32419
rect 21131 32385 21143 32419
rect 21085 32379 21143 32385
rect 22002 32376 22008 32428
rect 22060 32416 22066 32428
rect 22097 32419 22155 32425
rect 22097 32416 22109 32419
rect 22060 32388 22109 32416
rect 22060 32376 22066 32388
rect 22097 32385 22109 32388
rect 22143 32385 22155 32419
rect 22278 32416 22284 32428
rect 22239 32388 22284 32416
rect 22097 32379 22155 32385
rect 22278 32376 22284 32388
rect 22336 32376 22342 32428
rect 22480 32425 22508 32524
rect 22646 32512 22652 32524
rect 22704 32512 22710 32564
rect 23652 32487 23710 32493
rect 23652 32453 23664 32487
rect 23698 32484 23710 32487
rect 24210 32484 24216 32496
rect 23698 32456 24216 32484
rect 23698 32453 23710 32456
rect 23652 32447 23710 32453
rect 24210 32444 24216 32456
rect 24268 32444 24274 32496
rect 22465 32419 22523 32425
rect 22465 32385 22477 32419
rect 22511 32416 22523 32419
rect 22554 32416 22560 32428
rect 22511 32388 22560 32416
rect 22511 32385 22523 32388
rect 22465 32379 22523 32385
rect 22554 32376 22560 32388
rect 22612 32376 22618 32428
rect 23385 32419 23443 32425
rect 23385 32385 23397 32419
rect 23431 32416 23443 32419
rect 23474 32416 23480 32428
rect 23431 32388 23480 32416
rect 23431 32385 23443 32388
rect 23385 32379 23443 32385
rect 23474 32376 23480 32388
rect 23532 32376 23538 32428
rect 25406 32416 25412 32428
rect 25367 32388 25412 32416
rect 25406 32376 25412 32388
rect 25464 32376 25470 32428
rect 20622 32348 20628 32360
rect 19444 32320 20628 32348
rect 20622 32308 20628 32320
rect 20680 32308 20686 32360
rect 18325 32215 18383 32221
rect 18325 32181 18337 32215
rect 18371 32212 18383 32215
rect 18414 32212 18420 32224
rect 18371 32184 18420 32212
rect 18371 32181 18383 32184
rect 18325 32175 18383 32181
rect 18414 32172 18420 32184
rect 18472 32212 18478 32224
rect 18874 32212 18880 32224
rect 18472 32184 18880 32212
rect 18472 32172 18478 32184
rect 18874 32172 18880 32184
rect 18932 32172 18938 32224
rect 23566 32172 23572 32224
rect 23624 32212 23630 32224
rect 24765 32215 24823 32221
rect 24765 32212 24777 32215
rect 23624 32184 24777 32212
rect 23624 32172 23630 32184
rect 24765 32181 24777 32184
rect 24811 32181 24823 32215
rect 25222 32212 25228 32224
rect 25183 32184 25228 32212
rect 24765 32175 24823 32181
rect 25222 32172 25228 32184
rect 25280 32172 25286 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 17034 31968 17040 32020
rect 17092 32008 17098 32020
rect 17681 32011 17739 32017
rect 17681 32008 17693 32011
rect 17092 31980 17693 32008
rect 17092 31968 17098 31980
rect 17681 31977 17693 31980
rect 17727 31977 17739 32011
rect 17681 31971 17739 31977
rect 18506 31968 18512 32020
rect 18564 32008 18570 32020
rect 19797 32011 19855 32017
rect 19797 32008 19809 32011
rect 18564 31980 19809 32008
rect 18564 31968 18570 31980
rect 19797 31977 19809 31980
rect 19843 31977 19855 32011
rect 21450 32008 21456 32020
rect 21411 31980 21456 32008
rect 19797 31971 19855 31977
rect 21450 31968 21456 31980
rect 21508 31968 21514 32020
rect 21913 32011 21971 32017
rect 21913 31977 21925 32011
rect 21959 32008 21971 32011
rect 22278 32008 22284 32020
rect 21959 31980 22284 32008
rect 21959 31977 21971 31980
rect 21913 31971 21971 31977
rect 22278 31968 22284 31980
rect 22336 31968 22342 32020
rect 23661 32011 23719 32017
rect 23661 31977 23673 32011
rect 23707 32008 23719 32011
rect 24578 32008 24584 32020
rect 23707 31980 24584 32008
rect 23707 31977 23719 31980
rect 23661 31971 23719 31977
rect 24578 31968 24584 31980
rect 24636 31968 24642 32020
rect 18693 31943 18751 31949
rect 18693 31909 18705 31943
rect 18739 31909 18751 31943
rect 18693 31903 18751 31909
rect 18708 31872 18736 31903
rect 23474 31900 23480 31952
rect 23532 31900 23538 31952
rect 17512 31844 18736 31872
rect 18892 31844 19656 31872
rect 17402 31804 17408 31816
rect 17363 31776 17408 31804
rect 17402 31764 17408 31776
rect 17460 31764 17466 31816
rect 17512 31813 17540 31844
rect 17497 31807 17555 31813
rect 17497 31773 17509 31807
rect 17543 31773 17555 31807
rect 17497 31767 17555 31773
rect 18141 31807 18199 31813
rect 18141 31773 18153 31807
rect 18187 31773 18199 31807
rect 18506 31804 18512 31816
rect 18419 31776 18512 31804
rect 18141 31767 18199 31773
rect 17954 31628 17960 31680
rect 18012 31668 18018 31680
rect 18156 31668 18184 31767
rect 18506 31764 18512 31776
rect 18564 31804 18570 31816
rect 18892 31804 18920 31844
rect 19628 31816 19656 31844
rect 20714 31832 20720 31884
rect 20772 31872 20778 31884
rect 22002 31872 22008 31884
rect 20772 31844 22008 31872
rect 20772 31832 20778 31844
rect 19242 31804 19248 31816
rect 18564 31776 18920 31804
rect 19203 31776 19248 31804
rect 18564 31764 18570 31776
rect 19242 31764 19248 31776
rect 19300 31764 19306 31816
rect 19426 31804 19432 31816
rect 19387 31776 19432 31804
rect 19426 31764 19432 31776
rect 19484 31764 19490 31816
rect 19610 31804 19616 31816
rect 19571 31776 19616 31804
rect 19610 31764 19616 31776
rect 19668 31764 19674 31816
rect 19978 31804 19984 31816
rect 19720 31776 19984 31804
rect 18322 31736 18328 31748
rect 18283 31708 18328 31736
rect 18322 31696 18328 31708
rect 18380 31696 18386 31748
rect 18414 31696 18420 31748
rect 18472 31736 18478 31748
rect 19521 31739 19579 31745
rect 18472 31708 18517 31736
rect 18472 31696 18478 31708
rect 19521 31705 19533 31739
rect 19567 31736 19579 31739
rect 19720 31736 19748 31776
rect 19978 31764 19984 31776
rect 20036 31804 20042 31816
rect 20438 31804 20444 31816
rect 20036 31776 20444 31804
rect 20036 31764 20042 31776
rect 20438 31764 20444 31776
rect 20496 31764 20502 31816
rect 20916 31813 20944 31844
rect 22002 31832 22008 31844
rect 22060 31832 22066 31884
rect 22462 31872 22468 31884
rect 22423 31844 22468 31872
rect 22462 31832 22468 31844
rect 22520 31832 22526 31884
rect 23382 31872 23388 31884
rect 23032 31844 23388 31872
rect 20901 31807 20959 31813
rect 20901 31773 20913 31807
rect 20947 31773 20959 31807
rect 20901 31767 20959 31773
rect 21177 31807 21235 31813
rect 21177 31773 21189 31807
rect 21223 31773 21235 31807
rect 21177 31767 21235 31773
rect 21269 31807 21327 31813
rect 21269 31773 21281 31807
rect 21315 31804 21327 31807
rect 22554 31804 22560 31816
rect 21315 31776 22560 31804
rect 21315 31773 21327 31776
rect 21269 31767 21327 31773
rect 21082 31736 21088 31748
rect 19567 31708 19748 31736
rect 21043 31708 21088 31736
rect 19567 31705 19579 31708
rect 19521 31699 19579 31705
rect 21082 31696 21088 31708
rect 21140 31696 21146 31748
rect 19242 31668 19248 31680
rect 18012 31640 19248 31668
rect 18012 31628 18018 31640
rect 19242 31628 19248 31640
rect 19300 31628 19306 31680
rect 21192 31668 21220 31767
rect 22554 31764 22560 31776
rect 22612 31804 22618 31816
rect 23032 31804 23060 31844
rect 23382 31832 23388 31844
rect 23440 31832 23446 31884
rect 23492 31872 23520 31900
rect 24394 31872 24400 31884
rect 23492 31844 24400 31872
rect 24394 31832 24400 31844
rect 24452 31832 24458 31884
rect 22612 31776 23060 31804
rect 23109 31807 23167 31813
rect 22612 31764 22618 31776
rect 23109 31773 23121 31807
rect 23155 31773 23167 31807
rect 23109 31767 23167 31773
rect 21542 31696 21548 31748
rect 21600 31736 21606 31748
rect 22002 31736 22008 31748
rect 21600 31708 22008 31736
rect 21600 31696 21606 31708
rect 22002 31696 22008 31708
rect 22060 31736 22066 31748
rect 23124 31736 23152 31767
rect 23198 31764 23204 31816
rect 23256 31804 23262 31816
rect 23293 31807 23351 31813
rect 23293 31804 23305 31807
rect 23256 31776 23305 31804
rect 23256 31764 23262 31776
rect 23293 31773 23305 31776
rect 23339 31773 23351 31807
rect 23400 31804 23428 31832
rect 23477 31807 23535 31813
rect 23477 31804 23489 31807
rect 23400 31776 23489 31804
rect 23293 31767 23351 31773
rect 23477 31773 23489 31776
rect 23523 31804 23535 31807
rect 24664 31807 24722 31813
rect 23523 31776 24624 31804
rect 23523 31773 23535 31776
rect 23477 31767 23535 31773
rect 24596 31748 24624 31776
rect 24664 31773 24676 31807
rect 24710 31804 24722 31807
rect 25222 31804 25228 31816
rect 24710 31776 25228 31804
rect 24710 31773 24722 31776
rect 24664 31767 24722 31773
rect 25222 31764 25228 31776
rect 25280 31764 25286 31816
rect 22060 31708 23152 31736
rect 22060 31696 22066 31708
rect 21818 31668 21824 31680
rect 21192 31640 21824 31668
rect 21818 31628 21824 31640
rect 21876 31628 21882 31680
rect 22278 31668 22284 31680
rect 22239 31640 22284 31668
rect 22278 31628 22284 31640
rect 22336 31628 22342 31680
rect 22370 31628 22376 31680
rect 22428 31668 22434 31680
rect 23124 31668 23152 31708
rect 23385 31739 23443 31745
rect 23385 31705 23397 31739
rect 23431 31736 23443 31739
rect 23566 31736 23572 31748
rect 23431 31708 23572 31736
rect 23431 31705 23443 31708
rect 23385 31699 23443 31705
rect 23566 31696 23572 31708
rect 23624 31696 23630 31748
rect 24578 31696 24584 31748
rect 24636 31696 24642 31748
rect 24210 31668 24216 31680
rect 22428 31640 22473 31668
rect 23124 31640 24216 31668
rect 22428 31628 22434 31640
rect 24210 31628 24216 31640
rect 24268 31628 24274 31680
rect 25038 31628 25044 31680
rect 25096 31668 25102 31680
rect 25777 31671 25835 31677
rect 25777 31668 25789 31671
rect 25096 31640 25789 31668
rect 25096 31628 25102 31640
rect 25777 31637 25789 31640
rect 25823 31637 25835 31671
rect 25777 31631 25835 31637
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 18322 31424 18328 31476
rect 18380 31464 18386 31476
rect 18969 31467 19027 31473
rect 18969 31464 18981 31467
rect 18380 31436 18981 31464
rect 18380 31424 18386 31436
rect 18969 31433 18981 31436
rect 19015 31433 19027 31467
rect 18969 31427 19027 31433
rect 19334 31424 19340 31476
rect 19392 31464 19398 31476
rect 20257 31467 20315 31473
rect 20257 31464 20269 31467
rect 19392 31436 20269 31464
rect 19392 31424 19398 31436
rect 20257 31433 20269 31436
rect 20303 31433 20315 31467
rect 20257 31427 20315 31433
rect 21082 31424 21088 31476
rect 21140 31464 21146 31476
rect 21821 31467 21879 31473
rect 21821 31464 21833 31467
rect 21140 31436 21833 31464
rect 21140 31424 21146 31436
rect 21821 31433 21833 31436
rect 21867 31433 21879 31467
rect 21821 31427 21879 31433
rect 23017 31467 23075 31473
rect 23017 31433 23029 31467
rect 23063 31464 23075 31467
rect 23063 31436 24440 31464
rect 23063 31433 23075 31436
rect 23017 31427 23075 31433
rect 18046 31356 18052 31408
rect 18104 31396 18110 31408
rect 18233 31399 18291 31405
rect 18233 31396 18245 31399
rect 18104 31368 18245 31396
rect 18104 31356 18110 31368
rect 18233 31365 18245 31368
rect 18279 31365 18291 31399
rect 18233 31359 18291 31365
rect 20717 31399 20775 31405
rect 20717 31365 20729 31399
rect 20763 31396 20775 31399
rect 22370 31396 22376 31408
rect 20763 31368 22376 31396
rect 20763 31365 20775 31368
rect 20717 31359 20775 31365
rect 16850 31328 16856 31340
rect 16811 31300 16856 31328
rect 16850 31288 16856 31300
rect 16908 31288 16914 31340
rect 17954 31328 17960 31340
rect 17915 31300 17960 31328
rect 17954 31288 17960 31300
rect 18012 31288 18018 31340
rect 18138 31328 18144 31340
rect 18099 31300 18144 31328
rect 18138 31288 18144 31300
rect 18196 31288 18202 31340
rect 18325 31331 18383 31337
rect 18325 31297 18337 31331
rect 18371 31328 18383 31331
rect 18506 31328 18512 31340
rect 18371 31300 18512 31328
rect 18371 31297 18383 31300
rect 18325 31291 18383 31297
rect 18506 31288 18512 31300
rect 18564 31328 18570 31340
rect 18782 31328 18788 31340
rect 18564 31300 18788 31328
rect 18564 31288 18570 31300
rect 18782 31288 18788 31300
rect 18840 31288 18846 31340
rect 18874 31288 18880 31340
rect 18932 31328 18938 31340
rect 19337 31331 19395 31337
rect 19337 31328 19349 31331
rect 18932 31300 19349 31328
rect 18932 31288 18938 31300
rect 19337 31297 19349 31300
rect 19383 31297 19395 31331
rect 19337 31291 19395 31297
rect 19429 31331 19487 31337
rect 19429 31297 19441 31331
rect 19475 31328 19487 31331
rect 20254 31328 20260 31340
rect 19475 31300 20260 31328
rect 19475 31297 19487 31300
rect 19429 31291 19487 31297
rect 20254 31288 20260 31300
rect 20312 31288 20318 31340
rect 20622 31328 20628 31340
rect 20583 31300 20628 31328
rect 20622 31288 20628 31300
rect 20680 31288 20686 31340
rect 21818 31288 21824 31340
rect 21876 31328 21882 31340
rect 22296 31337 22324 31368
rect 22370 31356 22376 31368
rect 22428 31356 22434 31408
rect 24412 31405 24440 31436
rect 25406 31424 25412 31476
rect 25464 31464 25470 31476
rect 25593 31467 25651 31473
rect 25593 31464 25605 31467
rect 25464 31436 25605 31464
rect 25464 31424 25470 31436
rect 25593 31433 25605 31436
rect 25639 31433 25651 31467
rect 25593 31427 25651 31433
rect 23385 31399 23443 31405
rect 23385 31365 23397 31399
rect 23431 31396 23443 31399
rect 24397 31399 24455 31405
rect 23431 31368 24348 31396
rect 23431 31365 23443 31368
rect 23385 31359 23443 31365
rect 22189 31331 22247 31337
rect 22189 31328 22201 31331
rect 21876 31300 22201 31328
rect 21876 31288 21882 31300
rect 22189 31297 22201 31300
rect 22235 31297 22247 31331
rect 22189 31291 22247 31297
rect 22281 31331 22339 31337
rect 22281 31297 22293 31331
rect 22327 31328 22339 31331
rect 24210 31328 24216 31340
rect 22327 31300 23336 31328
rect 24171 31300 24216 31328
rect 22327 31297 22339 31300
rect 22281 31291 22339 31297
rect 23308 31272 23336 31300
rect 24210 31288 24216 31300
rect 24268 31288 24274 31340
rect 24320 31328 24348 31368
rect 24397 31365 24409 31399
rect 24443 31365 24455 31399
rect 24397 31359 24455 31365
rect 24489 31399 24547 31405
rect 24489 31365 24501 31399
rect 24535 31396 24547 31399
rect 25038 31396 25044 31408
rect 24535 31368 25044 31396
rect 24535 31365 24547 31368
rect 24489 31359 24547 31365
rect 24504 31328 24532 31359
rect 25038 31356 25044 31368
rect 25096 31356 25102 31408
rect 24320 31300 24532 31328
rect 24578 31288 24584 31340
rect 24636 31328 24642 31340
rect 24636 31300 24681 31328
rect 24636 31288 24642 31300
rect 24762 31288 24768 31340
rect 24820 31288 24826 31340
rect 25409 31331 25467 31337
rect 25409 31297 25421 31331
rect 25455 31297 25467 31331
rect 26234 31328 26240 31340
rect 26195 31300 26240 31328
rect 25409 31291 25467 31297
rect 19613 31263 19671 31269
rect 19613 31229 19625 31263
rect 19659 31260 19671 31263
rect 20714 31260 20720 31272
rect 19659 31232 20720 31260
rect 19659 31229 19671 31232
rect 19613 31223 19671 31229
rect 20714 31220 20720 31232
rect 20772 31220 20778 31272
rect 20898 31260 20904 31272
rect 20859 31232 20904 31260
rect 20898 31220 20904 31232
rect 20956 31220 20962 31272
rect 22370 31220 22376 31272
rect 22428 31260 22434 31272
rect 22428 31232 22473 31260
rect 22428 31220 22434 31232
rect 23290 31220 23296 31272
rect 23348 31260 23354 31272
rect 23477 31263 23535 31269
rect 23477 31260 23489 31263
rect 23348 31232 23489 31260
rect 23348 31220 23354 31232
rect 23477 31229 23489 31232
rect 23523 31229 23535 31263
rect 23477 31223 23535 31229
rect 23569 31263 23627 31269
rect 23569 31229 23581 31263
rect 23615 31229 23627 31263
rect 23569 31223 23627 31229
rect 23014 31152 23020 31204
rect 23072 31192 23078 31204
rect 23584 31192 23612 31223
rect 24026 31220 24032 31272
rect 24084 31260 24090 31272
rect 24780 31260 24808 31288
rect 25225 31263 25283 31269
rect 25225 31260 25237 31263
rect 24084 31232 25237 31260
rect 24084 31220 24090 31232
rect 25225 31229 25237 31232
rect 25271 31229 25283 31263
rect 25225 31223 25283 31229
rect 23072 31164 23612 31192
rect 24765 31195 24823 31201
rect 23072 31152 23078 31164
rect 24765 31161 24777 31195
rect 24811 31192 24823 31195
rect 25424 31192 25452 31291
rect 26234 31288 26240 31300
rect 26292 31288 26298 31340
rect 24811 31164 25452 31192
rect 24811 31161 24823 31164
rect 24765 31155 24823 31161
rect 16574 31084 16580 31136
rect 16632 31124 16638 31136
rect 16669 31127 16727 31133
rect 16669 31124 16681 31127
rect 16632 31096 16681 31124
rect 16632 31084 16638 31096
rect 16669 31093 16681 31096
rect 16715 31093 16727 31127
rect 16669 31087 16727 31093
rect 16758 31084 16764 31136
rect 16816 31124 16822 31136
rect 18509 31127 18567 31133
rect 18509 31124 18521 31127
rect 16816 31096 18521 31124
rect 16816 31084 16822 31096
rect 18509 31093 18521 31096
rect 18555 31093 18567 31127
rect 26050 31124 26056 31136
rect 26011 31096 26056 31124
rect 18509 31087 18567 31093
rect 26050 31084 26056 31096
rect 26108 31084 26114 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 23290 30880 23296 30932
rect 23348 30920 23354 30932
rect 24397 30923 24455 30929
rect 24397 30920 24409 30923
rect 23348 30892 24409 30920
rect 23348 30880 23354 30892
rect 24397 30889 24409 30892
rect 24443 30889 24455 30923
rect 24397 30883 24455 30889
rect 17402 30852 17408 30864
rect 16776 30824 17408 30852
rect 16776 30793 16804 30824
rect 17402 30812 17408 30824
rect 17460 30812 17466 30864
rect 18693 30855 18751 30861
rect 18693 30821 18705 30855
rect 18739 30821 18751 30855
rect 18693 30815 18751 30821
rect 16761 30787 16819 30793
rect 16761 30753 16773 30787
rect 16807 30753 16819 30787
rect 18708 30784 18736 30815
rect 21269 30787 21327 30793
rect 21269 30784 21281 30787
rect 16761 30747 16819 30753
rect 16960 30756 18736 30784
rect 19260 30756 21281 30784
rect 16960 30725 16988 30756
rect 16945 30719 17003 30725
rect 16945 30685 16957 30719
rect 16991 30685 17003 30719
rect 16945 30679 17003 30685
rect 18141 30719 18199 30725
rect 18141 30685 18153 30719
rect 18187 30685 18199 30719
rect 18141 30679 18199 30685
rect 16942 30540 16948 30592
rect 17000 30580 17006 30592
rect 17129 30583 17187 30589
rect 17129 30580 17141 30583
rect 17000 30552 17141 30580
rect 17000 30540 17006 30552
rect 17129 30549 17141 30552
rect 17175 30549 17187 30583
rect 18156 30580 18184 30679
rect 18230 30676 18236 30728
rect 18288 30716 18294 30728
rect 18417 30719 18475 30725
rect 18417 30716 18429 30719
rect 18288 30688 18429 30716
rect 18288 30676 18294 30688
rect 18417 30685 18429 30688
rect 18463 30685 18475 30719
rect 18417 30679 18475 30685
rect 18509 30719 18567 30725
rect 18509 30685 18521 30719
rect 18555 30716 18567 30719
rect 18782 30716 18788 30728
rect 18555 30688 18788 30716
rect 18555 30685 18567 30688
rect 18509 30679 18567 30685
rect 18782 30676 18788 30688
rect 18840 30676 18846 30728
rect 19150 30676 19156 30728
rect 19208 30716 19214 30728
rect 19260 30725 19288 30756
rect 21269 30753 21281 30756
rect 21315 30753 21327 30787
rect 21542 30784 21548 30796
rect 21503 30756 21548 30784
rect 21269 30747 21327 30753
rect 19245 30719 19303 30725
rect 19245 30716 19257 30719
rect 19208 30688 19257 30716
rect 19208 30676 19214 30688
rect 19245 30685 19257 30688
rect 19291 30685 19303 30719
rect 19245 30679 19303 30685
rect 19521 30719 19579 30725
rect 19521 30685 19533 30719
rect 19567 30685 19579 30719
rect 19521 30679 19579 30685
rect 18322 30648 18328 30660
rect 18283 30620 18328 30648
rect 18322 30608 18328 30620
rect 18380 30608 18386 30660
rect 19242 30580 19248 30592
rect 18156 30552 19248 30580
rect 17129 30543 17187 30549
rect 19242 30540 19248 30552
rect 19300 30580 19306 30592
rect 19536 30580 19564 30679
rect 19300 30552 19564 30580
rect 19300 30540 19306 30552
rect 20070 30540 20076 30592
rect 20128 30580 20134 30592
rect 20622 30580 20628 30592
rect 20128 30552 20628 30580
rect 20128 30540 20134 30552
rect 20622 30540 20628 30552
rect 20680 30540 20686 30592
rect 21284 30580 21312 30747
rect 21542 30744 21548 30756
rect 21600 30744 21606 30796
rect 23293 30787 23351 30793
rect 23293 30753 23305 30787
rect 23339 30784 23351 30787
rect 23382 30784 23388 30796
rect 23339 30756 23388 30784
rect 23339 30753 23351 30756
rect 23293 30747 23351 30753
rect 23382 30744 23388 30756
rect 23440 30744 23446 30796
rect 24394 30744 24400 30796
rect 24452 30784 24458 30796
rect 25041 30787 25099 30793
rect 25041 30784 25053 30787
rect 24452 30756 25053 30784
rect 24452 30744 24458 30756
rect 25041 30753 25053 30756
rect 25087 30753 25099 30787
rect 25041 30747 25099 30753
rect 22094 30676 22100 30728
rect 22152 30716 22158 30728
rect 23017 30719 23075 30725
rect 23017 30716 23029 30719
rect 22152 30688 23029 30716
rect 22152 30676 22158 30688
rect 23017 30685 23029 30688
rect 23063 30685 23075 30719
rect 24578 30716 24584 30728
rect 24539 30688 24584 30716
rect 23017 30679 23075 30685
rect 24578 30676 24584 30688
rect 24636 30676 24642 30728
rect 25056 30716 25084 30747
rect 26418 30716 26424 30728
rect 25056 30688 26424 30716
rect 26418 30676 26424 30688
rect 26476 30676 26482 30728
rect 25308 30651 25366 30657
rect 25308 30617 25320 30651
rect 25354 30648 25366 30651
rect 26050 30648 26056 30660
rect 25354 30620 26056 30648
rect 25354 30617 25366 30620
rect 25308 30611 25366 30617
rect 26050 30608 26056 30620
rect 26108 30608 26114 30660
rect 23474 30580 23480 30592
rect 21284 30552 23480 30580
rect 23474 30540 23480 30552
rect 23532 30540 23538 30592
rect 26421 30583 26479 30589
rect 26421 30549 26433 30583
rect 26467 30580 26479 30583
rect 26602 30580 26608 30592
rect 26467 30552 26608 30580
rect 26467 30549 26479 30552
rect 26421 30543 26479 30549
rect 26602 30540 26608 30552
rect 26660 30540 26666 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 16758 30376 16764 30388
rect 16040 30348 16764 30376
rect 15933 30243 15991 30249
rect 15933 30209 15945 30243
rect 15979 30240 15991 30243
rect 16040 30240 16068 30348
rect 16758 30336 16764 30348
rect 16816 30336 16822 30388
rect 16850 30336 16856 30388
rect 16908 30336 16914 30388
rect 20254 30376 20260 30388
rect 20215 30348 20260 30376
rect 20254 30336 20260 30348
rect 20312 30336 20318 30388
rect 23290 30376 23296 30388
rect 23251 30348 23296 30376
rect 23290 30336 23296 30348
rect 23348 30336 23354 30388
rect 24026 30376 24032 30388
rect 23987 30348 24032 30376
rect 24026 30336 24032 30348
rect 24084 30336 24090 30388
rect 26234 30336 26240 30388
rect 26292 30376 26298 30388
rect 26329 30379 26387 30385
rect 26329 30376 26341 30379
rect 26292 30348 26341 30376
rect 26292 30336 26298 30348
rect 26329 30345 26341 30348
rect 26375 30345 26387 30379
rect 26329 30339 26387 30345
rect 16117 30311 16175 30317
rect 16117 30277 16129 30311
rect 16163 30308 16175 30311
rect 16868 30308 16896 30336
rect 16163 30280 16896 30308
rect 20165 30311 20223 30317
rect 16163 30277 16175 30280
rect 16117 30271 16175 30277
rect 20165 30277 20177 30311
rect 20211 30308 20223 30311
rect 20438 30308 20444 30320
rect 20211 30280 20444 30308
rect 20211 30277 20223 30280
rect 20165 30271 20223 30277
rect 20438 30268 20444 30280
rect 20496 30268 20502 30320
rect 22554 30308 22560 30320
rect 21836 30280 22560 30308
rect 15979 30212 16068 30240
rect 15979 30209 15991 30212
rect 15933 30203 15991 30209
rect 16758 30200 16764 30252
rect 16816 30240 16822 30252
rect 16925 30243 16983 30249
rect 16925 30240 16937 30243
rect 16816 30212 16937 30240
rect 16816 30200 16822 30212
rect 16925 30209 16937 30212
rect 16971 30209 16983 30243
rect 18782 30240 18788 30252
rect 18743 30212 18788 30240
rect 16925 30203 16983 30209
rect 18782 30200 18788 30212
rect 18840 30200 18846 30252
rect 21836 30249 21864 30280
rect 22554 30268 22560 30280
rect 22612 30268 22618 30320
rect 25225 30311 25283 30317
rect 25225 30277 25237 30311
rect 25271 30308 25283 30311
rect 26602 30308 26608 30320
rect 25271 30280 26608 30308
rect 25271 30277 25283 30280
rect 25225 30271 25283 30277
rect 26602 30268 26608 30280
rect 26660 30268 26666 30320
rect 21821 30243 21879 30249
rect 21821 30209 21833 30243
rect 21867 30209 21879 30243
rect 21821 30203 21879 30209
rect 22005 30243 22063 30249
rect 22005 30209 22017 30243
rect 22051 30240 22063 30243
rect 22186 30240 22192 30252
rect 22051 30212 22192 30240
rect 22051 30209 22063 30212
rect 22005 30203 22063 30209
rect 22186 30200 22192 30212
rect 22244 30200 22250 30252
rect 23201 30243 23259 30249
rect 23201 30209 23213 30243
rect 23247 30240 23259 30243
rect 23290 30240 23296 30252
rect 23247 30212 23296 30240
rect 23247 30209 23259 30212
rect 23201 30203 23259 30209
rect 23290 30200 23296 30212
rect 23348 30200 23354 30252
rect 24026 30200 24032 30252
rect 24084 30240 24090 30252
rect 24213 30243 24271 30249
rect 24213 30240 24225 30243
rect 24084 30212 24225 30240
rect 24084 30200 24090 30212
rect 24213 30209 24225 30212
rect 24259 30209 24271 30243
rect 24213 30203 24271 30209
rect 24854 30200 24860 30252
rect 24912 30240 24918 30252
rect 24949 30243 25007 30249
rect 24949 30240 24961 30243
rect 24912 30212 24961 30240
rect 24912 30200 24918 30212
rect 24949 30209 24961 30212
rect 24995 30209 25007 30243
rect 25130 30240 25136 30252
rect 25091 30212 25136 30240
rect 24949 30203 25007 30209
rect 25130 30200 25136 30212
rect 25188 30200 25194 30252
rect 25314 30200 25320 30252
rect 25372 30240 25378 30252
rect 26145 30243 26203 30249
rect 26145 30240 26157 30243
rect 25372 30212 25417 30240
rect 25516 30212 26157 30240
rect 25372 30200 25378 30212
rect 15749 30175 15807 30181
rect 15749 30141 15761 30175
rect 15795 30141 15807 30175
rect 16666 30172 16672 30184
rect 16627 30144 16672 30172
rect 15749 30135 15807 30141
rect 14734 29996 14740 30048
rect 14792 30036 14798 30048
rect 15764 30036 15792 30135
rect 16666 30132 16672 30144
rect 16724 30132 16730 30184
rect 18506 30172 18512 30184
rect 18419 30144 18512 30172
rect 18506 30132 18512 30144
rect 18564 30172 18570 30184
rect 20441 30175 20499 30181
rect 18564 30144 20024 30172
rect 18564 30132 18570 30144
rect 19426 30064 19432 30116
rect 19484 30104 19490 30116
rect 19797 30107 19855 30113
rect 19797 30104 19809 30107
rect 19484 30076 19809 30104
rect 19484 30064 19490 30076
rect 19797 30073 19809 30076
rect 19843 30073 19855 30107
rect 19996 30104 20024 30144
rect 20441 30141 20453 30175
rect 20487 30172 20499 30175
rect 21913 30175 21971 30181
rect 21913 30172 21925 30175
rect 20487 30144 21925 30172
rect 20487 30141 20499 30144
rect 20441 30135 20499 30141
rect 21913 30141 21925 30144
rect 21959 30141 21971 30175
rect 21913 30135 21971 30141
rect 23382 30132 23388 30184
rect 23440 30172 23446 30184
rect 23440 30144 23485 30172
rect 23440 30132 23446 30144
rect 22094 30104 22100 30116
rect 19996 30076 22100 30104
rect 19797 30067 19855 30073
rect 22094 30064 22100 30076
rect 22152 30064 22158 30116
rect 22833 30107 22891 30113
rect 22833 30073 22845 30107
rect 22879 30104 22891 30107
rect 23198 30104 23204 30116
rect 22879 30076 23204 30104
rect 22879 30073 22891 30076
rect 22833 30067 22891 30073
rect 23198 30064 23204 30076
rect 23256 30064 23262 30116
rect 25516 30113 25544 30212
rect 26145 30209 26157 30212
rect 26191 30209 26203 30243
rect 26145 30203 26203 30209
rect 27157 30243 27215 30249
rect 27157 30209 27169 30243
rect 27203 30240 27215 30243
rect 27522 30240 27528 30252
rect 27203 30212 27528 30240
rect 27203 30209 27215 30212
rect 27157 30203 27215 30209
rect 27522 30200 27528 30212
rect 27580 30200 27586 30252
rect 25961 30175 26019 30181
rect 25961 30172 25973 30175
rect 25884 30144 25973 30172
rect 25501 30107 25559 30113
rect 25501 30073 25513 30107
rect 25547 30073 25559 30107
rect 25501 30067 25559 30073
rect 17402 30036 17408 30048
rect 14792 30008 17408 30036
rect 14792 29996 14798 30008
rect 17402 29996 17408 30008
rect 17460 29996 17466 30048
rect 18049 30039 18107 30045
rect 18049 30005 18061 30039
rect 18095 30036 18107 30039
rect 18230 30036 18236 30048
rect 18095 30008 18236 30036
rect 18095 30005 18107 30008
rect 18049 29999 18107 30005
rect 18230 29996 18236 30008
rect 18288 29996 18294 30048
rect 23658 29996 23664 30048
rect 23716 30036 23722 30048
rect 25884 30036 25912 30144
rect 25961 30141 25973 30144
rect 26007 30172 26019 30175
rect 26970 30172 26976 30184
rect 26007 30144 26976 30172
rect 26007 30141 26019 30144
rect 25961 30135 26019 30141
rect 26970 30132 26976 30144
rect 27028 30132 27034 30184
rect 23716 30008 25912 30036
rect 27341 30039 27399 30045
rect 23716 29996 23722 30008
rect 27341 30005 27353 30039
rect 27387 30036 27399 30039
rect 28442 30036 28448 30048
rect 27387 30008 28448 30036
rect 27387 30005 27399 30008
rect 27341 29999 27399 30005
rect 28442 29996 28448 30008
rect 28500 29996 28506 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 14734 29832 14740 29844
rect 14695 29804 14740 29832
rect 14734 29792 14740 29804
rect 14792 29792 14798 29844
rect 16666 29832 16672 29844
rect 16408 29804 16672 29832
rect 15381 29767 15439 29773
rect 15381 29733 15393 29767
rect 15427 29764 15439 29767
rect 15562 29764 15568 29776
rect 15427 29736 15568 29764
rect 15427 29733 15439 29736
rect 15381 29727 15439 29733
rect 15562 29724 15568 29736
rect 15620 29724 15626 29776
rect 14642 29656 14648 29708
rect 14700 29696 14706 29708
rect 16408 29705 16436 29804
rect 16666 29792 16672 29804
rect 16724 29792 16730 29844
rect 18322 29792 18328 29844
rect 18380 29832 18386 29844
rect 19245 29835 19303 29841
rect 19245 29832 19257 29835
rect 18380 29804 19257 29832
rect 18380 29792 18386 29804
rect 19245 29801 19257 29804
rect 19291 29801 19303 29835
rect 20530 29832 20536 29844
rect 20491 29804 20536 29832
rect 19245 29795 19303 29801
rect 20530 29792 20536 29804
rect 20588 29792 20594 29844
rect 21913 29835 21971 29841
rect 21913 29801 21925 29835
rect 21959 29801 21971 29835
rect 21913 29795 21971 29801
rect 22097 29835 22155 29841
rect 22097 29801 22109 29835
rect 22143 29832 22155 29835
rect 22370 29832 22376 29844
rect 22143 29804 22376 29832
rect 22143 29801 22155 29804
rect 22097 29795 22155 29801
rect 21928 29764 21956 29795
rect 22370 29792 22376 29804
rect 22428 29792 22434 29844
rect 22741 29835 22799 29841
rect 22741 29801 22753 29835
rect 22787 29832 22799 29835
rect 23382 29832 23388 29844
rect 22787 29804 22821 29832
rect 23343 29804 23388 29832
rect 22787 29801 22799 29804
rect 22741 29795 22799 29801
rect 22756 29764 22784 29795
rect 23382 29792 23388 29804
rect 23440 29792 23446 29844
rect 24673 29835 24731 29841
rect 24673 29801 24685 29835
rect 24719 29832 24731 29835
rect 25130 29832 25136 29844
rect 24719 29804 25136 29832
rect 24719 29801 24731 29804
rect 24673 29795 24731 29801
rect 25130 29792 25136 29804
rect 25188 29792 25194 29844
rect 22830 29764 22836 29776
rect 21928 29736 22836 29764
rect 22830 29724 22836 29736
rect 22888 29724 22894 29776
rect 16393 29699 16451 29705
rect 16393 29696 16405 29699
rect 14700 29668 16405 29696
rect 14700 29656 14706 29668
rect 16393 29665 16405 29668
rect 16439 29665 16451 29699
rect 16393 29659 16451 29665
rect 19889 29699 19947 29705
rect 19889 29665 19901 29699
rect 19935 29696 19947 29699
rect 20622 29696 20628 29708
rect 19935 29668 20628 29696
rect 19935 29665 19947 29668
rect 19889 29659 19947 29665
rect 20622 29656 20628 29668
rect 20680 29656 20686 29708
rect 20990 29656 20996 29708
rect 21048 29696 21054 29708
rect 21085 29699 21143 29705
rect 21085 29696 21097 29699
rect 21048 29668 21097 29696
rect 21048 29656 21054 29668
rect 21085 29665 21097 29668
rect 21131 29665 21143 29699
rect 25222 29696 25228 29708
rect 25183 29668 25228 29696
rect 21085 29659 21143 29665
rect 25222 29656 25228 29668
rect 25280 29656 25286 29708
rect 26418 29696 26424 29708
rect 26379 29668 26424 29696
rect 26418 29656 26424 29668
rect 26476 29656 26482 29708
rect 14734 29588 14740 29640
rect 14792 29628 14798 29640
rect 16666 29637 16672 29640
rect 14921 29631 14979 29637
rect 14921 29628 14933 29631
rect 14792 29600 14933 29628
rect 14792 29588 14798 29600
rect 14921 29597 14933 29600
rect 14967 29597 14979 29631
rect 14921 29591 14979 29597
rect 15657 29631 15715 29637
rect 15657 29597 15669 29631
rect 15703 29597 15715 29631
rect 16660 29628 16672 29637
rect 16627 29600 16672 29628
rect 15657 29591 15715 29597
rect 16660 29591 16672 29600
rect 15286 29520 15292 29572
rect 15344 29560 15350 29572
rect 15381 29563 15439 29569
rect 15381 29560 15393 29563
rect 15344 29532 15393 29560
rect 15344 29520 15350 29532
rect 15381 29529 15393 29532
rect 15427 29529 15439 29563
rect 15672 29560 15700 29591
rect 16666 29588 16672 29591
rect 16724 29588 16730 29640
rect 19613 29631 19671 29637
rect 19613 29597 19625 29631
rect 19659 29628 19671 29631
rect 20254 29628 20260 29640
rect 19659 29600 20260 29628
rect 19659 29597 19671 29600
rect 19613 29591 19671 29597
rect 20254 29588 20260 29600
rect 20312 29628 20318 29640
rect 20901 29631 20959 29637
rect 20901 29628 20913 29631
rect 20312 29600 20913 29628
rect 20312 29588 20318 29600
rect 20901 29597 20913 29600
rect 20947 29597 20959 29631
rect 20901 29591 20959 29597
rect 23290 29588 23296 29640
rect 23348 29628 23354 29640
rect 23385 29631 23443 29637
rect 23385 29628 23397 29631
rect 23348 29600 23397 29628
rect 23348 29588 23354 29600
rect 23385 29597 23397 29600
rect 23431 29597 23443 29631
rect 23385 29591 23443 29597
rect 23569 29631 23627 29637
rect 23569 29597 23581 29631
rect 23615 29597 23627 29631
rect 28442 29628 28448 29640
rect 28403 29600 28448 29628
rect 23569 29591 23627 29597
rect 16574 29560 16580 29572
rect 15672 29532 16580 29560
rect 15381 29523 15439 29529
rect 16574 29520 16580 29532
rect 16632 29520 16638 29572
rect 21729 29563 21787 29569
rect 21729 29529 21741 29563
rect 21775 29560 21787 29563
rect 22557 29563 22615 29569
rect 22557 29560 22569 29563
rect 21775 29532 22569 29560
rect 21775 29529 21787 29532
rect 21729 29523 21787 29529
rect 22112 29504 22140 29532
rect 22557 29529 22569 29532
rect 22603 29529 22615 29563
rect 22557 29523 22615 29529
rect 23106 29520 23112 29572
rect 23164 29560 23170 29572
rect 23584 29560 23612 29591
rect 28442 29588 28448 29600
rect 28500 29588 28506 29640
rect 23164 29532 23612 29560
rect 25041 29563 25099 29569
rect 23164 29520 23170 29532
rect 25041 29529 25053 29563
rect 25087 29560 25099 29563
rect 26688 29563 26746 29569
rect 25087 29532 26648 29560
rect 25087 29529 25099 29532
rect 25041 29523 25099 29529
rect 26620 29504 26648 29532
rect 26688 29529 26700 29563
rect 26734 29560 26746 29563
rect 26734 29532 28304 29560
rect 26734 29529 26746 29532
rect 26688 29523 26746 29529
rect 14918 29452 14924 29504
rect 14976 29492 14982 29504
rect 15565 29495 15623 29501
rect 15565 29492 15577 29495
rect 14976 29464 15577 29492
rect 14976 29452 14982 29464
rect 15565 29461 15577 29464
rect 15611 29461 15623 29495
rect 15565 29455 15623 29461
rect 17773 29495 17831 29501
rect 17773 29461 17785 29495
rect 17819 29492 17831 29495
rect 18046 29492 18052 29504
rect 17819 29464 18052 29492
rect 17819 29461 17831 29464
rect 17773 29455 17831 29461
rect 18046 29452 18052 29464
rect 18104 29452 18110 29504
rect 18230 29452 18236 29504
rect 18288 29492 18294 29504
rect 19705 29495 19763 29501
rect 19705 29492 19717 29495
rect 18288 29464 19717 29492
rect 18288 29452 18294 29464
rect 19705 29461 19717 29464
rect 19751 29492 19763 29495
rect 20438 29492 20444 29504
rect 19751 29464 20444 29492
rect 19751 29461 19763 29464
rect 19705 29455 19763 29461
rect 20438 29452 20444 29464
rect 20496 29452 20502 29504
rect 20993 29495 21051 29501
rect 20993 29461 21005 29495
rect 21039 29492 21051 29495
rect 21082 29492 21088 29504
rect 21039 29464 21088 29492
rect 21039 29461 21051 29464
rect 20993 29455 21051 29461
rect 21082 29452 21088 29464
rect 21140 29492 21146 29504
rect 21634 29492 21640 29504
rect 21140 29464 21640 29492
rect 21140 29452 21146 29464
rect 21634 29452 21640 29464
rect 21692 29452 21698 29504
rect 21910 29452 21916 29504
rect 21968 29501 21974 29504
rect 21968 29495 21987 29501
rect 21975 29461 21987 29495
rect 21968 29455 21987 29461
rect 21968 29452 21974 29455
rect 22094 29452 22100 29504
rect 22152 29452 22158 29504
rect 22738 29452 22744 29504
rect 22796 29501 22802 29504
rect 22796 29495 22815 29501
rect 22803 29461 22815 29495
rect 22796 29455 22815 29461
rect 22925 29495 22983 29501
rect 22925 29461 22937 29495
rect 22971 29492 22983 29495
rect 24946 29492 24952 29504
rect 22971 29464 24952 29492
rect 22971 29461 22983 29464
rect 22925 29455 22983 29461
rect 22796 29452 22802 29455
rect 24946 29452 24952 29464
rect 25004 29452 25010 29504
rect 25133 29495 25191 29501
rect 25133 29461 25145 29495
rect 25179 29492 25191 29495
rect 25866 29492 25872 29504
rect 25179 29464 25872 29492
rect 25179 29461 25191 29464
rect 25133 29455 25191 29461
rect 25866 29452 25872 29464
rect 25924 29452 25930 29504
rect 26602 29452 26608 29504
rect 26660 29452 26666 29504
rect 27246 29452 27252 29504
rect 27304 29492 27310 29504
rect 28276 29501 28304 29532
rect 27801 29495 27859 29501
rect 27801 29492 27813 29495
rect 27304 29464 27813 29492
rect 27304 29452 27310 29464
rect 27801 29461 27813 29464
rect 27847 29461 27859 29495
rect 27801 29455 27859 29461
rect 28261 29495 28319 29501
rect 28261 29461 28273 29495
rect 28307 29461 28319 29495
rect 28261 29455 28319 29461
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 4614 29248 4620 29300
rect 4672 29288 4678 29300
rect 16758 29288 16764 29300
rect 4672 29260 16620 29288
rect 16719 29260 16764 29288
rect 4672 29248 4678 29260
rect 14642 29220 14648 29232
rect 14200 29192 14648 29220
rect 13078 29152 13084 29164
rect 13039 29124 13084 29152
rect 13078 29112 13084 29124
rect 13136 29112 13142 29164
rect 14200 29161 14228 29192
rect 14642 29180 14648 29192
rect 14700 29180 14706 29232
rect 16592 29220 16620 29260
rect 16758 29248 16764 29260
rect 16816 29248 16822 29300
rect 18138 29248 18144 29300
rect 18196 29288 18202 29300
rect 18601 29291 18659 29297
rect 18601 29288 18613 29291
rect 18196 29260 18613 29288
rect 18196 29248 18202 29260
rect 18601 29257 18613 29260
rect 18647 29257 18659 29291
rect 18601 29251 18659 29257
rect 19061 29291 19119 29297
rect 19061 29257 19073 29291
rect 19107 29288 19119 29291
rect 19889 29291 19947 29297
rect 19889 29288 19901 29291
rect 19107 29260 19901 29288
rect 19107 29257 19119 29260
rect 19061 29251 19119 29257
rect 19889 29257 19901 29260
rect 19935 29288 19947 29291
rect 20254 29288 20260 29300
rect 19935 29260 20260 29288
rect 19935 29257 19947 29260
rect 19889 29251 19947 29257
rect 20254 29248 20260 29260
rect 20312 29248 20318 29300
rect 20898 29248 20904 29300
rect 20956 29288 20962 29300
rect 21177 29291 21235 29297
rect 21177 29288 21189 29291
rect 20956 29260 21189 29288
rect 20956 29248 20962 29260
rect 21177 29257 21189 29260
rect 21223 29257 21235 29291
rect 22186 29288 22192 29300
rect 21177 29251 21235 29257
rect 21284 29260 22192 29288
rect 16592 29192 20116 29220
rect 14458 29161 14464 29164
rect 13265 29155 13323 29161
rect 13265 29121 13277 29155
rect 13311 29121 13323 29155
rect 13265 29115 13323 29121
rect 14185 29155 14243 29161
rect 14185 29121 14197 29155
rect 14231 29121 14243 29155
rect 14185 29115 14243 29121
rect 14452 29115 14464 29161
rect 14516 29152 14522 29164
rect 16942 29152 16948 29164
rect 14516 29124 14552 29152
rect 16903 29124 16948 29152
rect 12618 29044 12624 29096
rect 12676 29084 12682 29096
rect 13280 29084 13308 29115
rect 14458 29112 14464 29115
rect 14516 29112 14522 29124
rect 16942 29112 16948 29124
rect 17000 29112 17006 29164
rect 18046 29112 18052 29164
rect 18104 29152 18110 29164
rect 20088 29161 20116 29192
rect 18969 29155 19027 29161
rect 18969 29152 18981 29155
rect 18104 29124 18981 29152
rect 18104 29112 18110 29124
rect 18969 29121 18981 29124
rect 19015 29121 19027 29155
rect 18969 29115 19027 29121
rect 20073 29155 20131 29161
rect 20073 29121 20085 29155
rect 20119 29121 20131 29155
rect 20073 29115 20131 29121
rect 12676 29056 13308 29084
rect 12676 29044 12682 29056
rect 13280 29016 13308 29056
rect 19245 29087 19303 29093
rect 19245 29053 19257 29087
rect 19291 29053 19303 29087
rect 20088 29084 20116 29115
rect 20898 29112 20904 29164
rect 20956 29152 20962 29164
rect 21284 29161 21312 29260
rect 22186 29248 22192 29260
rect 22244 29288 22250 29300
rect 22849 29291 22907 29297
rect 22849 29288 22861 29291
rect 22244 29260 22861 29288
rect 22244 29248 22250 29260
rect 22849 29257 22861 29260
rect 22895 29288 22907 29291
rect 23014 29288 23020 29300
rect 22895 29257 22908 29288
rect 22975 29260 23020 29288
rect 22849 29251 22908 29257
rect 21821 29223 21879 29229
rect 21821 29189 21833 29223
rect 21867 29189 21879 29223
rect 21821 29183 21879 29189
rect 22037 29223 22095 29229
rect 22037 29189 22049 29223
rect 22083 29220 22095 29223
rect 22278 29220 22284 29232
rect 22083 29192 22284 29220
rect 22083 29189 22095 29192
rect 22037 29183 22095 29189
rect 21085 29155 21143 29161
rect 21085 29152 21097 29155
rect 20956 29124 21097 29152
rect 20956 29112 20962 29124
rect 21085 29121 21097 29124
rect 21131 29121 21143 29155
rect 21085 29115 21143 29121
rect 21269 29155 21327 29161
rect 21269 29121 21281 29155
rect 21315 29121 21327 29155
rect 21836 29152 21864 29183
rect 22278 29180 22284 29192
rect 22336 29180 22342 29232
rect 22649 29223 22707 29229
rect 22649 29189 22661 29223
rect 22695 29189 22707 29223
rect 22880 29220 22908 29251
rect 23014 29248 23020 29260
rect 23072 29248 23078 29300
rect 23658 29288 23664 29300
rect 23619 29260 23664 29288
rect 23658 29248 23664 29260
rect 23716 29248 23722 29300
rect 25593 29291 25651 29297
rect 25593 29257 25605 29291
rect 25639 29288 25651 29291
rect 27522 29288 27528 29300
rect 25639 29260 27200 29288
rect 27483 29260 27528 29288
rect 25639 29257 25651 29260
rect 25593 29251 25651 29257
rect 23106 29220 23112 29232
rect 22880 29192 23112 29220
rect 22649 29183 22707 29189
rect 22186 29152 22192 29164
rect 21836 29124 22192 29152
rect 21269 29115 21327 29121
rect 22186 29112 22192 29124
rect 22244 29152 22250 29164
rect 22664 29152 22692 29183
rect 23106 29180 23112 29192
rect 23164 29180 23170 29232
rect 24578 29220 24584 29232
rect 23768 29192 24584 29220
rect 22244 29124 22692 29152
rect 22244 29112 22250 29124
rect 23768 29084 23796 29192
rect 24578 29180 24584 29192
rect 24636 29180 24642 29232
rect 24946 29180 24952 29232
rect 25004 29220 25010 29232
rect 25004 29192 26280 29220
rect 25004 29180 25010 29192
rect 23845 29155 23903 29161
rect 23845 29121 23857 29155
rect 23891 29152 23903 29155
rect 24026 29152 24032 29164
rect 23891 29124 24032 29152
rect 23891 29121 23903 29124
rect 23845 29115 23903 29121
rect 24026 29112 24032 29124
rect 24084 29112 24090 29164
rect 25958 29152 25964 29164
rect 25919 29124 25964 29152
rect 25958 29112 25964 29124
rect 26016 29112 26022 29164
rect 20088 29056 23796 29084
rect 24305 29087 24363 29093
rect 19245 29047 19303 29053
rect 24305 29053 24317 29087
rect 24351 29053 24363 29087
rect 24305 29047 24363 29053
rect 24581 29087 24639 29093
rect 24581 29053 24593 29087
rect 24627 29084 24639 29087
rect 24854 29084 24860 29096
rect 24627 29056 24860 29084
rect 24627 29053 24639 29056
rect 24581 29047 24639 29053
rect 15565 29019 15623 29025
rect 13280 28988 14228 29016
rect 12434 28908 12440 28960
rect 12492 28948 12498 28960
rect 13081 28951 13139 28957
rect 13081 28948 13093 28951
rect 12492 28920 13093 28948
rect 12492 28908 12498 28920
rect 13081 28917 13093 28920
rect 13127 28917 13139 28951
rect 14200 28948 14228 28988
rect 15565 28985 15577 29019
rect 15611 29016 15623 29019
rect 16666 29016 16672 29028
rect 15611 28988 16672 29016
rect 15611 28985 15623 28988
rect 15565 28979 15623 28985
rect 16666 28976 16672 28988
rect 16724 28976 16730 29028
rect 19260 29016 19288 29047
rect 22189 29019 22247 29025
rect 22189 29016 22201 29019
rect 19260 28988 22201 29016
rect 22189 28985 22201 28988
rect 22235 28985 22247 29019
rect 22189 28979 22247 28985
rect 23474 28976 23480 29028
rect 23532 29016 23538 29028
rect 24320 29016 24348 29047
rect 24854 29044 24860 29056
rect 24912 29084 24918 29096
rect 24912 29056 25728 29084
rect 24912 29044 24918 29056
rect 25700 29028 25728 29056
rect 26050 29044 26056 29096
rect 26108 29084 26114 29096
rect 26252 29093 26280 29192
rect 26326 29180 26332 29232
rect 26384 29220 26390 29232
rect 26694 29220 26700 29232
rect 26384 29192 26700 29220
rect 26384 29180 26390 29192
rect 26694 29180 26700 29192
rect 26752 29220 26758 29232
rect 27172 29229 27200 29260
rect 27522 29248 27528 29260
rect 27580 29248 27586 29300
rect 27157 29223 27215 29229
rect 26752 29192 27108 29220
rect 26752 29180 26758 29192
rect 26973 29155 27031 29161
rect 26973 29152 26985 29155
rect 26804 29124 26985 29152
rect 26237 29087 26295 29093
rect 26108 29056 26153 29084
rect 26108 29044 26114 29056
rect 26237 29053 26249 29087
rect 26283 29053 26295 29087
rect 26237 29047 26295 29053
rect 24394 29016 24400 29028
rect 23532 28988 24400 29016
rect 23532 28976 23538 28988
rect 24394 28976 24400 28988
rect 24452 28976 24458 29028
rect 25682 28976 25688 29028
rect 25740 29016 25746 29028
rect 26804 29016 26832 29124
rect 26973 29121 26985 29124
rect 27019 29121 27031 29155
rect 27080 29152 27108 29192
rect 27157 29189 27169 29223
rect 27203 29189 27215 29223
rect 27157 29183 27215 29189
rect 27246 29152 27252 29164
rect 27080 29124 27252 29152
rect 26973 29115 27031 29121
rect 27246 29112 27252 29124
rect 27304 29112 27310 29164
rect 27341 29155 27399 29161
rect 27341 29121 27353 29155
rect 27387 29121 27399 29155
rect 27341 29115 27399 29121
rect 27356 29084 27384 29115
rect 25740 28988 26832 29016
rect 27264 29056 27384 29084
rect 25740 28976 25746 28988
rect 15654 28948 15660 28960
rect 14200 28920 15660 28948
rect 13081 28911 13139 28917
rect 15654 28908 15660 28920
rect 15712 28908 15718 28960
rect 22005 28951 22063 28957
rect 22005 28917 22017 28951
rect 22051 28948 22063 28951
rect 22830 28948 22836 28960
rect 22051 28920 22836 28948
rect 22051 28917 22063 28920
rect 22005 28911 22063 28917
rect 22830 28908 22836 28920
rect 22888 28908 22894 28960
rect 26142 28908 26148 28960
rect 26200 28948 26206 28960
rect 27264 28948 27292 29056
rect 26200 28920 27292 28948
rect 26200 28908 26206 28920
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 16574 28704 16580 28756
rect 16632 28744 16638 28756
rect 16669 28747 16727 28753
rect 16669 28744 16681 28747
rect 16632 28716 16681 28744
rect 16632 28704 16638 28716
rect 16669 28713 16681 28716
rect 16715 28713 16727 28747
rect 16669 28707 16727 28713
rect 20714 28704 20720 28756
rect 20772 28744 20778 28756
rect 20993 28747 21051 28753
rect 20993 28744 21005 28747
rect 20772 28716 21005 28744
rect 20772 28704 20778 28716
rect 20993 28713 21005 28716
rect 21039 28713 21051 28747
rect 20993 28707 21051 28713
rect 22097 28747 22155 28753
rect 22097 28713 22109 28747
rect 22143 28744 22155 28747
rect 22462 28744 22468 28756
rect 22143 28716 22468 28744
rect 22143 28713 22155 28716
rect 22097 28707 22155 28713
rect 22462 28704 22468 28716
rect 22520 28704 22526 28756
rect 23569 28747 23627 28753
rect 23569 28713 23581 28747
rect 23615 28744 23627 28747
rect 25222 28744 25228 28756
rect 23615 28716 25228 28744
rect 23615 28713 23627 28716
rect 23569 28707 23627 28713
rect 25222 28704 25228 28716
rect 25280 28704 25286 28756
rect 26326 28704 26332 28756
rect 26384 28744 26390 28756
rect 28537 28747 28595 28753
rect 28537 28744 28549 28747
rect 26384 28716 28549 28744
rect 26384 28704 26390 28716
rect 28537 28713 28549 28716
rect 28583 28713 28595 28747
rect 28537 28707 28595 28713
rect 20806 28676 20812 28688
rect 20732 28648 20812 28676
rect 12161 28611 12219 28617
rect 12161 28608 12173 28611
rect 9968 28580 12173 28608
rect 9968 28552 9996 28580
rect 12161 28577 12173 28580
rect 12207 28577 12219 28611
rect 12161 28571 12219 28577
rect 15838 28568 15844 28620
rect 15896 28608 15902 28620
rect 16761 28611 16819 28617
rect 16761 28608 16773 28611
rect 15896 28580 16773 28608
rect 15896 28568 15902 28580
rect 16761 28577 16773 28580
rect 16807 28577 16819 28611
rect 16761 28571 16819 28577
rect 19242 28568 19248 28620
rect 19300 28608 19306 28620
rect 19300 28580 19840 28608
rect 19300 28568 19306 28580
rect 8941 28543 8999 28549
rect 8941 28509 8953 28543
rect 8987 28540 8999 28543
rect 9950 28540 9956 28552
rect 8987 28512 9956 28540
rect 8987 28509 8999 28512
rect 8941 28503 8999 28509
rect 9950 28500 9956 28512
rect 10008 28500 10014 28552
rect 11054 28540 11060 28552
rect 11015 28512 11060 28540
rect 11054 28500 11060 28512
rect 11112 28500 11118 28552
rect 11146 28543 11204 28549
rect 11146 28509 11158 28543
rect 11192 28509 11204 28543
rect 11146 28503 11204 28509
rect 8386 28432 8392 28484
rect 8444 28472 8450 28484
rect 9186 28475 9244 28481
rect 9186 28472 9198 28475
rect 8444 28444 9198 28472
rect 8444 28432 8450 28444
rect 9186 28441 9198 28444
rect 9232 28441 9244 28475
rect 9186 28435 9244 28441
rect 9582 28432 9588 28484
rect 9640 28472 9646 28484
rect 11164 28472 11192 28503
rect 11238 28500 11244 28552
rect 11296 28540 11302 28552
rect 12434 28549 12440 28552
rect 11425 28543 11483 28549
rect 11296 28512 11341 28540
rect 11296 28500 11302 28512
rect 11425 28509 11437 28543
rect 11471 28509 11483 28543
rect 11425 28503 11483 28509
rect 12428 28503 12440 28549
rect 12492 28540 12498 28552
rect 14642 28540 14648 28552
rect 12492 28512 12528 28540
rect 14603 28512 14648 28540
rect 11330 28472 11336 28484
rect 9640 28444 10916 28472
rect 11164 28444 11336 28472
rect 9640 28432 9646 28444
rect 9766 28364 9772 28416
rect 9824 28404 9830 28416
rect 10321 28407 10379 28413
rect 10321 28404 10333 28407
rect 9824 28376 10333 28404
rect 9824 28364 9830 28376
rect 10321 28373 10333 28376
rect 10367 28373 10379 28407
rect 10778 28404 10784 28416
rect 10739 28376 10784 28404
rect 10321 28367 10379 28373
rect 10778 28364 10784 28376
rect 10836 28364 10842 28416
rect 10888 28404 10916 28444
rect 11330 28432 11336 28444
rect 11388 28432 11394 28484
rect 11440 28404 11468 28503
rect 12434 28500 12440 28503
rect 12492 28500 12498 28512
rect 14642 28500 14648 28512
rect 14700 28500 14706 28552
rect 16485 28543 16543 28549
rect 16485 28509 16497 28543
rect 16531 28509 16543 28543
rect 16485 28503 16543 28509
rect 14912 28475 14970 28481
rect 14912 28441 14924 28475
rect 14958 28472 14970 28475
rect 15102 28472 15108 28484
rect 14958 28444 15108 28472
rect 14958 28441 14970 28444
rect 14912 28435 14970 28441
rect 15102 28432 15108 28444
rect 15160 28432 15166 28484
rect 16500 28472 16528 28503
rect 16574 28500 16580 28552
rect 16632 28540 16638 28552
rect 19812 28549 19840 28580
rect 20732 28549 20760 28648
rect 20806 28636 20812 28648
rect 20864 28636 20870 28688
rect 21910 28676 21916 28688
rect 20916 28648 21916 28676
rect 20916 28608 20944 28648
rect 21910 28636 21916 28648
rect 21968 28636 21974 28688
rect 22002 28636 22008 28688
rect 22060 28676 22066 28688
rect 22060 28648 24716 28676
rect 22060 28636 22066 28648
rect 20824 28580 20944 28608
rect 20824 28549 20852 28580
rect 21450 28568 21456 28620
rect 21508 28608 21514 28620
rect 22646 28608 22652 28620
rect 21508 28580 22652 28608
rect 21508 28568 21514 28580
rect 22646 28568 22652 28580
rect 22704 28568 22710 28620
rect 24688 28617 24716 28648
rect 24673 28611 24731 28617
rect 24673 28577 24685 28611
rect 24719 28608 24731 28611
rect 24762 28608 24768 28620
rect 24719 28580 24768 28608
rect 24719 28577 24731 28580
rect 24673 28571 24731 28577
rect 24762 28568 24768 28580
rect 24820 28568 24826 28620
rect 26513 28611 26571 28617
rect 26513 28608 26525 28611
rect 24872 28580 26525 28608
rect 19613 28543 19671 28549
rect 16632 28512 16677 28540
rect 16632 28500 16638 28512
rect 19613 28509 19625 28543
rect 19659 28509 19671 28543
rect 19613 28503 19671 28509
rect 19797 28543 19855 28549
rect 19797 28509 19809 28543
rect 19843 28509 19855 28543
rect 19797 28503 19855 28509
rect 20717 28543 20775 28549
rect 20717 28509 20729 28543
rect 20763 28509 20775 28543
rect 20717 28503 20775 28509
rect 20809 28543 20867 28549
rect 20809 28509 20821 28543
rect 20855 28509 20867 28543
rect 20809 28503 20867 28509
rect 21821 28543 21879 28549
rect 21821 28509 21833 28543
rect 21867 28540 21879 28543
rect 22094 28540 22100 28552
rect 21867 28512 22100 28540
rect 21867 28509 21879 28512
rect 21821 28503 21879 28509
rect 17494 28472 17500 28484
rect 16040 28444 17500 28472
rect 16040 28416 16068 28444
rect 17494 28432 17500 28444
rect 17552 28432 17558 28484
rect 19628 28472 19656 28503
rect 22094 28500 22100 28512
rect 22152 28540 22158 28552
rect 22152 28512 22692 28540
rect 22152 28500 22158 28512
rect 19978 28472 19984 28484
rect 19628 28444 19984 28472
rect 19978 28432 19984 28444
rect 20036 28432 20042 28484
rect 20441 28475 20499 28481
rect 20441 28441 20453 28475
rect 20487 28472 20499 28475
rect 21082 28472 21088 28484
rect 20487 28444 21088 28472
rect 20487 28441 20499 28444
rect 20441 28435 20499 28441
rect 21082 28432 21088 28444
rect 21140 28472 21146 28484
rect 21545 28475 21603 28481
rect 21545 28472 21557 28475
rect 21140 28444 21557 28472
rect 21140 28432 21146 28444
rect 21545 28441 21557 28444
rect 21591 28472 21603 28475
rect 22557 28475 22615 28481
rect 22557 28472 22569 28475
rect 21591 28444 22569 28472
rect 21591 28441 21603 28444
rect 21545 28435 21603 28441
rect 22557 28441 22569 28444
rect 22603 28441 22615 28475
rect 22664 28472 22692 28512
rect 22738 28500 22744 28552
rect 22796 28540 22802 28552
rect 22925 28543 22983 28549
rect 22925 28540 22937 28543
rect 22796 28512 22937 28540
rect 22796 28500 22802 28512
rect 22925 28509 22937 28512
rect 22971 28509 22983 28543
rect 22925 28503 22983 28509
rect 23290 28500 23296 28552
rect 23348 28540 23354 28552
rect 23569 28543 23627 28549
rect 23569 28540 23581 28543
rect 23348 28512 23581 28540
rect 23348 28500 23354 28512
rect 23569 28509 23581 28512
rect 23615 28509 23627 28543
rect 23569 28503 23627 28509
rect 23658 28500 23664 28552
rect 23716 28540 23722 28552
rect 23753 28543 23811 28549
rect 23753 28540 23765 28543
rect 23716 28512 23765 28540
rect 23716 28500 23722 28512
rect 23753 28509 23765 28512
rect 23799 28509 23811 28543
rect 23753 28503 23811 28509
rect 23842 28500 23848 28552
rect 23900 28540 23906 28552
rect 24872 28540 24900 28580
rect 26513 28577 26525 28580
rect 26559 28577 26571 28611
rect 26513 28571 26571 28577
rect 23900 28512 24900 28540
rect 24949 28543 25007 28549
rect 23900 28500 23906 28512
rect 24949 28509 24961 28543
rect 24995 28540 25007 28543
rect 25314 28540 25320 28552
rect 24995 28512 25320 28540
rect 24995 28509 25007 28512
rect 24949 28503 25007 28509
rect 25314 28500 25320 28512
rect 25372 28500 25378 28552
rect 26418 28500 26424 28552
rect 26476 28540 26482 28552
rect 26878 28540 26884 28552
rect 26476 28512 26884 28540
rect 26476 28500 26482 28512
rect 26878 28500 26884 28512
rect 26936 28540 26942 28552
rect 27157 28543 27215 28549
rect 27157 28540 27169 28543
rect 26936 28512 27169 28540
rect 26936 28500 26942 28512
rect 27157 28509 27169 28512
rect 27203 28509 27215 28543
rect 27157 28503 27215 28509
rect 23109 28475 23167 28481
rect 22664 28444 22876 28472
rect 22557 28435 22615 28441
rect 13538 28404 13544 28416
rect 10888 28376 11468 28404
rect 13499 28376 13544 28404
rect 13538 28364 13544 28376
rect 13596 28364 13602 28416
rect 16022 28404 16028 28416
rect 15935 28376 16028 28404
rect 16022 28364 16028 28376
rect 16080 28364 16086 28416
rect 19705 28407 19763 28413
rect 19705 28373 19717 28407
rect 19751 28404 19763 28407
rect 20162 28404 20168 28416
rect 19751 28376 20168 28404
rect 19751 28373 19763 28376
rect 19705 28367 19763 28373
rect 20162 28364 20168 28376
rect 20220 28364 20226 28416
rect 20254 28364 20260 28416
rect 20312 28404 20318 28416
rect 20625 28407 20683 28413
rect 20625 28404 20637 28407
rect 20312 28376 20637 28404
rect 20312 28364 20318 28376
rect 20625 28373 20637 28376
rect 20671 28404 20683 28407
rect 21450 28404 21456 28416
rect 20671 28376 21456 28404
rect 20671 28373 20683 28376
rect 20625 28367 20683 28373
rect 21450 28364 21456 28376
rect 21508 28404 21514 28416
rect 21729 28407 21787 28413
rect 21729 28404 21741 28407
rect 21508 28376 21741 28404
rect 21508 28364 21514 28376
rect 21729 28373 21741 28376
rect 21775 28373 21787 28407
rect 21910 28404 21916 28416
rect 21871 28376 21916 28404
rect 21729 28367 21787 28373
rect 21910 28364 21916 28376
rect 21968 28364 21974 28416
rect 22646 28364 22652 28416
rect 22704 28404 22710 28416
rect 22848 28413 22876 28444
rect 23109 28441 23121 28475
rect 23155 28472 23167 28475
rect 23934 28472 23940 28484
rect 23155 28444 23940 28472
rect 23155 28441 23167 28444
rect 23109 28435 23167 28441
rect 23934 28432 23940 28444
rect 23992 28432 23998 28484
rect 25866 28432 25872 28484
rect 25924 28472 25930 28484
rect 27424 28475 27482 28481
rect 25924 28444 26464 28472
rect 25924 28432 25930 28444
rect 22741 28407 22799 28413
rect 22741 28404 22753 28407
rect 22704 28376 22753 28404
rect 22704 28364 22710 28376
rect 22741 28373 22753 28376
rect 22787 28373 22799 28407
rect 22741 28367 22799 28373
rect 22833 28407 22891 28413
rect 22833 28373 22845 28407
rect 22879 28404 22891 28407
rect 23014 28404 23020 28416
rect 22879 28376 23020 28404
rect 22879 28373 22891 28376
rect 22833 28367 22891 28373
rect 23014 28364 23020 28376
rect 23072 28364 23078 28416
rect 25961 28407 26019 28413
rect 25961 28373 25973 28407
rect 26007 28404 26019 28407
rect 26050 28404 26056 28416
rect 26007 28376 26056 28404
rect 26007 28373 26019 28376
rect 25961 28367 26019 28373
rect 26050 28364 26056 28376
rect 26108 28364 26114 28416
rect 26326 28404 26332 28416
rect 26287 28376 26332 28404
rect 26326 28364 26332 28376
rect 26384 28364 26390 28416
rect 26436 28413 26464 28444
rect 27424 28441 27436 28475
rect 27470 28472 27482 28475
rect 27798 28472 27804 28484
rect 27470 28444 27804 28472
rect 27470 28441 27482 28444
rect 27424 28435 27482 28441
rect 27798 28432 27804 28444
rect 27856 28432 27862 28484
rect 26421 28407 26479 28413
rect 26421 28373 26433 28407
rect 26467 28373 26479 28407
rect 26421 28367 26479 28373
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 13081 28203 13139 28209
rect 13081 28169 13093 28203
rect 13127 28169 13139 28203
rect 15102 28200 15108 28212
rect 15063 28172 15108 28200
rect 13081 28163 13139 28169
rect 9484 28135 9542 28141
rect 9484 28101 9496 28135
rect 9530 28132 9542 28135
rect 9674 28132 9680 28144
rect 9530 28104 9680 28132
rect 9530 28101 9542 28104
rect 9484 28095 9542 28101
rect 9674 28092 9680 28104
rect 9732 28092 9738 28144
rect 12710 28092 12716 28144
rect 12768 28132 12774 28144
rect 13096 28132 13124 28163
rect 15102 28160 15108 28172
rect 15160 28160 15166 28212
rect 17313 28203 17371 28209
rect 17313 28169 17325 28203
rect 17359 28200 17371 28203
rect 18506 28200 18512 28212
rect 17359 28172 18512 28200
rect 17359 28169 17371 28172
rect 17313 28163 17371 28169
rect 18506 28160 18512 28172
rect 18564 28160 18570 28212
rect 20622 28200 20628 28212
rect 20583 28172 20628 28200
rect 20622 28160 20628 28172
rect 20680 28160 20686 28212
rect 25314 28160 25320 28212
rect 25372 28200 25378 28212
rect 26142 28200 26148 28212
rect 25372 28172 26148 28200
rect 25372 28160 25378 28172
rect 26142 28160 26148 28172
rect 26200 28160 26206 28212
rect 27798 28200 27804 28212
rect 27759 28172 27804 28200
rect 27798 28160 27804 28172
rect 27856 28160 27862 28212
rect 13541 28135 13599 28141
rect 13541 28132 13553 28135
rect 12768 28104 13553 28132
rect 12768 28092 12774 28104
rect 13541 28101 13553 28104
rect 13587 28101 13599 28135
rect 13541 28095 13599 28101
rect 14182 28092 14188 28144
rect 14240 28132 14246 28144
rect 16022 28132 16028 28144
rect 14240 28104 14688 28132
rect 14240 28092 14246 28104
rect 8570 28064 8576 28076
rect 8531 28036 8576 28064
rect 8570 28024 8576 28036
rect 8628 28024 8634 28076
rect 8754 28064 8760 28076
rect 8715 28036 8760 28064
rect 8754 28024 8760 28036
rect 8812 28024 8818 28076
rect 11974 28073 11980 28076
rect 11968 28027 11980 28073
rect 12032 28064 12038 28076
rect 14660 28073 14688 28104
rect 15396 28104 16028 28132
rect 13725 28067 13783 28073
rect 12032 28036 12068 28064
rect 11974 28024 11980 28027
rect 12032 28024 12038 28036
rect 13725 28033 13737 28067
rect 13771 28033 13783 28067
rect 13725 28027 13783 28033
rect 14461 28067 14519 28073
rect 14461 28033 14473 28067
rect 14507 28033 14519 28067
rect 14461 28027 14519 28033
rect 14645 28067 14703 28073
rect 14645 28033 14657 28067
rect 14691 28033 14703 28067
rect 15286 28064 15292 28076
rect 15247 28036 15292 28064
rect 14645 28027 14703 28033
rect 9217 27999 9275 28005
rect 9217 27965 9229 27999
rect 9263 27965 9275 27999
rect 11701 27999 11759 28005
rect 11701 27996 11713 27999
rect 9217 27959 9275 27965
rect 10520 27968 11713 27996
rect 8573 27863 8631 27869
rect 8573 27829 8585 27863
rect 8619 27860 8631 27863
rect 9122 27860 9128 27872
rect 8619 27832 9128 27860
rect 8619 27829 8631 27832
rect 8573 27823 8631 27829
rect 9122 27820 9128 27832
rect 9180 27820 9186 27872
rect 9232 27860 9260 27959
rect 10520 27872 10548 27968
rect 11701 27965 11713 27968
rect 11747 27965 11759 27999
rect 11701 27959 11759 27965
rect 13538 27956 13544 28008
rect 13596 27996 13602 28008
rect 13740 27996 13768 28027
rect 13596 27968 13768 27996
rect 13596 27956 13602 27968
rect 14476 27928 14504 28027
rect 15286 28024 15292 28036
rect 15344 28024 15350 28076
rect 15396 28073 15424 28104
rect 16022 28092 16028 28104
rect 16080 28092 16086 28144
rect 23658 28132 23664 28144
rect 22296 28104 23664 28132
rect 22296 28076 22324 28104
rect 23658 28092 23664 28104
rect 23716 28092 23722 28144
rect 26050 28132 26056 28144
rect 26011 28104 26056 28132
rect 26050 28092 26056 28104
rect 26108 28092 26114 28144
rect 26160 28132 26188 28160
rect 26160 28104 26280 28132
rect 15381 28067 15439 28073
rect 15381 28033 15393 28067
rect 15427 28033 15439 28067
rect 15562 28064 15568 28076
rect 15523 28036 15568 28064
rect 15381 28027 15439 28033
rect 15562 28024 15568 28036
rect 15620 28024 15626 28076
rect 15654 28024 15660 28076
rect 15712 28064 15718 28076
rect 15712 28036 15757 28064
rect 15712 28024 15718 28036
rect 15930 28024 15936 28076
rect 15988 28064 15994 28076
rect 16669 28067 16727 28073
rect 16669 28064 16681 28067
rect 15988 28036 16681 28064
rect 15988 28024 15994 28036
rect 16669 28033 16681 28036
rect 16715 28033 16727 28067
rect 16850 28064 16856 28076
rect 16811 28036 16856 28064
rect 16669 28027 16727 28033
rect 16850 28024 16856 28036
rect 16908 28024 16914 28076
rect 17126 28024 17132 28076
rect 17184 28064 17190 28076
rect 17497 28067 17555 28073
rect 17497 28064 17509 28067
rect 17184 28036 17509 28064
rect 17184 28024 17190 28036
rect 17497 28033 17509 28036
rect 17543 28033 17555 28067
rect 18598 28064 18604 28076
rect 18559 28036 18604 28064
rect 17497 28027 17555 28033
rect 18598 28024 18604 28036
rect 18656 28024 18662 28076
rect 18785 28067 18843 28073
rect 18785 28033 18797 28067
rect 18831 28033 18843 28067
rect 19334 28064 19340 28076
rect 19295 28036 19340 28064
rect 18785 28027 18843 28033
rect 14553 27999 14611 28005
rect 14553 27965 14565 27999
rect 14599 27996 14611 27999
rect 15304 27996 15332 28024
rect 17770 27996 17776 28008
rect 14599 27968 15332 27996
rect 17731 27968 17776 27996
rect 14599 27965 14611 27968
rect 14553 27959 14611 27965
rect 17770 27956 17776 27968
rect 17828 27956 17834 28008
rect 18800 27996 18828 28027
rect 19334 28024 19340 28036
rect 19392 28024 19398 28076
rect 20162 28064 20168 28076
rect 20075 28036 20168 28064
rect 20162 28024 20168 28036
rect 20220 28064 20226 28076
rect 20441 28067 20499 28073
rect 20220 28036 20392 28064
rect 20220 28024 20226 28036
rect 19242 27996 19248 28008
rect 17972 27968 19248 27996
rect 15562 27928 15568 27940
rect 14476 27900 15568 27928
rect 15562 27888 15568 27900
rect 15620 27888 15626 27940
rect 17972 27872 18000 27968
rect 19242 27956 19248 27968
rect 19300 27996 19306 28008
rect 19521 27999 19579 28005
rect 19521 27996 19533 27999
rect 19300 27968 19533 27996
rect 19300 27956 19306 27968
rect 19521 27965 19533 27968
rect 19567 27965 19579 27999
rect 19521 27959 19579 27965
rect 20257 27999 20315 28005
rect 20257 27965 20269 27999
rect 20303 27965 20315 27999
rect 20364 27996 20392 28036
rect 20441 28033 20453 28067
rect 20487 28064 20499 28067
rect 21082 28064 21088 28076
rect 20487 28036 21088 28064
rect 20487 28033 20499 28036
rect 20441 28027 20499 28033
rect 21082 28024 21088 28036
rect 21140 28024 21146 28076
rect 21266 28064 21272 28076
rect 21227 28036 21272 28064
rect 21266 28024 21272 28036
rect 21324 28024 21330 28076
rect 22097 28067 22155 28073
rect 22097 28033 22109 28067
rect 22143 28064 22155 28067
rect 22278 28064 22284 28076
rect 22143 28036 22284 28064
rect 22143 28033 22155 28036
rect 22097 28027 22155 28033
rect 22278 28024 22284 28036
rect 22336 28024 22342 28076
rect 23750 28064 23756 28076
rect 23711 28036 23756 28064
rect 23750 28024 23756 28036
rect 23808 28024 23814 28076
rect 23845 28067 23903 28073
rect 23845 28033 23857 28067
rect 23891 28064 23903 28067
rect 24578 28064 24584 28076
rect 23891 28036 24584 28064
rect 23891 28033 23903 28036
rect 23845 28027 23903 28033
rect 24578 28024 24584 28036
rect 24636 28024 24642 28076
rect 25682 28024 25688 28076
rect 25740 28064 25746 28076
rect 26252 28073 26280 28104
rect 25869 28067 25927 28073
rect 25869 28064 25881 28067
rect 25740 28036 25881 28064
rect 25740 28024 25746 28036
rect 25869 28033 25881 28036
rect 25915 28033 25927 28067
rect 25869 28027 25927 28033
rect 26145 28067 26203 28073
rect 26145 28033 26157 28067
rect 26191 28033 26203 28067
rect 26145 28027 26203 28033
rect 26237 28067 26295 28073
rect 26237 28033 26249 28067
rect 26283 28033 26295 28067
rect 26970 28064 26976 28076
rect 26931 28036 26976 28064
rect 26237 28027 26295 28033
rect 20622 27996 20628 28008
rect 20364 27968 20628 27996
rect 20257 27959 20315 27965
rect 18601 27931 18659 27937
rect 18601 27897 18613 27931
rect 18647 27928 18659 27931
rect 18647 27900 19334 27928
rect 18647 27897 18659 27900
rect 18601 27891 18659 27897
rect 9950 27860 9956 27872
rect 9232 27832 9956 27860
rect 9950 27820 9956 27832
rect 10008 27860 10014 27872
rect 10502 27860 10508 27872
rect 10008 27832 10508 27860
rect 10008 27820 10014 27832
rect 10502 27820 10508 27832
rect 10560 27820 10566 27872
rect 10594 27820 10600 27872
rect 10652 27860 10658 27872
rect 13909 27863 13967 27869
rect 10652 27832 10697 27860
rect 10652 27820 10658 27832
rect 13909 27829 13921 27863
rect 13955 27860 13967 27863
rect 13998 27860 14004 27872
rect 13955 27832 14004 27860
rect 13955 27829 13967 27832
rect 13909 27823 13967 27829
rect 13998 27820 14004 27832
rect 14056 27820 14062 27872
rect 14550 27820 14556 27872
rect 14608 27860 14614 27872
rect 16761 27863 16819 27869
rect 16761 27860 16773 27863
rect 14608 27832 16773 27860
rect 14608 27820 14614 27832
rect 16761 27829 16773 27832
rect 16807 27829 16819 27863
rect 16761 27823 16819 27829
rect 17681 27863 17739 27869
rect 17681 27829 17693 27863
rect 17727 27860 17739 27863
rect 17954 27860 17960 27872
rect 17727 27832 17960 27860
rect 17727 27829 17739 27832
rect 17681 27823 17739 27829
rect 17954 27820 17960 27832
rect 18012 27820 18018 27872
rect 19306 27860 19334 27900
rect 20070 27860 20076 27872
rect 19306 27832 20076 27860
rect 20070 27820 20076 27832
rect 20128 27860 20134 27872
rect 20165 27863 20223 27869
rect 20165 27860 20177 27863
rect 20128 27832 20177 27860
rect 20128 27820 20134 27832
rect 20165 27829 20177 27832
rect 20211 27829 20223 27863
rect 20272 27860 20300 27959
rect 20622 27956 20628 27968
rect 20680 27956 20686 28008
rect 21726 27956 21732 28008
rect 21784 27996 21790 28008
rect 21821 27999 21879 28005
rect 21821 27996 21833 27999
rect 21784 27968 21833 27996
rect 21784 27956 21790 27968
rect 21821 27965 21833 27968
rect 21867 27996 21879 27999
rect 21910 27996 21916 28008
rect 21867 27968 21916 27996
rect 21867 27965 21879 27968
rect 21821 27959 21879 27965
rect 21910 27956 21916 27968
rect 21968 27956 21974 28008
rect 23934 27956 23940 28008
rect 23992 27996 23998 28008
rect 24857 27999 24915 28005
rect 23992 27968 24037 27996
rect 23992 27956 23998 27968
rect 24857 27965 24869 27999
rect 24903 27996 24915 27999
rect 25774 27996 25780 28008
rect 24903 27968 25780 27996
rect 24903 27965 24915 27968
rect 24857 27959 24915 27965
rect 25774 27956 25780 27968
rect 25832 27956 25838 28008
rect 26160 27996 26188 28027
rect 26970 28024 26976 28036
rect 27028 28024 27034 28076
rect 27157 28067 27215 28073
rect 27157 28033 27169 28067
rect 27203 28033 27215 28067
rect 27157 28027 27215 28033
rect 27341 28067 27399 28073
rect 27341 28033 27353 28067
rect 27387 28064 27399 28067
rect 27985 28067 28043 28073
rect 27985 28064 27997 28067
rect 27387 28036 27997 28064
rect 27387 28033 27399 28036
rect 27341 28027 27399 28033
rect 27985 28033 27997 28036
rect 28031 28033 28043 28067
rect 27985 28027 28043 28033
rect 26326 27996 26332 28008
rect 26160 27968 26332 27996
rect 26326 27956 26332 27968
rect 26384 27956 26390 28008
rect 26421 27931 26479 27937
rect 26421 27897 26433 27931
rect 26467 27928 26479 27931
rect 27172 27928 27200 28027
rect 26467 27900 27200 27928
rect 26467 27897 26479 27900
rect 26421 27891 26479 27897
rect 20714 27860 20720 27872
rect 20272 27832 20720 27860
rect 20165 27823 20223 27829
rect 20714 27820 20720 27832
rect 20772 27820 20778 27872
rect 21082 27860 21088 27872
rect 21043 27832 21088 27860
rect 21082 27820 21088 27832
rect 21140 27820 21146 27872
rect 23385 27863 23443 27869
rect 23385 27829 23397 27863
rect 23431 27860 23443 27863
rect 24578 27860 24584 27872
rect 23431 27832 24584 27860
rect 23431 27829 23443 27832
rect 23385 27823 23443 27829
rect 24578 27820 24584 27832
rect 24636 27820 24642 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 8386 27656 8392 27668
rect 8347 27628 8392 27656
rect 8386 27616 8392 27628
rect 8444 27616 8450 27668
rect 15838 27656 15844 27668
rect 15799 27628 15844 27656
rect 15838 27616 15844 27628
rect 15896 27616 15902 27668
rect 17954 27656 17960 27668
rect 16500 27628 17960 27656
rect 9674 27588 9680 27600
rect 9635 27560 9680 27588
rect 9674 27548 9680 27560
rect 9732 27548 9738 27600
rect 14185 27591 14243 27597
rect 14185 27557 14197 27591
rect 14231 27588 14243 27591
rect 16500 27588 16528 27628
rect 17954 27616 17960 27628
rect 18012 27616 18018 27668
rect 20070 27616 20076 27668
rect 20128 27656 20134 27668
rect 20533 27659 20591 27665
rect 20533 27656 20545 27659
rect 20128 27628 20545 27656
rect 20128 27616 20134 27628
rect 20533 27625 20545 27628
rect 20579 27656 20591 27659
rect 21726 27656 21732 27668
rect 20579 27628 21732 27656
rect 20579 27625 20591 27628
rect 20533 27619 20591 27625
rect 21726 27616 21732 27628
rect 21784 27616 21790 27668
rect 22186 27616 22192 27668
rect 22244 27656 22250 27668
rect 22925 27659 22983 27665
rect 22925 27656 22937 27659
rect 22244 27628 22937 27656
rect 22244 27616 22250 27628
rect 22925 27625 22937 27628
rect 22971 27625 22983 27659
rect 23290 27656 23296 27668
rect 23251 27628 23296 27656
rect 22925 27619 22983 27625
rect 23290 27616 23296 27628
rect 23348 27616 23354 27668
rect 14231 27560 16528 27588
rect 14231 27557 14243 27560
rect 14185 27551 14243 27557
rect 8110 27480 8116 27532
rect 8168 27520 8174 27532
rect 8205 27523 8263 27529
rect 8205 27520 8217 27523
rect 8168 27492 8217 27520
rect 8168 27480 8174 27492
rect 8205 27489 8217 27492
rect 8251 27520 8263 27523
rect 9309 27523 9367 27529
rect 9309 27520 9321 27523
rect 8251 27492 9321 27520
rect 8251 27489 8263 27492
rect 8205 27483 8263 27489
rect 9309 27489 9321 27492
rect 9355 27489 9367 27523
rect 10318 27520 10324 27532
rect 9309 27483 9367 27489
rect 9508 27492 10324 27520
rect 8018 27452 8024 27464
rect 7979 27424 8024 27452
rect 8018 27412 8024 27424
rect 8076 27412 8082 27464
rect 8389 27455 8447 27461
rect 8389 27421 8401 27455
rect 8435 27421 8447 27455
rect 8938 27452 8944 27464
rect 8899 27424 8944 27452
rect 8389 27415 8447 27421
rect 8404 27384 8432 27415
rect 8938 27412 8944 27424
rect 8996 27412 9002 27464
rect 9122 27452 9128 27464
rect 9083 27424 9128 27452
rect 9122 27412 9128 27424
rect 9180 27412 9186 27464
rect 9214 27412 9220 27464
rect 9272 27452 9278 27464
rect 9508 27461 9536 27492
rect 10318 27480 10324 27492
rect 10376 27520 10382 27532
rect 10594 27520 10600 27532
rect 10376 27492 10600 27520
rect 10376 27480 10382 27492
rect 10594 27480 10600 27492
rect 10652 27480 10658 27532
rect 12710 27520 12716 27532
rect 12671 27492 12716 27520
rect 12710 27480 12716 27492
rect 12768 27480 12774 27532
rect 13538 27480 13544 27532
rect 13596 27520 13602 27532
rect 14369 27523 14427 27529
rect 14369 27520 14381 27523
rect 13596 27492 14381 27520
rect 13596 27480 13602 27492
rect 14369 27489 14381 27492
rect 14415 27489 14427 27523
rect 14369 27483 14427 27489
rect 15286 27480 15292 27532
rect 15344 27520 15350 27532
rect 15749 27523 15807 27529
rect 15749 27520 15761 27523
rect 15344 27492 15761 27520
rect 15344 27480 15350 27492
rect 15749 27489 15761 27492
rect 15795 27489 15807 27523
rect 17972 27520 18000 27616
rect 19426 27548 19432 27600
rect 19484 27548 19490 27600
rect 20990 27588 20996 27600
rect 20951 27560 20996 27588
rect 20990 27548 20996 27560
rect 21048 27548 21054 27600
rect 21082 27548 21088 27600
rect 21140 27588 21146 27600
rect 21913 27591 21971 27597
rect 21913 27588 21925 27591
rect 21140 27560 21925 27588
rect 21140 27548 21146 27560
rect 21913 27557 21925 27560
rect 21959 27557 21971 27591
rect 21913 27551 21971 27557
rect 22465 27591 22523 27597
rect 22465 27557 22477 27591
rect 22511 27588 22523 27591
rect 23842 27588 23848 27600
rect 22511 27560 23848 27588
rect 22511 27557 22523 27560
rect 22465 27551 22523 27557
rect 23842 27548 23848 27560
rect 23900 27548 23906 27600
rect 28166 27588 28172 27600
rect 25976 27560 28172 27588
rect 18693 27523 18751 27529
rect 15749 27483 15807 27489
rect 16316 27492 16614 27520
rect 17972 27492 18552 27520
rect 9493 27455 9551 27461
rect 9272 27424 9317 27452
rect 9272 27412 9278 27424
rect 9493 27421 9505 27455
rect 9539 27421 9551 27455
rect 9493 27415 9551 27421
rect 10502 27412 10508 27464
rect 10560 27452 10566 27464
rect 10689 27455 10747 27461
rect 10689 27452 10701 27455
rect 10560 27424 10701 27452
rect 10560 27412 10566 27424
rect 10689 27421 10701 27424
rect 10735 27421 10747 27455
rect 10689 27415 10747 27421
rect 10778 27412 10784 27464
rect 10836 27452 10842 27464
rect 10945 27455 11003 27461
rect 10945 27452 10957 27455
rect 10836 27424 10957 27452
rect 10836 27412 10842 27424
rect 10945 27421 10957 27424
rect 10991 27421 11003 27455
rect 12986 27452 12992 27464
rect 12947 27424 12992 27452
rect 10945 27415 11003 27421
rect 12986 27412 12992 27424
rect 13044 27452 13050 27464
rect 14093 27455 14151 27461
rect 14093 27452 14105 27455
rect 13044 27424 14105 27452
rect 13044 27412 13050 27424
rect 14093 27421 14105 27424
rect 14139 27421 14151 27455
rect 14093 27415 14151 27421
rect 14829 27455 14887 27461
rect 14829 27421 14841 27455
rect 14875 27421 14887 27455
rect 14829 27415 14887 27421
rect 15473 27455 15531 27461
rect 15473 27421 15485 27455
rect 15519 27452 15531 27455
rect 16316 27452 16344 27492
rect 16482 27452 16488 27464
rect 15519 27424 16344 27452
rect 16443 27424 16488 27452
rect 15519 27421 15531 27424
rect 15473 27415 15531 27421
rect 9858 27384 9864 27396
rect 8404 27356 9864 27384
rect 9858 27344 9864 27356
rect 9916 27344 9922 27396
rect 12250 27344 12256 27396
rect 12308 27384 12314 27396
rect 14844 27384 14872 27415
rect 16482 27412 16488 27424
rect 16540 27412 16546 27464
rect 16586 27452 16614 27492
rect 16586 27424 16896 27452
rect 16868 27396 16896 27424
rect 17310 27412 17316 27464
rect 17368 27452 17374 27464
rect 17770 27452 17776 27464
rect 17368 27424 17776 27452
rect 17368 27412 17374 27424
rect 17770 27412 17776 27424
rect 17828 27452 17834 27464
rect 18524 27461 18552 27492
rect 18693 27489 18705 27523
rect 18739 27520 18751 27523
rect 19150 27520 19156 27532
rect 18739 27492 19156 27520
rect 18739 27489 18751 27492
rect 18693 27483 18751 27489
rect 19150 27480 19156 27492
rect 19208 27480 19214 27532
rect 19444 27520 19472 27548
rect 19521 27523 19579 27529
rect 19521 27520 19533 27523
rect 19444 27492 19533 27520
rect 19521 27489 19533 27492
rect 19567 27489 19579 27523
rect 19521 27483 19579 27489
rect 19797 27523 19855 27529
rect 19797 27489 19809 27523
rect 19843 27520 19855 27523
rect 19978 27520 19984 27532
rect 19843 27492 19984 27520
rect 19843 27489 19855 27492
rect 19797 27483 19855 27489
rect 19978 27480 19984 27492
rect 20036 27480 20042 27532
rect 22002 27480 22008 27532
rect 22060 27520 22066 27532
rect 23017 27523 23075 27529
rect 23017 27520 23029 27523
rect 22060 27492 23029 27520
rect 22060 27480 22066 27492
rect 23017 27489 23029 27492
rect 23063 27489 23075 27523
rect 23017 27483 23075 27489
rect 18325 27455 18383 27461
rect 18325 27452 18337 27455
rect 17828 27424 18337 27452
rect 17828 27412 17834 27424
rect 18325 27421 18337 27424
rect 18371 27421 18383 27455
rect 18325 27415 18383 27421
rect 18509 27455 18567 27461
rect 18509 27421 18521 27455
rect 18555 27421 18567 27455
rect 18509 27415 18567 27421
rect 18966 27412 18972 27464
rect 19024 27452 19030 27464
rect 19429 27455 19487 27461
rect 19429 27452 19441 27455
rect 19024 27424 19441 27452
rect 19024 27412 19030 27424
rect 19429 27421 19441 27424
rect 19475 27421 19487 27455
rect 20714 27452 20720 27464
rect 20675 27424 20720 27452
rect 19429 27415 19487 27421
rect 20714 27412 20720 27424
rect 20772 27412 20778 27464
rect 20809 27455 20867 27461
rect 20809 27421 20821 27455
rect 20855 27452 20867 27455
rect 21082 27452 21088 27464
rect 20855 27424 21088 27452
rect 20855 27421 20867 27424
rect 20809 27415 20867 27421
rect 21082 27412 21088 27424
rect 21140 27452 21146 27464
rect 21266 27452 21272 27464
rect 21140 27424 21272 27452
rect 21140 27412 21146 27424
rect 21266 27412 21272 27424
rect 21324 27412 21330 27464
rect 22186 27452 22192 27464
rect 22147 27424 22192 27452
rect 22186 27412 22192 27424
rect 22244 27412 22250 27464
rect 22281 27455 22339 27461
rect 22281 27421 22293 27455
rect 22327 27452 22339 27455
rect 22738 27452 22744 27464
rect 22327 27424 22744 27452
rect 22327 27421 22339 27424
rect 22281 27415 22339 27421
rect 22738 27412 22744 27424
rect 22796 27412 22802 27464
rect 22922 27452 22928 27464
rect 22883 27424 22928 27452
rect 22922 27412 22928 27424
rect 22980 27412 22986 27464
rect 24394 27452 24400 27464
rect 24355 27424 24400 27452
rect 24394 27412 24400 27424
rect 24452 27412 24458 27464
rect 24578 27452 24584 27464
rect 24539 27424 24584 27452
rect 24578 27412 24584 27424
rect 24636 27412 24642 27464
rect 24762 27452 24768 27464
rect 24723 27424 24768 27452
rect 24762 27412 24768 27424
rect 24820 27412 24826 27464
rect 25682 27452 25688 27464
rect 25643 27424 25688 27452
rect 25682 27412 25688 27424
rect 25740 27412 25746 27464
rect 25774 27412 25780 27464
rect 25832 27452 25838 27464
rect 25976 27461 26004 27560
rect 28166 27548 28172 27560
rect 28224 27548 28230 27600
rect 26697 27523 26755 27529
rect 26697 27489 26709 27523
rect 26743 27520 26755 27523
rect 26970 27520 26976 27532
rect 26743 27492 26976 27520
rect 26743 27489 26755 27492
rect 26697 27483 26755 27489
rect 26970 27480 26976 27492
rect 27028 27480 27034 27532
rect 25961 27455 26019 27461
rect 25961 27452 25973 27455
rect 25832 27424 25973 27452
rect 25832 27412 25838 27424
rect 25961 27421 25973 27424
rect 26007 27421 26019 27455
rect 25961 27415 26019 27421
rect 26053 27455 26111 27461
rect 26053 27421 26065 27455
rect 26099 27452 26111 27455
rect 26142 27452 26148 27464
rect 26099 27424 26148 27452
rect 26099 27421 26111 27424
rect 26053 27415 26111 27421
rect 26142 27412 26148 27424
rect 26200 27412 26206 27464
rect 26881 27455 26939 27461
rect 26881 27421 26893 27455
rect 26927 27421 26939 27455
rect 26881 27415 26939 27421
rect 27709 27455 27767 27461
rect 27709 27421 27721 27455
rect 27755 27452 27767 27455
rect 28350 27452 28356 27464
rect 27755 27424 28356 27452
rect 27755 27421 27767 27424
rect 27709 27415 27767 27421
rect 12308 27356 14872 27384
rect 12308 27344 12314 27356
rect 16114 27344 16120 27396
rect 16172 27384 16178 27396
rect 16730 27387 16788 27393
rect 16730 27384 16742 27387
rect 16172 27356 16742 27384
rect 16172 27344 16178 27356
rect 16730 27353 16742 27356
rect 16776 27353 16788 27387
rect 16730 27347 16788 27353
rect 16850 27344 16856 27396
rect 16908 27344 16914 27396
rect 20533 27387 20591 27393
rect 20533 27353 20545 27387
rect 20579 27384 20591 27387
rect 20622 27384 20628 27396
rect 20579 27356 20628 27384
rect 20579 27353 20591 27356
rect 20533 27347 20591 27353
rect 20622 27344 20628 27356
rect 20680 27344 20686 27396
rect 22097 27387 22155 27393
rect 22097 27353 22109 27387
rect 22143 27384 22155 27387
rect 22646 27384 22652 27396
rect 22143 27356 22652 27384
rect 22143 27353 22155 27356
rect 22097 27347 22155 27353
rect 22646 27344 22652 27356
rect 22704 27344 22710 27396
rect 23750 27344 23756 27396
rect 23808 27384 23814 27396
rect 24673 27387 24731 27393
rect 24673 27384 24685 27387
rect 23808 27356 24685 27384
rect 23808 27344 23814 27356
rect 24673 27353 24685 27356
rect 24719 27384 24731 27387
rect 25222 27384 25228 27396
rect 24719 27356 25228 27384
rect 24719 27353 24731 27356
rect 24673 27347 24731 27353
rect 25222 27344 25228 27356
rect 25280 27344 25286 27396
rect 25498 27344 25504 27396
rect 25556 27384 25562 27396
rect 25869 27387 25927 27393
rect 25869 27384 25881 27387
rect 25556 27356 25881 27384
rect 25556 27344 25562 27356
rect 25869 27353 25881 27356
rect 25915 27353 25927 27387
rect 26896 27384 26924 27415
rect 28350 27412 28356 27424
rect 28408 27412 28414 27464
rect 25869 27347 25927 27353
rect 26252 27356 26924 27384
rect 8113 27319 8171 27325
rect 8113 27285 8125 27319
rect 8159 27316 8171 27319
rect 8754 27316 8760 27328
rect 8159 27288 8760 27316
rect 8159 27285 8171 27288
rect 8113 27279 8171 27285
rect 8754 27276 8760 27288
rect 8812 27276 8818 27328
rect 11054 27276 11060 27328
rect 11112 27316 11118 27328
rect 11606 27316 11612 27328
rect 11112 27288 11612 27316
rect 11112 27276 11118 27288
rect 11606 27276 11612 27288
rect 11664 27316 11670 27328
rect 12069 27319 12127 27325
rect 12069 27316 12081 27319
rect 11664 27288 12081 27316
rect 11664 27276 11670 27288
rect 12069 27285 12081 27288
rect 12115 27285 12127 27319
rect 12069 27279 12127 27285
rect 14090 27276 14096 27328
rect 14148 27316 14154 27328
rect 14369 27319 14427 27325
rect 14369 27316 14381 27319
rect 14148 27288 14381 27316
rect 14148 27276 14154 27288
rect 14369 27285 14381 27288
rect 14415 27285 14427 27319
rect 14369 27279 14427 27285
rect 14826 27276 14832 27328
rect 14884 27316 14890 27328
rect 14921 27319 14979 27325
rect 14921 27316 14933 27319
rect 14884 27288 14933 27316
rect 14884 27276 14890 27288
rect 14921 27285 14933 27288
rect 14967 27285 14979 27319
rect 14921 27279 14979 27285
rect 16025 27319 16083 27325
rect 16025 27285 16037 27319
rect 16071 27316 16083 27319
rect 16390 27316 16396 27328
rect 16071 27288 16396 27316
rect 16071 27285 16083 27288
rect 16025 27279 16083 27285
rect 16390 27276 16396 27288
rect 16448 27276 16454 27328
rect 17865 27319 17923 27325
rect 17865 27285 17877 27319
rect 17911 27316 17923 27319
rect 17954 27316 17960 27328
rect 17911 27288 17960 27316
rect 17911 27285 17923 27288
rect 17865 27279 17923 27285
rect 17954 27276 17960 27288
rect 18012 27276 18018 27328
rect 24946 27316 24952 27328
rect 24907 27288 24952 27316
rect 24946 27276 24952 27288
rect 25004 27276 25010 27328
rect 26252 27325 26280 27356
rect 26237 27319 26295 27325
rect 26237 27285 26249 27319
rect 26283 27285 26295 27319
rect 27062 27316 27068 27328
rect 27023 27288 27068 27316
rect 26237 27279 26295 27285
rect 27062 27276 27068 27288
rect 27120 27276 27126 27328
rect 27522 27316 27528 27328
rect 27483 27288 27528 27316
rect 27522 27276 27528 27288
rect 27580 27276 27586 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 8018 27112 8024 27124
rect 7979 27084 8024 27112
rect 8018 27072 8024 27084
rect 8076 27072 8082 27124
rect 9125 27115 9183 27121
rect 9125 27081 9137 27115
rect 9171 27112 9183 27115
rect 9214 27112 9220 27124
rect 9171 27084 9220 27112
rect 9171 27081 9183 27084
rect 9125 27075 9183 27081
rect 9214 27072 9220 27084
rect 9272 27072 9278 27124
rect 9858 27112 9864 27124
rect 9819 27084 9864 27112
rect 9858 27072 9864 27084
rect 9916 27072 9922 27124
rect 10965 27115 11023 27121
rect 10965 27081 10977 27115
rect 11011 27112 11023 27115
rect 11238 27112 11244 27124
rect 11011 27084 11244 27112
rect 11011 27081 11023 27084
rect 10965 27075 11023 27081
rect 11238 27072 11244 27084
rect 11296 27072 11302 27124
rect 13078 27072 13084 27124
rect 13136 27112 13142 27124
rect 13449 27115 13507 27121
rect 13449 27112 13461 27115
rect 13136 27084 13461 27112
rect 13136 27072 13142 27084
rect 13449 27081 13461 27084
rect 13495 27081 13507 27115
rect 13449 27075 13507 27081
rect 13633 27115 13691 27121
rect 13633 27081 13645 27115
rect 13679 27081 13691 27115
rect 13633 27075 13691 27081
rect 8938 27004 8944 27056
rect 8996 27044 9002 27056
rect 8996 27016 12756 27044
rect 8996 27004 9002 27016
rect 7745 26979 7803 26985
rect 7745 26945 7757 26979
rect 7791 26976 7803 26979
rect 8386 26976 8392 26988
rect 7791 26948 8392 26976
rect 7791 26945 7803 26948
rect 7745 26939 7803 26945
rect 8386 26936 8392 26948
rect 8444 26936 8450 26988
rect 8754 26936 8760 26988
rect 8812 26976 8818 26988
rect 8849 26979 8907 26985
rect 8849 26976 8861 26979
rect 8812 26948 8861 26976
rect 8812 26936 8818 26948
rect 8849 26945 8861 26948
rect 8895 26945 8907 26979
rect 8849 26939 8907 26945
rect 9585 26979 9643 26985
rect 9585 26945 9597 26979
rect 9631 26976 9643 26979
rect 9766 26976 9772 26988
rect 9631 26948 9772 26976
rect 9631 26945 9643 26948
rect 9585 26939 9643 26945
rect 9766 26936 9772 26948
rect 9824 26936 9830 26988
rect 8021 26911 8079 26917
rect 8021 26877 8033 26911
rect 8067 26908 8079 26911
rect 8294 26908 8300 26920
rect 8067 26880 8300 26908
rect 8067 26877 8079 26880
rect 8021 26871 8079 26877
rect 8294 26868 8300 26880
rect 8352 26868 8358 26920
rect 8481 26911 8539 26917
rect 8481 26877 8493 26911
rect 8527 26877 8539 26911
rect 8481 26871 8539 26877
rect 8496 26840 8524 26871
rect 8570 26868 8576 26920
rect 8628 26908 8634 26920
rect 8938 26908 8944 26920
rect 8628 26880 8944 26908
rect 8628 26868 8634 26880
rect 8938 26868 8944 26880
rect 8996 26868 9002 26920
rect 9876 26917 9904 27016
rect 10594 26936 10600 26988
rect 10652 26976 10658 26988
rect 11517 26979 11575 26985
rect 11517 26976 11529 26979
rect 10652 26948 11529 26976
rect 10652 26936 10658 26948
rect 11517 26945 11529 26948
rect 11563 26945 11575 26979
rect 11517 26939 11575 26945
rect 12437 26979 12495 26985
rect 12437 26945 12449 26979
rect 12483 26945 12495 26979
rect 12437 26939 12495 26945
rect 9861 26911 9919 26917
rect 9861 26877 9873 26911
rect 9907 26877 9919 26911
rect 9861 26871 9919 26877
rect 10321 26911 10379 26917
rect 10321 26877 10333 26911
rect 10367 26877 10379 26911
rect 10686 26908 10692 26920
rect 10647 26880 10692 26908
rect 10321 26871 10379 26877
rect 8846 26840 8852 26852
rect 8496 26812 8852 26840
rect 8846 26800 8852 26812
rect 8904 26800 8910 26852
rect 9677 26843 9735 26849
rect 9677 26809 9689 26843
rect 9723 26840 9735 26843
rect 10336 26840 10364 26871
rect 10686 26868 10692 26880
rect 10744 26868 10750 26920
rect 10781 26911 10839 26917
rect 10781 26877 10793 26911
rect 10827 26908 10839 26911
rect 11146 26908 11152 26920
rect 10827 26880 11152 26908
rect 10827 26877 10839 26880
rect 10781 26871 10839 26877
rect 11146 26868 11152 26880
rect 11204 26868 11210 26920
rect 12158 26908 12164 26920
rect 12119 26880 12164 26908
rect 12158 26868 12164 26880
rect 12216 26868 12222 26920
rect 12452 26840 12480 26939
rect 12728 26908 12756 27016
rect 12802 27004 12808 27056
rect 12860 27044 12866 27056
rect 13648 27044 13676 27075
rect 14458 27072 14464 27124
rect 14516 27112 14522 27124
rect 14645 27115 14703 27121
rect 14645 27112 14657 27115
rect 14516 27084 14657 27112
rect 14516 27072 14522 27084
rect 14645 27081 14657 27084
rect 14691 27081 14703 27115
rect 15194 27112 15200 27124
rect 14645 27075 14703 27081
rect 14752 27084 15200 27112
rect 12860 27016 13676 27044
rect 12860 27004 12866 27016
rect 13262 26936 13268 26988
rect 13320 26976 13326 26988
rect 13574 26979 13632 26985
rect 13574 26976 13586 26979
rect 13320 26948 13586 26976
rect 13320 26936 13326 26948
rect 13574 26945 13586 26948
rect 13620 26945 13632 26979
rect 14090 26976 14096 26988
rect 14051 26948 14096 26976
rect 13574 26939 13632 26945
rect 14090 26936 14096 26948
rect 14148 26936 14154 26988
rect 14752 26908 14780 27084
rect 15194 27072 15200 27084
rect 15252 27072 15258 27124
rect 15838 27072 15844 27124
rect 15896 27112 15902 27124
rect 16025 27115 16083 27121
rect 16025 27112 16037 27115
rect 15896 27084 16037 27112
rect 15896 27072 15902 27084
rect 16025 27081 16037 27084
rect 16071 27081 16083 27115
rect 16025 27075 16083 27081
rect 17497 27115 17555 27121
rect 17497 27081 17509 27115
rect 17543 27112 17555 27115
rect 18598 27112 18604 27124
rect 17543 27084 18604 27112
rect 17543 27081 17555 27084
rect 17497 27075 17555 27081
rect 18598 27072 18604 27084
rect 18656 27072 18662 27124
rect 20070 27112 20076 27124
rect 20031 27084 20076 27112
rect 20070 27072 20076 27084
rect 20128 27072 20134 27124
rect 20533 27115 20591 27121
rect 20533 27081 20545 27115
rect 20579 27112 20591 27115
rect 22186 27112 22192 27124
rect 20579 27084 22192 27112
rect 20579 27081 20591 27084
rect 20533 27075 20591 27081
rect 22186 27072 22192 27084
rect 22244 27072 22250 27124
rect 22738 27072 22744 27124
rect 22796 27112 22802 27124
rect 25498 27112 25504 27124
rect 22796 27084 22876 27112
rect 25459 27084 25504 27112
rect 22796 27072 22802 27084
rect 15010 27044 15016 27056
rect 14844 27016 15016 27044
rect 14844 26985 14872 27016
rect 15010 27004 15016 27016
rect 15068 27004 15074 27056
rect 16853 27047 16911 27053
rect 15948 27016 16804 27044
rect 14829 26979 14887 26985
rect 14829 26945 14841 26979
rect 14875 26945 14887 26979
rect 14829 26939 14887 26945
rect 14918 26936 14924 26988
rect 14976 26976 14982 26988
rect 14976 26948 15021 26976
rect 15102 26960 15108 27012
rect 15160 26960 15166 27012
rect 15948 26988 15976 27016
rect 14976 26936 14982 26948
rect 15105 26945 15117 26960
rect 15151 26945 15163 26960
rect 15105 26939 15163 26945
rect 15194 26936 15200 26988
rect 15252 26976 15258 26988
rect 15289 26979 15347 26985
rect 15289 26976 15301 26979
rect 15252 26948 15301 26976
rect 15252 26936 15258 26948
rect 15289 26945 15301 26948
rect 15335 26976 15347 26979
rect 15470 26976 15476 26988
rect 15335 26948 15476 26976
rect 15335 26945 15347 26948
rect 15289 26939 15347 26945
rect 15470 26936 15476 26948
rect 15528 26936 15534 26988
rect 15930 26976 15936 26988
rect 15891 26948 15936 26976
rect 15930 26936 15936 26948
rect 15988 26936 15994 26988
rect 16117 26979 16175 26985
rect 16117 26945 16129 26979
rect 16163 26976 16175 26979
rect 16206 26976 16212 26988
rect 16163 26948 16212 26976
rect 16163 26945 16175 26948
rect 16117 26939 16175 26945
rect 16206 26936 16212 26948
rect 16264 26936 16270 26988
rect 16776 26976 16804 27016
rect 16853 27013 16865 27047
rect 16899 27044 16911 27047
rect 17954 27044 17960 27056
rect 16899 27016 17960 27044
rect 16899 27013 16911 27016
rect 16853 27007 16911 27013
rect 17954 27004 17960 27016
rect 18012 27004 18018 27056
rect 18616 27044 18644 27072
rect 18616 27016 19012 27044
rect 17218 26976 17224 26988
rect 16776 26948 17224 26976
rect 17218 26936 17224 26948
rect 17276 26936 17282 26988
rect 17862 26976 17868 26988
rect 17823 26948 17868 26976
rect 17862 26936 17868 26948
rect 17920 26936 17926 26988
rect 18877 26979 18935 26985
rect 18877 26976 18889 26979
rect 18064 26948 18889 26976
rect 12728 26880 14780 26908
rect 15013 26911 15071 26917
rect 15013 26877 15025 26911
rect 15059 26908 15071 26911
rect 15562 26908 15568 26920
rect 15059 26880 15568 26908
rect 15059 26877 15071 26880
rect 15013 26871 15071 26877
rect 15562 26868 15568 26880
rect 15620 26868 15626 26920
rect 16022 26868 16028 26920
rect 16080 26908 16086 26920
rect 17957 26911 18015 26917
rect 17957 26908 17969 26911
rect 16080 26880 17969 26908
rect 16080 26868 16086 26880
rect 17957 26877 17969 26880
rect 18003 26877 18015 26911
rect 17957 26871 18015 26877
rect 13262 26840 13268 26852
rect 9723 26812 13268 26840
rect 9723 26809 9735 26812
rect 9677 26803 9735 26809
rect 13262 26800 13268 26812
rect 13320 26800 13326 26852
rect 14001 26843 14059 26849
rect 14001 26809 14013 26843
rect 14047 26809 14059 26843
rect 14001 26803 14059 26809
rect 7837 26775 7895 26781
rect 7837 26741 7849 26775
rect 7883 26772 7895 26775
rect 8018 26772 8024 26784
rect 7883 26744 8024 26772
rect 7883 26741 7895 26744
rect 7837 26735 7895 26741
rect 8018 26732 8024 26744
rect 8076 26732 8082 26784
rect 10410 26732 10416 26784
rect 10468 26772 10474 26784
rect 11609 26775 11667 26781
rect 11609 26772 11621 26775
rect 10468 26744 11621 26772
rect 10468 26732 10474 26744
rect 11609 26741 11621 26744
rect 11655 26741 11667 26775
rect 14016 26772 14044 26803
rect 15194 26800 15200 26852
rect 15252 26840 15258 26852
rect 16482 26840 16488 26852
rect 15252 26812 16488 26840
rect 15252 26800 15258 26812
rect 16482 26800 16488 26812
rect 16540 26800 16546 26852
rect 16850 26800 16856 26852
rect 16908 26840 16914 26852
rect 17037 26843 17095 26849
rect 17037 26840 17049 26843
rect 16908 26812 17049 26840
rect 16908 26800 16914 26812
rect 17037 26809 17049 26812
rect 17083 26840 17095 26843
rect 18064 26840 18092 26948
rect 18877 26945 18889 26948
rect 18923 26945 18935 26979
rect 18984 26976 19012 27016
rect 19334 27004 19340 27056
rect 19392 27044 19398 27056
rect 22848 27053 22876 27084
rect 25498 27072 25504 27084
rect 25556 27072 25562 27124
rect 25774 27072 25780 27124
rect 25832 27112 25838 27124
rect 25869 27115 25927 27121
rect 25869 27112 25881 27115
rect 25832 27084 25881 27112
rect 25832 27072 25838 27084
rect 25869 27081 25881 27084
rect 25915 27081 25927 27115
rect 25869 27075 25927 27081
rect 25961 27115 26019 27121
rect 25961 27081 25973 27115
rect 26007 27112 26019 27115
rect 26050 27112 26056 27124
rect 26007 27084 26056 27112
rect 26007 27081 26019 27084
rect 25961 27075 26019 27081
rect 26050 27072 26056 27084
rect 26108 27072 26114 27124
rect 28350 27112 28356 27124
rect 28311 27084 28356 27112
rect 28350 27072 28356 27084
rect 28408 27072 28414 27124
rect 19889 27047 19947 27053
rect 19889 27044 19901 27047
rect 19392 27016 19901 27044
rect 19392 27004 19398 27016
rect 19889 27013 19901 27016
rect 19935 27013 19947 27047
rect 19889 27007 19947 27013
rect 22833 27047 22891 27053
rect 22833 27013 22845 27047
rect 22879 27013 22891 27047
rect 26878 27044 26884 27056
rect 22833 27007 22891 27013
rect 23676 27016 26884 27044
rect 19705 26979 19763 26985
rect 19705 26976 19717 26979
rect 18984 26948 19717 26976
rect 18877 26939 18935 26945
rect 19705 26945 19717 26948
rect 19751 26945 19763 26979
rect 19705 26939 19763 26945
rect 18141 26911 18199 26917
rect 18141 26877 18153 26911
rect 18187 26908 18199 26911
rect 18785 26911 18843 26917
rect 18785 26908 18797 26911
rect 18187 26880 18797 26908
rect 18187 26877 18199 26880
rect 18141 26871 18199 26877
rect 18785 26877 18797 26880
rect 18831 26877 18843 26911
rect 18892 26908 18920 26939
rect 19978 26936 19984 26988
rect 20036 26976 20042 26988
rect 20717 26979 20775 26985
rect 20717 26976 20729 26979
rect 20036 26948 20729 26976
rect 20036 26936 20042 26948
rect 20717 26945 20729 26948
rect 20763 26945 20775 26979
rect 20717 26939 20775 26945
rect 21913 26979 21971 26985
rect 21913 26945 21925 26979
rect 21959 26976 21971 26979
rect 22738 26976 22744 26988
rect 21959 26948 22744 26976
rect 21959 26945 21971 26948
rect 21913 26939 21971 26945
rect 22738 26936 22744 26948
rect 22796 26976 22802 26988
rect 22922 26976 22928 26988
rect 22796 26948 22928 26976
rect 22796 26936 22802 26948
rect 22922 26936 22928 26948
rect 22980 26936 22986 26988
rect 23106 26936 23112 26988
rect 23164 26976 23170 26988
rect 23676 26985 23704 27016
rect 26878 27004 26884 27016
rect 26936 27004 26942 27056
rect 27249 27047 27307 27053
rect 27249 27013 27261 27047
rect 27295 27044 27307 27047
rect 28442 27044 28448 27056
rect 27295 27016 28448 27044
rect 27295 27013 27307 27016
rect 27249 27007 27307 27013
rect 28442 27004 28448 27016
rect 28500 27004 28506 27056
rect 23661 26979 23719 26985
rect 23164 26948 23244 26976
rect 23164 26936 23170 26948
rect 18966 26908 18972 26920
rect 18892 26880 18972 26908
rect 18785 26871 18843 26877
rect 17083 26812 18092 26840
rect 17083 26809 17095 26812
rect 17037 26803 17095 26809
rect 14274 26772 14280 26784
rect 14016 26744 14280 26772
rect 11609 26735 11667 26741
rect 14274 26732 14280 26744
rect 14332 26772 14338 26784
rect 14918 26772 14924 26784
rect 14332 26744 14924 26772
rect 14332 26732 14338 26744
rect 14918 26732 14924 26744
rect 14976 26772 14982 26784
rect 16942 26772 16948 26784
rect 14976 26744 16948 26772
rect 14976 26732 14982 26744
rect 16942 26732 16948 26744
rect 17000 26732 17006 26784
rect 18800 26772 18828 26871
rect 18966 26868 18972 26880
rect 19024 26868 19030 26920
rect 22002 26908 22008 26920
rect 21963 26880 22008 26908
rect 22002 26868 22008 26880
rect 22060 26868 22066 26920
rect 19245 26843 19303 26849
rect 19245 26809 19257 26843
rect 19291 26840 19303 26843
rect 19426 26840 19432 26852
rect 19291 26812 19432 26840
rect 19291 26809 19303 26812
rect 19245 26803 19303 26809
rect 19426 26800 19432 26812
rect 19484 26800 19490 26852
rect 20622 26800 20628 26852
rect 20680 26840 20686 26852
rect 23106 26840 23112 26852
rect 20680 26812 23112 26840
rect 20680 26800 20686 26812
rect 23106 26800 23112 26812
rect 23164 26800 23170 26852
rect 19518 26772 19524 26784
rect 18800 26744 19524 26772
rect 19518 26732 19524 26744
rect 19576 26772 19582 26784
rect 19978 26772 19984 26784
rect 19576 26744 19984 26772
rect 19576 26732 19582 26744
rect 19978 26732 19984 26744
rect 20036 26732 20042 26784
rect 22094 26732 22100 26784
rect 22152 26772 22158 26784
rect 22281 26775 22339 26781
rect 22152 26744 22197 26772
rect 22152 26732 22158 26744
rect 22281 26741 22293 26775
rect 22327 26772 22339 26775
rect 22554 26772 22560 26784
rect 22327 26744 22560 26772
rect 22327 26741 22339 26744
rect 22281 26735 22339 26741
rect 22554 26732 22560 26744
rect 22612 26732 22618 26784
rect 22922 26772 22928 26784
rect 22883 26744 22928 26772
rect 22922 26732 22928 26744
rect 22980 26772 22986 26784
rect 23216 26772 23244 26948
rect 23661 26945 23673 26979
rect 23707 26945 23719 26979
rect 23661 26939 23719 26945
rect 23928 26979 23986 26985
rect 23928 26945 23940 26979
rect 23974 26976 23986 26979
rect 25774 26976 25780 26988
rect 23974 26948 25780 26976
rect 23974 26945 23986 26948
rect 23928 26939 23986 26945
rect 25774 26936 25780 26948
rect 25832 26936 25838 26988
rect 26973 26979 27031 26985
rect 26973 26976 26985 26979
rect 25976 26948 26985 26976
rect 25682 26868 25688 26920
rect 25740 26908 25746 26920
rect 25976 26908 26004 26948
rect 26973 26945 26985 26948
rect 27019 26945 27031 26979
rect 27154 26976 27160 26988
rect 27115 26948 27160 26976
rect 26973 26939 27031 26945
rect 27154 26936 27160 26948
rect 27212 26936 27218 26988
rect 27341 26979 27399 26985
rect 27341 26945 27353 26979
rect 27387 26945 27399 26979
rect 28169 26979 28227 26985
rect 28169 26976 28181 26979
rect 27341 26939 27399 26945
rect 27540 26948 28181 26976
rect 25740 26880 26004 26908
rect 26053 26911 26111 26917
rect 25740 26868 25746 26880
rect 26053 26877 26065 26911
rect 26099 26877 26111 26911
rect 26053 26871 26111 26877
rect 24670 26800 24676 26852
rect 24728 26840 24734 26852
rect 26068 26840 26096 26871
rect 26142 26868 26148 26920
rect 26200 26908 26206 26920
rect 27356 26908 27384 26939
rect 26200 26880 27384 26908
rect 26200 26868 26206 26880
rect 27540 26849 27568 26948
rect 28169 26945 28181 26948
rect 28215 26945 28227 26979
rect 28169 26939 28227 26945
rect 27985 26911 28043 26917
rect 27985 26908 27997 26911
rect 27632 26880 27997 26908
rect 24728 26812 26096 26840
rect 27525 26843 27583 26849
rect 24728 26800 24734 26812
rect 27525 26809 27537 26843
rect 27571 26809 27583 26843
rect 27525 26803 27583 26809
rect 22980 26744 23244 26772
rect 25041 26775 25099 26781
rect 22980 26732 22986 26744
rect 25041 26741 25053 26775
rect 25087 26772 25099 26775
rect 25222 26772 25228 26784
rect 25087 26744 25228 26772
rect 25087 26741 25099 26744
rect 25041 26735 25099 26741
rect 25222 26732 25228 26744
rect 25280 26732 25286 26784
rect 26970 26732 26976 26784
rect 27028 26772 27034 26784
rect 27632 26772 27660 26880
rect 27985 26877 27997 26880
rect 28031 26877 28043 26911
rect 27985 26871 28043 26877
rect 27028 26744 27660 26772
rect 27028 26732 27034 26744
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 8018 26568 8024 26580
rect 7979 26540 8024 26568
rect 8018 26528 8024 26540
rect 8076 26528 8082 26580
rect 8389 26571 8447 26577
rect 8389 26537 8401 26571
rect 8435 26568 8447 26571
rect 8754 26568 8760 26580
rect 8435 26540 8760 26568
rect 8435 26537 8447 26540
rect 8389 26531 8447 26537
rect 8754 26528 8760 26540
rect 8812 26528 8818 26580
rect 8941 26571 8999 26577
rect 8941 26537 8953 26571
rect 8987 26537 8999 26571
rect 8941 26531 8999 26537
rect 9401 26571 9459 26577
rect 9401 26537 9413 26571
rect 9447 26568 9459 26571
rect 10686 26568 10692 26580
rect 9447 26540 10692 26568
rect 9447 26537 9459 26540
rect 9401 26531 9459 26537
rect 8036 26500 8064 26528
rect 8662 26500 8668 26512
rect 8036 26472 8668 26500
rect 8662 26460 8668 26472
rect 8720 26500 8726 26512
rect 8956 26500 8984 26531
rect 10686 26528 10692 26540
rect 10744 26528 10750 26580
rect 11146 26568 11152 26580
rect 11107 26540 11152 26568
rect 11146 26528 11152 26540
rect 11204 26528 11210 26580
rect 11974 26528 11980 26580
rect 12032 26568 12038 26580
rect 12069 26571 12127 26577
rect 12069 26568 12081 26571
rect 12032 26540 12081 26568
rect 12032 26528 12038 26540
rect 12069 26537 12081 26540
rect 12115 26537 12127 26571
rect 12069 26531 12127 26537
rect 14829 26571 14887 26577
rect 14829 26537 14841 26571
rect 14875 26568 14887 26571
rect 15838 26568 15844 26580
rect 14875 26540 15844 26568
rect 14875 26537 14887 26540
rect 14829 26531 14887 26537
rect 15838 26528 15844 26540
rect 15896 26528 15902 26580
rect 17037 26571 17095 26577
rect 17037 26537 17049 26571
rect 17083 26537 17095 26571
rect 17037 26531 17095 26537
rect 8720 26472 8984 26500
rect 8720 26460 8726 26472
rect 9030 26460 9036 26512
rect 9088 26500 9094 26512
rect 9953 26503 10011 26509
rect 9953 26500 9965 26503
rect 9088 26472 9965 26500
rect 9088 26460 9094 26472
rect 9953 26469 9965 26472
rect 9999 26469 10011 26503
rect 11330 26500 11336 26512
rect 9953 26463 10011 26469
rect 10244 26472 11336 26500
rect 8294 26432 8300 26444
rect 8036 26404 8300 26432
rect 8036 26373 8064 26404
rect 8294 26392 8300 26404
rect 8352 26432 8358 26444
rect 8352 26404 9168 26432
rect 8352 26392 8358 26404
rect 9140 26376 9168 26404
rect 9306 26392 9312 26444
rect 9364 26432 9370 26444
rect 10244 26432 10272 26472
rect 11330 26460 11336 26472
rect 11388 26500 11394 26512
rect 11388 26472 12572 26500
rect 11388 26460 11394 26472
rect 10410 26432 10416 26444
rect 9364 26404 10272 26432
rect 10371 26404 10416 26432
rect 9364 26392 9370 26404
rect 10410 26392 10416 26404
rect 10468 26392 10474 26444
rect 10597 26435 10655 26441
rect 10597 26401 10609 26435
rect 10643 26432 10655 26435
rect 10778 26432 10784 26444
rect 10643 26404 10784 26432
rect 10643 26401 10655 26404
rect 10597 26395 10655 26401
rect 10778 26392 10784 26404
rect 10836 26392 10842 26444
rect 12544 26432 12572 26472
rect 14090 26460 14096 26512
rect 14148 26500 14154 26512
rect 14369 26503 14427 26509
rect 14369 26500 14381 26503
rect 14148 26472 14381 26500
rect 14148 26460 14154 26472
rect 14369 26469 14381 26472
rect 14415 26500 14427 26503
rect 14642 26500 14648 26512
rect 14415 26472 14648 26500
rect 14415 26469 14427 26472
rect 14369 26463 14427 26469
rect 14642 26460 14648 26472
rect 14700 26500 14706 26512
rect 15194 26500 15200 26512
rect 14700 26472 15200 26500
rect 14700 26460 14706 26472
rect 15194 26460 15200 26472
rect 15252 26460 15258 26512
rect 17052 26500 17080 26531
rect 17402 26528 17408 26580
rect 17460 26568 17466 26580
rect 17862 26568 17868 26580
rect 17460 26540 17868 26568
rect 17460 26528 17466 26540
rect 17862 26528 17868 26540
rect 17920 26568 17926 26580
rect 18141 26571 18199 26577
rect 18141 26568 18153 26571
rect 17920 26540 18153 26568
rect 17920 26528 17926 26540
rect 18141 26537 18153 26540
rect 18187 26537 18199 26571
rect 19334 26568 19340 26580
rect 19295 26540 19340 26568
rect 18141 26531 18199 26537
rect 19334 26528 19340 26540
rect 19392 26528 19398 26580
rect 20165 26571 20223 26577
rect 20165 26537 20177 26571
rect 20211 26568 20223 26571
rect 20254 26568 20260 26580
rect 20211 26540 20260 26568
rect 20211 26537 20223 26540
rect 20165 26531 20223 26537
rect 20254 26528 20260 26540
rect 20312 26528 20318 26580
rect 20806 26568 20812 26580
rect 20767 26540 20812 26568
rect 20806 26528 20812 26540
rect 20864 26528 20870 26580
rect 20898 26528 20904 26580
rect 20956 26568 20962 26580
rect 21177 26571 21235 26577
rect 21177 26568 21189 26571
rect 20956 26540 21189 26568
rect 20956 26528 20962 26540
rect 21177 26537 21189 26540
rect 21223 26537 21235 26571
rect 21177 26531 21235 26537
rect 22649 26571 22707 26577
rect 22649 26537 22661 26571
rect 22695 26568 22707 26571
rect 22830 26568 22836 26580
rect 22695 26540 22836 26568
rect 22695 26537 22707 26540
rect 22649 26531 22707 26537
rect 22830 26528 22836 26540
rect 22888 26528 22894 26580
rect 25501 26571 25559 26577
rect 25501 26537 25513 26571
rect 25547 26568 25559 26571
rect 27154 26568 27160 26580
rect 25547 26540 27160 26568
rect 25547 26537 25559 26540
rect 25501 26531 25559 26537
rect 27154 26528 27160 26540
rect 27212 26528 27218 26580
rect 16776 26472 17080 26500
rect 13449 26435 13507 26441
rect 13449 26432 13461 26435
rect 12544 26404 13461 26432
rect 8021 26367 8079 26373
rect 8021 26333 8033 26367
rect 8067 26333 8079 26367
rect 8021 26327 8079 26333
rect 8205 26367 8263 26373
rect 8205 26333 8217 26367
rect 8251 26333 8263 26367
rect 8938 26364 8944 26376
rect 8899 26336 8944 26364
rect 8205 26327 8263 26333
rect 8220 26296 8248 26327
rect 8938 26324 8944 26336
rect 8996 26324 9002 26376
rect 9122 26364 9128 26376
rect 9083 26336 9128 26364
rect 9122 26324 9128 26336
rect 9180 26324 9186 26376
rect 9217 26367 9275 26373
rect 9217 26333 9229 26367
rect 9263 26333 9275 26367
rect 10318 26364 10324 26376
rect 10279 26336 10324 26364
rect 9217 26327 9275 26333
rect 8294 26296 8300 26308
rect 8220 26268 8300 26296
rect 8294 26256 8300 26268
rect 8352 26296 8358 26308
rect 9232 26296 9260 26327
rect 10318 26324 10324 26336
rect 10376 26324 10382 26376
rect 11330 26364 11336 26376
rect 11291 26336 11336 26364
rect 11330 26324 11336 26336
rect 11388 26324 11394 26376
rect 11514 26364 11520 26376
rect 11475 26336 11520 26364
rect 11514 26324 11520 26336
rect 11572 26324 11578 26376
rect 11606 26324 11612 26376
rect 11664 26364 11670 26376
rect 12253 26367 12311 26373
rect 11664 26336 11709 26364
rect 11664 26324 11670 26336
rect 12253 26333 12265 26367
rect 12299 26364 12311 26367
rect 12434 26364 12440 26376
rect 12299 26336 12440 26364
rect 12299 26333 12311 26336
rect 12253 26327 12311 26333
rect 12434 26324 12440 26336
rect 12492 26324 12498 26376
rect 12544 26373 12572 26404
rect 13449 26401 13461 26404
rect 13495 26401 13507 26435
rect 13449 26395 13507 26401
rect 14918 26392 14924 26444
rect 14976 26432 14982 26444
rect 14976 26404 15240 26432
rect 14976 26392 14982 26404
rect 12529 26367 12587 26373
rect 12529 26333 12541 26367
rect 12575 26333 12587 26367
rect 12529 26327 12587 26333
rect 12713 26367 12771 26373
rect 12713 26333 12725 26367
rect 12759 26364 12771 26367
rect 12986 26364 12992 26376
rect 12759 26336 12992 26364
rect 12759 26333 12771 26336
rect 12713 26327 12771 26333
rect 12986 26324 12992 26336
rect 13044 26324 13050 26376
rect 13262 26364 13268 26376
rect 13223 26336 13268 26364
rect 13262 26324 13268 26336
rect 13320 26324 13326 26376
rect 14642 26324 14648 26376
rect 14700 26364 14706 26376
rect 15013 26367 15071 26373
rect 15013 26364 15025 26367
rect 14700 26336 15025 26364
rect 14700 26324 14706 26336
rect 15013 26333 15025 26336
rect 15059 26333 15071 26367
rect 15013 26327 15071 26333
rect 15105 26367 15163 26373
rect 15105 26333 15117 26367
rect 15151 26361 15163 26367
rect 15212 26361 15240 26404
rect 15286 26392 15292 26444
rect 15344 26432 15350 26444
rect 15473 26435 15531 26441
rect 15473 26432 15485 26435
rect 15344 26404 15485 26432
rect 15344 26392 15350 26404
rect 15473 26401 15485 26404
rect 15519 26401 15531 26435
rect 16776 26432 16804 26472
rect 22094 26460 22100 26512
rect 22152 26500 22158 26512
rect 23014 26500 23020 26512
rect 22152 26472 23020 26500
rect 22152 26460 22158 26472
rect 23014 26460 23020 26472
rect 23072 26500 23078 26512
rect 23293 26503 23351 26509
rect 23293 26500 23305 26503
rect 23072 26472 23305 26500
rect 23072 26460 23078 26472
rect 23293 26469 23305 26472
rect 23339 26469 23351 26503
rect 23293 26463 23351 26469
rect 28166 26460 28172 26512
rect 28224 26500 28230 26512
rect 28261 26503 28319 26509
rect 28261 26500 28273 26503
rect 28224 26472 28273 26500
rect 28224 26460 28230 26472
rect 28261 26469 28273 26472
rect 28307 26469 28319 26503
rect 28261 26463 28319 26469
rect 15473 26395 15531 26401
rect 16316 26404 16804 26432
rect 15151 26333 15240 26361
rect 15381 26367 15439 26373
rect 15381 26333 15393 26367
rect 15427 26364 15439 26367
rect 15838 26364 15844 26376
rect 15427 26336 15844 26364
rect 15427 26333 15439 26336
rect 15105 26327 15163 26333
rect 15381 26327 15439 26333
rect 15838 26324 15844 26336
rect 15896 26324 15902 26376
rect 16114 26364 16120 26376
rect 16040 26336 16120 26364
rect 8352 26268 9260 26296
rect 14185 26299 14243 26305
rect 8352 26256 8358 26268
rect 14185 26265 14197 26299
rect 14231 26296 14243 26299
rect 15286 26296 15292 26308
rect 14231 26268 15292 26296
rect 14231 26265 14243 26268
rect 14185 26259 14243 26265
rect 15286 26256 15292 26268
rect 15344 26256 15350 26308
rect 7742 26188 7748 26240
rect 7800 26228 7806 26240
rect 12342 26228 12348 26240
rect 7800 26200 12348 26228
rect 7800 26188 7806 26200
rect 12342 26188 12348 26200
rect 12400 26188 12406 26240
rect 12526 26188 12532 26240
rect 12584 26228 12590 26240
rect 13722 26228 13728 26240
rect 12584 26200 13728 26228
rect 12584 26188 12590 26200
rect 13722 26188 13728 26200
rect 13780 26188 13786 26240
rect 15933 26231 15991 26237
rect 15933 26197 15945 26231
rect 15979 26228 15991 26231
rect 16040 26228 16068 26336
rect 16114 26324 16120 26336
rect 16172 26324 16178 26376
rect 16316 26373 16344 26404
rect 16942 26392 16948 26444
rect 17000 26432 17006 26444
rect 17497 26435 17555 26441
rect 17497 26432 17509 26435
rect 17000 26404 17509 26432
rect 17000 26392 17006 26404
rect 17497 26401 17509 26404
rect 17543 26401 17555 26435
rect 20990 26432 20996 26444
rect 17497 26395 17555 26401
rect 20824 26404 20996 26432
rect 16209 26367 16267 26373
rect 16209 26333 16221 26367
rect 16255 26333 16267 26367
rect 16209 26327 16267 26333
rect 16301 26367 16359 26373
rect 16301 26333 16313 26367
rect 16347 26333 16359 26367
rect 16301 26327 16359 26333
rect 16224 26296 16252 26327
rect 16390 26324 16396 26376
rect 16448 26364 16454 26376
rect 16577 26367 16635 26373
rect 16448 26336 16493 26364
rect 16448 26324 16454 26336
rect 16577 26333 16589 26367
rect 16623 26364 16635 26367
rect 16666 26364 16672 26376
rect 16623 26336 16672 26364
rect 16623 26333 16635 26336
rect 16577 26327 16635 26333
rect 16666 26324 16672 26336
rect 16724 26324 16730 26376
rect 17218 26364 17224 26376
rect 17179 26336 17224 26364
rect 17218 26324 17224 26336
rect 17276 26324 17282 26376
rect 17405 26367 17463 26373
rect 17405 26333 17417 26367
rect 17451 26333 17463 26367
rect 19242 26364 19248 26376
rect 19203 26336 19248 26364
rect 17405 26327 17463 26333
rect 16850 26296 16856 26308
rect 16224 26268 16856 26296
rect 16850 26256 16856 26268
rect 16908 26256 16914 26308
rect 17034 26256 17040 26308
rect 17092 26296 17098 26308
rect 17420 26296 17448 26327
rect 19242 26324 19248 26336
rect 19300 26324 19306 26376
rect 19334 26324 19340 26376
rect 19392 26364 19398 26376
rect 19429 26367 19487 26373
rect 19429 26364 19441 26367
rect 19392 26336 19441 26364
rect 19392 26324 19398 26336
rect 19429 26333 19441 26336
rect 19475 26333 19487 26367
rect 19429 26327 19487 26333
rect 20349 26367 20407 26373
rect 20349 26333 20361 26367
rect 20395 26364 20407 26367
rect 20714 26364 20720 26376
rect 20395 26336 20720 26364
rect 20395 26333 20407 26336
rect 20349 26327 20407 26333
rect 20714 26324 20720 26336
rect 20772 26324 20778 26376
rect 20824 26373 20852 26404
rect 20990 26392 20996 26404
rect 21048 26392 21054 26444
rect 22002 26432 22008 26444
rect 21928 26404 22008 26432
rect 20809 26367 20867 26373
rect 20809 26333 20821 26367
rect 20855 26333 20867 26367
rect 20809 26327 20867 26333
rect 20901 26367 20959 26373
rect 20901 26333 20913 26367
rect 20947 26364 20959 26367
rect 21082 26364 21088 26376
rect 20947 26336 21088 26364
rect 20947 26333 20959 26336
rect 20901 26327 20959 26333
rect 21082 26324 21088 26336
rect 21140 26324 21146 26376
rect 21542 26324 21548 26376
rect 21600 26364 21606 26376
rect 21928 26373 21956 26404
rect 22002 26392 22008 26404
rect 22060 26392 22066 26444
rect 22189 26435 22247 26441
rect 22189 26401 22201 26435
rect 22235 26432 22247 26435
rect 22235 26404 22876 26432
rect 22235 26401 22247 26404
rect 22189 26395 22247 26401
rect 21913 26367 21971 26373
rect 21913 26364 21925 26367
rect 21600 26336 21925 26364
rect 21600 26324 21606 26336
rect 21913 26333 21925 26336
rect 21959 26333 21971 26367
rect 21913 26327 21971 26333
rect 22094 26324 22100 26376
rect 22152 26364 22158 26376
rect 22646 26364 22652 26376
rect 22152 26336 22197 26364
rect 22607 26336 22652 26364
rect 22152 26324 22158 26336
rect 22646 26324 22652 26336
rect 22704 26324 22710 26376
rect 22848 26373 22876 26404
rect 23658 26392 23664 26444
rect 23716 26432 23722 26444
rect 26053 26435 26111 26441
rect 26053 26432 26065 26435
rect 23716 26404 26065 26432
rect 23716 26392 23722 26404
rect 26053 26401 26065 26404
rect 26099 26401 26111 26435
rect 26878 26432 26884 26444
rect 26839 26404 26884 26432
rect 26053 26395 26111 26401
rect 26878 26392 26884 26404
rect 26936 26392 26942 26444
rect 22833 26367 22891 26373
rect 22833 26333 22845 26367
rect 22879 26364 22891 26367
rect 23290 26364 23296 26376
rect 22879 26336 23296 26364
rect 22879 26333 22891 26336
rect 22833 26327 22891 26333
rect 23290 26324 23296 26336
rect 23348 26324 23354 26376
rect 23477 26367 23535 26373
rect 23477 26333 23489 26367
rect 23523 26333 23535 26367
rect 24394 26364 24400 26376
rect 24355 26336 24400 26364
rect 23477 26327 23535 26333
rect 17954 26296 17960 26308
rect 17092 26268 17448 26296
rect 17915 26268 17960 26296
rect 17092 26256 17098 26268
rect 17954 26256 17960 26268
rect 18012 26256 18018 26308
rect 19518 26256 19524 26308
rect 19576 26296 19582 26308
rect 23492 26296 23520 26327
rect 24394 26324 24400 26336
rect 24452 26324 24458 26376
rect 24581 26367 24639 26373
rect 24581 26333 24593 26367
rect 24627 26364 24639 26367
rect 24946 26364 24952 26376
rect 24627 26336 24952 26364
rect 24627 26333 24639 26336
rect 24581 26327 24639 26333
rect 24946 26324 24952 26336
rect 25004 26324 25010 26376
rect 25866 26324 25872 26376
rect 25924 26364 25930 26376
rect 25961 26367 26019 26373
rect 25961 26364 25973 26367
rect 25924 26336 25973 26364
rect 25924 26324 25930 26336
rect 25961 26333 25973 26336
rect 26007 26333 26019 26367
rect 28442 26364 28448 26376
rect 25961 26327 26019 26333
rect 26896 26336 28448 26364
rect 19576 26268 23520 26296
rect 24765 26299 24823 26305
rect 19576 26256 19582 26268
rect 24765 26265 24777 26299
rect 24811 26296 24823 26299
rect 26142 26296 26148 26308
rect 24811 26268 26148 26296
rect 24811 26265 24823 26268
rect 24765 26259 24823 26265
rect 26142 26256 26148 26268
rect 26200 26256 26206 26308
rect 26896 26296 26924 26336
rect 28442 26324 28448 26336
rect 28500 26324 28506 26376
rect 26252 26268 26924 26296
rect 15979 26200 16068 26228
rect 15979 26197 15991 26200
rect 15933 26191 15991 26197
rect 17218 26188 17224 26240
rect 17276 26228 17282 26240
rect 17586 26228 17592 26240
rect 17276 26200 17592 26228
rect 17276 26188 17282 26200
rect 17586 26188 17592 26200
rect 17644 26228 17650 26240
rect 18157 26231 18215 26237
rect 18157 26228 18169 26231
rect 17644 26200 18169 26228
rect 17644 26188 17650 26200
rect 18157 26197 18169 26200
rect 18203 26197 18215 26231
rect 18322 26228 18328 26240
rect 18283 26200 18328 26228
rect 18157 26191 18215 26197
rect 18322 26188 18328 26200
rect 18380 26188 18386 26240
rect 20254 26188 20260 26240
rect 20312 26228 20318 26240
rect 20438 26228 20444 26240
rect 20312 26200 20444 26228
rect 20312 26188 20318 26200
rect 20438 26188 20444 26200
rect 20496 26188 20502 26240
rect 20898 26188 20904 26240
rect 20956 26228 20962 26240
rect 23474 26228 23480 26240
rect 20956 26200 23480 26228
rect 20956 26188 20962 26200
rect 23474 26188 23480 26200
rect 23532 26188 23538 26240
rect 25869 26231 25927 26237
rect 25869 26197 25881 26231
rect 25915 26228 25927 26231
rect 26252 26228 26280 26268
rect 26970 26256 26976 26308
rect 27028 26296 27034 26308
rect 27126 26299 27184 26305
rect 27126 26296 27138 26299
rect 27028 26268 27138 26296
rect 27028 26256 27034 26268
rect 27126 26265 27138 26268
rect 27172 26265 27184 26299
rect 27126 26259 27184 26265
rect 25915 26200 26280 26228
rect 25915 26197 25927 26200
rect 25869 26191 25927 26197
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 9030 26024 9036 26036
rect 7300 25996 9036 26024
rect 7300 25897 7328 25996
rect 9030 25984 9036 25996
rect 9088 25984 9094 26036
rect 9122 25984 9128 26036
rect 9180 26024 9186 26036
rect 9217 26027 9275 26033
rect 9217 26024 9229 26027
rect 9180 25996 9229 26024
rect 9180 25984 9186 25996
rect 9217 25993 9229 25996
rect 9263 25993 9275 26027
rect 11330 26024 11336 26036
rect 9217 25987 9275 25993
rect 9324 25996 11336 26024
rect 9324 25956 9352 25996
rect 11330 25984 11336 25996
rect 11388 25984 11394 26036
rect 12161 26027 12219 26033
rect 12161 25993 12173 26027
rect 12207 26024 12219 26027
rect 12250 26024 12256 26036
rect 12207 25996 12256 26024
rect 12207 25993 12219 25996
rect 12161 25987 12219 25993
rect 12250 25984 12256 25996
rect 12308 25984 12314 26036
rect 12434 25984 12440 26036
rect 12492 26024 12498 26036
rect 12713 26027 12771 26033
rect 12713 26024 12725 26027
rect 12492 25996 12725 26024
rect 12492 25984 12498 25996
rect 12713 25993 12725 25996
rect 12759 25993 12771 26027
rect 12713 25987 12771 25993
rect 15838 25984 15844 26036
rect 15896 26024 15902 26036
rect 16022 26024 16028 26036
rect 15896 25996 16028 26024
rect 15896 25984 15902 25996
rect 16022 25984 16028 25996
rect 16080 25984 16086 26036
rect 17957 26027 18015 26033
rect 17957 26024 17969 26027
rect 16132 25996 17969 26024
rect 7576 25928 9352 25956
rect 9585 25959 9643 25965
rect 7101 25891 7159 25897
rect 7101 25857 7113 25891
rect 7147 25857 7159 25891
rect 7101 25851 7159 25857
rect 7285 25891 7343 25897
rect 7285 25857 7297 25891
rect 7331 25857 7343 25891
rect 7285 25851 7343 25857
rect 7116 25684 7144 25851
rect 7193 25823 7251 25829
rect 7193 25789 7205 25823
rect 7239 25820 7251 25823
rect 7576 25820 7604 25928
rect 9585 25925 9597 25959
rect 9631 25956 9643 25959
rect 9766 25956 9772 25968
rect 9631 25928 9772 25956
rect 9631 25925 9643 25928
rect 9585 25919 9643 25925
rect 9766 25916 9772 25928
rect 9824 25916 9830 25968
rect 10965 25959 11023 25965
rect 10965 25925 10977 25959
rect 11011 25956 11023 25959
rect 11514 25956 11520 25968
rect 11011 25928 11520 25956
rect 11011 25925 11023 25928
rect 10965 25919 11023 25925
rect 11514 25916 11520 25928
rect 11572 25956 11578 25968
rect 14182 25956 14188 25968
rect 11572 25928 14188 25956
rect 11572 25916 11578 25928
rect 14182 25916 14188 25928
rect 14240 25916 14246 25968
rect 14360 25959 14418 25965
rect 14360 25925 14372 25959
rect 14406 25956 14418 25959
rect 16132 25956 16160 25996
rect 17957 25993 17969 25996
rect 18003 25993 18015 26027
rect 17957 25987 18015 25993
rect 19981 26027 20039 26033
rect 19981 25993 19993 26027
rect 20027 26024 20039 26027
rect 20990 26024 20996 26036
rect 20027 25996 20996 26024
rect 20027 25993 20039 25996
rect 19981 25987 20039 25993
rect 20990 25984 20996 25996
rect 21048 25984 21054 26036
rect 22278 25984 22284 26036
rect 22336 25984 22342 26036
rect 23569 26027 23627 26033
rect 23569 25993 23581 26027
rect 23615 26024 23627 26027
rect 23658 26024 23664 26036
rect 23615 25996 23664 26024
rect 23615 25993 23627 25996
rect 23569 25987 23627 25993
rect 23658 25984 23664 25996
rect 23716 25984 23722 26036
rect 25501 26027 25559 26033
rect 25501 25993 25513 26027
rect 25547 26024 25559 26027
rect 26234 26024 26240 26036
rect 25547 25996 26240 26024
rect 25547 25993 25559 25996
rect 25501 25987 25559 25993
rect 26234 25984 26240 25996
rect 26292 26024 26298 26036
rect 26878 26024 26884 26036
rect 26292 25996 26884 26024
rect 26292 25984 26298 25996
rect 26878 25984 26884 25996
rect 26936 25984 26942 26036
rect 14406 25928 16160 25956
rect 14406 25925 14418 25928
rect 14360 25919 14418 25925
rect 16298 25916 16304 25968
rect 16356 25956 16362 25968
rect 22296 25956 22324 25984
rect 23382 25956 23388 25968
rect 16356 25928 17908 25956
rect 22296 25928 23388 25956
rect 16356 25916 16362 25928
rect 7742 25888 7748 25900
rect 7703 25860 7748 25888
rect 7742 25848 7748 25860
rect 7800 25848 7806 25900
rect 7926 25888 7932 25900
rect 7887 25860 7932 25888
rect 7926 25848 7932 25860
rect 7984 25848 7990 25900
rect 8110 25888 8116 25900
rect 8071 25860 8116 25888
rect 8110 25848 8116 25860
rect 8168 25848 8174 25900
rect 8297 25891 8355 25897
rect 8297 25857 8309 25891
rect 8343 25888 8355 25891
rect 8386 25888 8392 25900
rect 8343 25860 8392 25888
rect 8343 25857 8355 25860
rect 8297 25851 8355 25857
rect 8386 25848 8392 25860
rect 8444 25848 8450 25900
rect 9398 25848 9404 25900
rect 9456 25888 9462 25900
rect 10778 25888 10784 25900
rect 9456 25860 9904 25888
rect 10739 25860 10784 25888
rect 9456 25848 9462 25860
rect 7239 25792 7604 25820
rect 7239 25789 7251 25792
rect 7193 25783 7251 25789
rect 8018 25780 8024 25832
rect 8076 25820 8082 25832
rect 9674 25820 9680 25832
rect 8076 25792 8121 25820
rect 9635 25792 9680 25820
rect 8076 25780 8082 25792
rect 9674 25780 9680 25792
rect 9732 25780 9738 25832
rect 9876 25829 9904 25860
rect 10778 25848 10784 25860
rect 10836 25848 10842 25900
rect 12069 25891 12127 25897
rect 12069 25857 12081 25891
rect 12115 25857 12127 25891
rect 12069 25851 12127 25857
rect 12897 25891 12955 25897
rect 12897 25857 12909 25891
rect 12943 25888 12955 25891
rect 13262 25888 13268 25900
rect 12943 25860 13268 25888
rect 12943 25857 12955 25860
rect 12897 25851 12955 25857
rect 9861 25823 9919 25829
rect 9861 25789 9873 25823
rect 9907 25820 9919 25823
rect 12084 25820 12112 25851
rect 13262 25848 13268 25860
rect 13320 25848 13326 25900
rect 14090 25888 14096 25900
rect 14051 25860 14096 25888
rect 14090 25848 14096 25860
rect 14148 25848 14154 25900
rect 17880 25897 17908 25928
rect 15933 25891 15991 25897
rect 14200 25860 15148 25888
rect 12986 25820 12992 25832
rect 9907 25792 12112 25820
rect 12947 25792 12992 25820
rect 9907 25789 9919 25792
rect 9861 25783 9919 25789
rect 12986 25780 12992 25792
rect 13044 25780 13050 25832
rect 13081 25823 13139 25829
rect 13081 25789 13093 25823
rect 13127 25789 13139 25823
rect 13081 25783 13139 25789
rect 10778 25752 10784 25764
rect 8312 25724 10784 25752
rect 8312 25684 8340 25724
rect 10778 25712 10784 25724
rect 10836 25752 10842 25764
rect 12342 25752 12348 25764
rect 10836 25724 12348 25752
rect 10836 25712 10842 25724
rect 12342 25712 12348 25724
rect 12400 25712 12406 25764
rect 13096 25752 13124 25783
rect 13170 25780 13176 25832
rect 13228 25820 13234 25832
rect 13228 25792 13273 25820
rect 13228 25780 13234 25792
rect 13722 25780 13728 25832
rect 13780 25820 13786 25832
rect 14200 25820 14228 25860
rect 13780 25792 14228 25820
rect 15120 25820 15148 25860
rect 15933 25857 15945 25891
rect 15979 25888 15991 25891
rect 17037 25891 17095 25897
rect 17037 25888 17049 25891
rect 15979 25860 17049 25888
rect 15979 25857 15991 25860
rect 15933 25851 15991 25857
rect 16114 25820 16120 25832
rect 15120 25792 16120 25820
rect 13780 25780 13786 25792
rect 16114 25780 16120 25792
rect 16172 25780 16178 25832
rect 13354 25752 13360 25764
rect 13096 25724 13360 25752
rect 13354 25712 13360 25724
rect 13412 25712 13418 25764
rect 15194 25712 15200 25764
rect 15252 25752 15258 25764
rect 15473 25755 15531 25761
rect 15473 25752 15485 25755
rect 15252 25724 15485 25752
rect 15252 25712 15258 25724
rect 15473 25721 15485 25724
rect 15519 25752 15531 25755
rect 16224 25752 16252 25860
rect 17037 25857 17049 25860
rect 17083 25857 17095 25891
rect 17037 25851 17095 25857
rect 17865 25891 17923 25897
rect 17865 25857 17877 25891
rect 17911 25857 17923 25891
rect 17865 25851 17923 25857
rect 17954 25848 17960 25900
rect 18012 25888 18018 25900
rect 18049 25891 18107 25897
rect 18049 25888 18061 25891
rect 18012 25860 18061 25888
rect 18012 25848 18018 25860
rect 18049 25857 18061 25860
rect 18095 25857 18107 25891
rect 18877 25891 18935 25897
rect 18877 25888 18889 25891
rect 18049 25851 18107 25857
rect 18156 25860 18889 25888
rect 16758 25780 16764 25832
rect 16816 25820 16822 25832
rect 16945 25823 17003 25829
rect 16945 25820 16957 25823
rect 16816 25792 16957 25820
rect 16816 25780 16822 25792
rect 16945 25789 16957 25792
rect 16991 25789 17003 25823
rect 16945 25783 17003 25789
rect 17494 25780 17500 25832
rect 17552 25820 17558 25832
rect 18156 25820 18184 25860
rect 18877 25857 18889 25860
rect 18923 25857 18935 25891
rect 18877 25851 18935 25857
rect 19426 25848 19432 25900
rect 19484 25888 19490 25900
rect 19797 25891 19855 25897
rect 19797 25888 19809 25891
rect 19484 25860 19809 25888
rect 19484 25848 19490 25860
rect 19797 25857 19809 25860
rect 19843 25857 19855 25891
rect 19797 25851 19855 25857
rect 19981 25891 20039 25897
rect 19981 25857 19993 25891
rect 20027 25857 20039 25891
rect 19981 25851 20039 25857
rect 20441 25891 20499 25897
rect 20441 25857 20453 25891
rect 20487 25888 20499 25891
rect 20806 25888 20812 25900
rect 20487 25860 20812 25888
rect 20487 25857 20499 25860
rect 20441 25851 20499 25857
rect 18782 25820 18788 25832
rect 17552 25792 18184 25820
rect 18743 25792 18788 25820
rect 17552 25780 17558 25792
rect 18782 25780 18788 25792
rect 18840 25780 18846 25832
rect 19996 25820 20024 25851
rect 20806 25848 20812 25860
rect 20864 25848 20870 25900
rect 22005 25891 22063 25897
rect 22005 25857 22017 25891
rect 22051 25857 22063 25891
rect 22005 25851 22063 25857
rect 19306 25792 20024 25820
rect 17402 25752 17408 25764
rect 15519 25724 16252 25752
rect 17363 25724 17408 25752
rect 15519 25721 15531 25724
rect 15473 25715 15531 25721
rect 17402 25712 17408 25724
rect 17460 25712 17466 25764
rect 17678 25712 17684 25764
rect 17736 25752 17742 25764
rect 19306 25752 19334 25792
rect 17736 25724 19334 25752
rect 19996 25752 20024 25792
rect 20622 25780 20628 25832
rect 20680 25820 20686 25832
rect 20717 25823 20775 25829
rect 20717 25820 20729 25823
rect 20680 25792 20729 25820
rect 20680 25780 20686 25792
rect 20717 25789 20729 25792
rect 20763 25820 20775 25823
rect 21450 25820 21456 25832
rect 20763 25792 21456 25820
rect 20763 25789 20775 25792
rect 20717 25783 20775 25789
rect 21450 25780 21456 25792
rect 21508 25780 21514 25832
rect 21910 25780 21916 25832
rect 21968 25780 21974 25832
rect 21266 25752 21272 25764
rect 19996 25724 21272 25752
rect 17736 25712 17742 25724
rect 21266 25712 21272 25724
rect 21324 25752 21330 25764
rect 21928 25752 21956 25780
rect 21324 25724 21956 25752
rect 22020 25752 22048 25851
rect 22094 25848 22100 25900
rect 22152 25888 22158 25900
rect 22278 25888 22284 25900
rect 22152 25860 22197 25888
rect 22239 25860 22284 25888
rect 22152 25848 22158 25860
rect 22278 25848 22284 25860
rect 22336 25848 22342 25900
rect 22388 25897 22416 25928
rect 22373 25891 22431 25897
rect 22373 25857 22385 25891
rect 22419 25857 22431 25891
rect 22373 25851 22431 25857
rect 22554 25848 22560 25900
rect 22612 25888 22618 25900
rect 23032 25897 23060 25928
rect 23382 25916 23388 25928
rect 23440 25916 23446 25968
rect 25409 25959 25467 25965
rect 25409 25925 25421 25959
rect 25455 25956 25467 25959
rect 26786 25956 26792 25968
rect 25455 25928 26792 25956
rect 25455 25925 25467 25928
rect 25409 25919 25467 25925
rect 26786 25916 26792 25928
rect 26844 25916 26850 25968
rect 22833 25891 22891 25897
rect 22833 25888 22845 25891
rect 22612 25860 22845 25888
rect 22612 25848 22618 25860
rect 22833 25857 22845 25860
rect 22879 25857 22891 25891
rect 22833 25851 22891 25857
rect 23017 25891 23075 25897
rect 23017 25857 23029 25891
rect 23063 25857 23075 25891
rect 23474 25888 23480 25900
rect 23435 25860 23480 25888
rect 23017 25851 23075 25857
rect 23474 25848 23480 25860
rect 23532 25848 23538 25900
rect 23658 25848 23664 25900
rect 23716 25897 23722 25900
rect 23716 25891 23731 25897
rect 23719 25857 23731 25891
rect 23716 25851 23731 25857
rect 23716 25848 23722 25851
rect 24026 25848 24032 25900
rect 24084 25888 24090 25900
rect 24305 25891 24363 25897
rect 24305 25888 24317 25891
rect 24084 25860 24317 25888
rect 24084 25848 24090 25860
rect 24305 25857 24317 25860
rect 24351 25857 24363 25891
rect 24305 25851 24363 25857
rect 26142 25848 26148 25900
rect 26200 25888 26206 25900
rect 26237 25891 26295 25897
rect 26237 25888 26249 25891
rect 26200 25860 26249 25888
rect 26200 25848 26206 25860
rect 26237 25857 26249 25860
rect 26283 25857 26295 25891
rect 26896 25888 26924 25984
rect 27424 25959 27482 25965
rect 27424 25925 27436 25959
rect 27470 25956 27482 25959
rect 27522 25956 27528 25968
rect 27470 25928 27528 25956
rect 27470 25925 27482 25928
rect 27424 25919 27482 25925
rect 27522 25916 27528 25928
rect 27580 25916 27586 25968
rect 27157 25891 27215 25897
rect 27157 25888 27169 25891
rect 26896 25860 27169 25888
rect 26237 25851 26295 25857
rect 27157 25857 27169 25860
rect 27203 25857 27215 25891
rect 27157 25851 27215 25857
rect 22925 25823 22983 25829
rect 22925 25789 22937 25823
rect 22971 25820 22983 25823
rect 24670 25820 24676 25832
rect 22971 25792 24676 25820
rect 22971 25789 22983 25792
rect 22925 25783 22983 25789
rect 24670 25780 24676 25792
rect 24728 25780 24734 25832
rect 25498 25752 25504 25764
rect 22020 25724 25504 25752
rect 21324 25712 21330 25724
rect 25498 25712 25504 25724
rect 25556 25712 25562 25764
rect 25774 25712 25780 25764
rect 25832 25752 25838 25764
rect 26053 25755 26111 25761
rect 26053 25752 26065 25755
rect 25832 25724 26065 25752
rect 25832 25712 25838 25724
rect 26053 25721 26065 25724
rect 26099 25721 26111 25755
rect 26053 25715 26111 25721
rect 8478 25684 8484 25696
rect 7116 25656 8340 25684
rect 8439 25656 8484 25684
rect 8478 25644 8484 25656
rect 8536 25644 8542 25696
rect 9030 25644 9036 25696
rect 9088 25684 9094 25696
rect 10042 25684 10048 25696
rect 9088 25656 10048 25684
rect 9088 25644 9094 25656
rect 10042 25644 10048 25656
rect 10100 25644 10106 25696
rect 13262 25644 13268 25696
rect 13320 25684 13326 25696
rect 17696 25684 17724 25712
rect 13320 25656 17724 25684
rect 19153 25687 19211 25693
rect 13320 25644 13326 25656
rect 19153 25653 19165 25687
rect 19199 25684 19211 25687
rect 19334 25684 19340 25696
rect 19199 25656 19340 25684
rect 19199 25653 19211 25656
rect 19153 25647 19211 25653
rect 19334 25644 19340 25656
rect 19392 25644 19398 25696
rect 20438 25644 20444 25696
rect 20496 25684 20502 25696
rect 21821 25687 21879 25693
rect 21821 25684 21833 25687
rect 20496 25656 21833 25684
rect 20496 25644 20502 25656
rect 21821 25653 21833 25656
rect 21867 25653 21879 25687
rect 21821 25647 21879 25653
rect 21910 25644 21916 25696
rect 21968 25684 21974 25696
rect 24026 25684 24032 25696
rect 21968 25656 24032 25684
rect 21968 25644 21974 25656
rect 24026 25644 24032 25656
rect 24084 25644 24090 25696
rect 24121 25687 24179 25693
rect 24121 25653 24133 25687
rect 24167 25684 24179 25687
rect 24394 25684 24400 25696
rect 24167 25656 24400 25684
rect 24167 25653 24179 25656
rect 24121 25647 24179 25653
rect 24394 25644 24400 25656
rect 24452 25644 24458 25696
rect 28442 25644 28448 25696
rect 28500 25684 28506 25696
rect 28537 25687 28595 25693
rect 28537 25684 28549 25687
rect 28500 25656 28549 25684
rect 28500 25644 28506 25656
rect 28537 25653 28549 25656
rect 28583 25653 28595 25687
rect 28537 25647 28595 25653
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 8018 25440 8024 25492
rect 8076 25480 8082 25492
rect 9585 25483 9643 25489
rect 9585 25480 9597 25483
rect 8076 25452 9597 25480
rect 8076 25440 8082 25452
rect 9585 25449 9597 25452
rect 9631 25449 9643 25483
rect 9585 25443 9643 25449
rect 9674 25440 9680 25492
rect 9732 25480 9738 25492
rect 10137 25483 10195 25489
rect 10137 25480 10149 25483
rect 9732 25452 10149 25480
rect 9732 25440 9738 25452
rect 10137 25449 10149 25452
rect 10183 25449 10195 25483
rect 10137 25443 10195 25449
rect 10318 25440 10324 25492
rect 10376 25480 10382 25492
rect 10686 25480 10692 25492
rect 10376 25452 10692 25480
rect 10376 25440 10382 25452
rect 10686 25440 10692 25452
rect 10744 25440 10750 25492
rect 11885 25483 11943 25489
rect 11885 25449 11897 25483
rect 11931 25449 11943 25483
rect 11885 25443 11943 25449
rect 8386 25412 8392 25424
rect 8347 25384 8392 25412
rect 8386 25372 8392 25384
rect 8444 25412 8450 25424
rect 9122 25412 9128 25424
rect 8444 25384 9128 25412
rect 8444 25372 8450 25384
rect 9122 25372 9128 25384
rect 9180 25372 9186 25424
rect 11149 25415 11207 25421
rect 11149 25381 11161 25415
rect 11195 25381 11207 25415
rect 11900 25412 11928 25443
rect 12158 25440 12164 25492
rect 12216 25480 12222 25492
rect 12529 25483 12587 25489
rect 12529 25480 12541 25483
rect 12216 25452 12541 25480
rect 12216 25440 12222 25452
rect 12529 25449 12541 25452
rect 12575 25449 12587 25483
rect 12529 25443 12587 25449
rect 14369 25483 14427 25489
rect 14369 25449 14381 25483
rect 14415 25480 14427 25483
rect 14918 25480 14924 25492
rect 14415 25452 14924 25480
rect 14415 25449 14427 25452
rect 14369 25443 14427 25449
rect 14918 25440 14924 25452
rect 14976 25440 14982 25492
rect 15102 25480 15108 25492
rect 15063 25452 15108 25480
rect 15102 25440 15108 25452
rect 15160 25440 15166 25492
rect 15562 25440 15568 25492
rect 15620 25480 15626 25492
rect 16022 25480 16028 25492
rect 15620 25452 16028 25480
rect 15620 25440 15626 25452
rect 16022 25440 16028 25452
rect 16080 25440 16086 25492
rect 17402 25480 17408 25492
rect 17363 25452 17408 25480
rect 17402 25440 17408 25452
rect 17460 25440 17466 25492
rect 17586 25480 17592 25492
rect 17547 25452 17592 25480
rect 17586 25440 17592 25452
rect 17644 25440 17650 25492
rect 19242 25440 19248 25492
rect 19300 25480 19306 25492
rect 19429 25483 19487 25489
rect 19429 25480 19441 25483
rect 19300 25452 19441 25480
rect 19300 25440 19306 25452
rect 19429 25449 19441 25452
rect 19475 25449 19487 25483
rect 19429 25443 19487 25449
rect 20441 25483 20499 25489
rect 20441 25449 20453 25483
rect 20487 25480 20499 25483
rect 21177 25483 21235 25489
rect 21177 25480 21189 25483
rect 20487 25452 21189 25480
rect 20487 25449 20499 25452
rect 20441 25443 20499 25449
rect 21177 25449 21189 25452
rect 21223 25449 21235 25483
rect 21177 25443 21235 25449
rect 22278 25440 22284 25492
rect 22336 25480 22342 25492
rect 22465 25483 22523 25489
rect 22465 25480 22477 25483
rect 22336 25452 22477 25480
rect 22336 25440 22342 25452
rect 22465 25449 22477 25452
rect 22511 25449 22523 25483
rect 22465 25443 22523 25449
rect 26881 25483 26939 25489
rect 26881 25449 26893 25483
rect 26927 25480 26939 25483
rect 26970 25480 26976 25492
rect 26927 25452 26976 25480
rect 26927 25449 26939 25452
rect 26881 25443 26939 25449
rect 26970 25440 26976 25452
rect 27028 25440 27034 25492
rect 13998 25412 14004 25424
rect 11900 25384 14004 25412
rect 11149 25375 11207 25381
rect 8662 25304 8668 25356
rect 8720 25344 8726 25356
rect 9401 25347 9459 25353
rect 9401 25344 9413 25347
rect 8720 25316 9413 25344
rect 8720 25304 8726 25316
rect 9401 25313 9413 25316
rect 9447 25313 9459 25347
rect 9401 25307 9459 25313
rect 9766 25304 9772 25356
rect 9824 25344 9830 25356
rect 10410 25344 10416 25356
rect 9824 25316 10416 25344
rect 9824 25304 9830 25316
rect 10410 25304 10416 25316
rect 10468 25344 10474 25356
rect 10781 25347 10839 25353
rect 10781 25344 10793 25347
rect 10468 25316 10793 25344
rect 10468 25304 10474 25316
rect 10781 25313 10793 25316
rect 10827 25313 10839 25347
rect 11164 25344 11192 25375
rect 13998 25372 14004 25384
rect 14056 25372 14062 25424
rect 15010 25372 15016 25424
rect 15068 25412 15074 25424
rect 15068 25384 15608 25412
rect 15068 25372 15074 25384
rect 12894 25344 12900 25356
rect 11164 25316 12900 25344
rect 10781 25307 10839 25313
rect 7006 25276 7012 25288
rect 6967 25248 7012 25276
rect 7006 25236 7012 25248
rect 7064 25236 7070 25288
rect 7276 25279 7334 25285
rect 7276 25245 7288 25279
rect 7322 25276 7334 25279
rect 8478 25276 8484 25288
rect 7322 25248 8484 25276
rect 7322 25245 7334 25248
rect 7276 25239 7334 25245
rect 8478 25236 8484 25248
rect 8536 25236 8542 25288
rect 9309 25279 9367 25285
rect 9309 25245 9321 25279
rect 9355 25245 9367 25279
rect 9309 25239 9367 25245
rect 8386 25168 8392 25220
rect 8444 25208 8450 25220
rect 9324 25208 9352 25239
rect 9950 25236 9956 25288
rect 10008 25276 10014 25288
rect 11716 25285 11744 25316
rect 12894 25304 12900 25316
rect 12952 25304 12958 25356
rect 14550 25344 14556 25356
rect 14384 25316 14556 25344
rect 10045 25279 10103 25285
rect 10045 25276 10057 25279
rect 10008 25248 10057 25276
rect 10008 25236 10014 25248
rect 10045 25245 10057 25248
rect 10091 25245 10103 25279
rect 10045 25239 10103 25245
rect 10965 25279 11023 25285
rect 10965 25245 10977 25279
rect 11011 25245 11023 25279
rect 10965 25239 11023 25245
rect 11701 25279 11759 25285
rect 11701 25245 11713 25279
rect 11747 25245 11759 25279
rect 11701 25239 11759 25245
rect 8444 25180 9352 25208
rect 8444 25168 8450 25180
rect 10134 25168 10140 25220
rect 10192 25208 10198 25220
rect 10689 25211 10747 25217
rect 10689 25208 10701 25211
rect 10192 25180 10701 25208
rect 10192 25168 10198 25180
rect 10689 25177 10701 25180
rect 10735 25177 10747 25211
rect 10980 25208 11008 25239
rect 11790 25236 11796 25288
rect 11848 25276 11854 25288
rect 11848 25248 11893 25276
rect 11848 25236 11854 25248
rect 12342 25236 12348 25288
rect 12400 25276 12406 25288
rect 14384 25285 14412 25316
rect 14550 25304 14556 25316
rect 14608 25344 14614 25356
rect 15102 25344 15108 25356
rect 14608 25316 15108 25344
rect 14608 25304 14614 25316
rect 15102 25304 15108 25316
rect 15160 25304 15166 25356
rect 12713 25279 12771 25285
rect 12713 25276 12725 25279
rect 12400 25248 12725 25276
rect 12400 25236 12406 25248
rect 12713 25245 12725 25248
rect 12759 25245 12771 25279
rect 12713 25239 12771 25245
rect 12989 25279 13047 25285
rect 12989 25245 13001 25279
rect 13035 25245 13047 25279
rect 12989 25239 13047 25245
rect 14369 25279 14427 25285
rect 14369 25245 14381 25279
rect 14415 25245 14427 25279
rect 14369 25239 14427 25245
rect 14645 25279 14703 25285
rect 14645 25245 14657 25279
rect 14691 25276 14703 25279
rect 15194 25276 15200 25288
rect 14691 25248 15200 25276
rect 14691 25245 14703 25248
rect 14645 25239 14703 25245
rect 11606 25208 11612 25220
rect 10980 25180 11612 25208
rect 10689 25171 10747 25177
rect 11606 25168 11612 25180
rect 11664 25208 11670 25220
rect 12250 25208 12256 25220
rect 11664 25180 12256 25208
rect 11664 25168 11670 25180
rect 12250 25168 12256 25180
rect 12308 25168 12314 25220
rect 13004 25208 13032 25239
rect 15194 25236 15200 25248
rect 15252 25236 15258 25288
rect 15289 25279 15347 25285
rect 15289 25245 15301 25279
rect 15335 25245 15347 25279
rect 15289 25239 15347 25245
rect 15381 25279 15439 25285
rect 15381 25245 15393 25279
rect 15427 25276 15439 25279
rect 15580 25276 15608 25384
rect 16114 25372 16120 25424
rect 16172 25412 16178 25424
rect 20625 25415 20683 25421
rect 20625 25412 20637 25415
rect 16172 25384 20637 25412
rect 16172 25372 16178 25384
rect 20625 25381 20637 25384
rect 20671 25381 20683 25415
rect 22922 25412 22928 25424
rect 20625 25375 20683 25381
rect 22572 25384 22928 25412
rect 17770 25344 17776 25356
rect 16684 25316 17776 25344
rect 16574 25276 16580 25288
rect 15427 25248 16580 25276
rect 15427 25245 15439 25248
rect 15381 25239 15439 25245
rect 12406 25180 13032 25208
rect 15304 25208 15332 25239
rect 16574 25236 16580 25248
rect 16632 25236 16638 25288
rect 16684 25285 16712 25316
rect 17770 25304 17776 25316
rect 17828 25304 17834 25356
rect 20990 25304 20996 25356
rect 21048 25344 21054 25356
rect 22094 25344 22100 25356
rect 21048 25316 22100 25344
rect 21048 25304 21054 25316
rect 16669 25279 16727 25285
rect 16669 25245 16681 25279
rect 16715 25245 16727 25279
rect 20714 25276 20720 25288
rect 16669 25239 16727 25245
rect 19996 25248 20720 25276
rect 15304 25180 15424 25208
rect 8846 25100 8852 25152
rect 8904 25140 8910 25152
rect 8941 25143 8999 25149
rect 8941 25140 8953 25143
rect 8904 25112 8953 25140
rect 8904 25100 8910 25112
rect 8941 25109 8953 25112
rect 8987 25140 8999 25143
rect 11974 25140 11980 25152
rect 8987 25112 11980 25140
rect 8987 25109 8999 25112
rect 8941 25103 8999 25109
rect 11974 25100 11980 25112
rect 12032 25100 12038 25152
rect 12069 25143 12127 25149
rect 12069 25109 12081 25143
rect 12115 25140 12127 25143
rect 12406 25140 12434 25180
rect 12115 25112 12434 25140
rect 12897 25143 12955 25149
rect 12115 25109 12127 25112
rect 12069 25103 12127 25109
rect 12897 25109 12909 25143
rect 12943 25140 12955 25143
rect 13262 25140 13268 25152
rect 12943 25112 13268 25140
rect 12943 25109 12955 25112
rect 12897 25103 12955 25109
rect 13262 25100 13268 25112
rect 13320 25100 13326 25152
rect 13354 25100 13360 25152
rect 13412 25140 13418 25152
rect 14553 25143 14611 25149
rect 14553 25140 14565 25143
rect 13412 25112 14565 25140
rect 13412 25100 13418 25112
rect 14553 25109 14565 25112
rect 14599 25140 14611 25143
rect 14918 25140 14924 25152
rect 14599 25112 14924 25140
rect 14599 25109 14611 25112
rect 14553 25103 14611 25109
rect 14918 25100 14924 25112
rect 14976 25100 14982 25152
rect 15396 25140 15424 25180
rect 15470 25168 15476 25220
rect 15528 25208 15534 25220
rect 15657 25211 15715 25217
rect 15657 25208 15669 25211
rect 15528 25180 15669 25208
rect 15528 25168 15534 25180
rect 15657 25177 15669 25180
rect 15703 25177 15715 25211
rect 15657 25171 15715 25177
rect 15746 25168 15752 25220
rect 15804 25208 15810 25220
rect 16592 25208 16620 25236
rect 17218 25208 17224 25220
rect 15804 25180 15849 25208
rect 16592 25180 16804 25208
rect 17179 25180 17224 25208
rect 15804 25168 15810 25180
rect 16206 25140 16212 25152
rect 15396 25112 16212 25140
rect 16206 25100 16212 25112
rect 16264 25140 16270 25152
rect 16669 25143 16727 25149
rect 16669 25140 16681 25143
rect 16264 25112 16681 25140
rect 16264 25100 16270 25112
rect 16669 25109 16681 25112
rect 16715 25109 16727 25143
rect 16776 25140 16804 25180
rect 17218 25168 17224 25180
rect 17276 25168 17282 25220
rect 18414 25168 18420 25220
rect 18472 25208 18478 25220
rect 19245 25211 19303 25217
rect 19245 25208 19257 25211
rect 18472 25180 19257 25208
rect 18472 25168 18478 25180
rect 19245 25177 19257 25180
rect 19291 25177 19303 25211
rect 19245 25171 19303 25177
rect 19334 25168 19340 25220
rect 19392 25208 19398 25220
rect 19461 25211 19519 25217
rect 19461 25208 19473 25211
rect 19392 25180 19473 25208
rect 19392 25168 19398 25180
rect 19461 25177 19473 25180
rect 19507 25208 19519 25211
rect 19996 25208 20024 25248
rect 20714 25236 20720 25248
rect 20772 25276 20778 25288
rect 20898 25276 20904 25288
rect 20772 25248 20904 25276
rect 20772 25236 20778 25248
rect 20898 25236 20904 25248
rect 20956 25236 20962 25288
rect 21358 25276 21364 25288
rect 21319 25248 21364 25276
rect 21358 25236 21364 25248
rect 21416 25236 21422 25288
rect 21468 25285 21496 25316
rect 22094 25304 22100 25316
rect 22152 25304 22158 25356
rect 21453 25279 21511 25285
rect 21453 25245 21465 25279
rect 21499 25245 21511 25279
rect 21453 25239 21511 25245
rect 21637 25279 21695 25285
rect 21637 25245 21649 25279
rect 21683 25245 21695 25279
rect 21637 25239 21695 25245
rect 21729 25279 21787 25285
rect 21729 25245 21741 25279
rect 21775 25276 21787 25279
rect 22572 25276 22600 25384
rect 22922 25372 22928 25384
rect 22980 25372 22986 25424
rect 26145 25415 26203 25421
rect 26145 25412 26157 25415
rect 23032 25384 26157 25412
rect 22738 25276 22744 25288
rect 21775 25248 22600 25276
rect 22699 25248 22744 25276
rect 21775 25245 21787 25248
rect 21729 25239 21787 25245
rect 19507 25180 20024 25208
rect 19507 25177 19519 25180
rect 19461 25171 19519 25177
rect 20070 25168 20076 25220
rect 20128 25208 20134 25220
rect 20128 25180 20173 25208
rect 20128 25168 20134 25180
rect 20438 25168 20444 25220
rect 20496 25217 20502 25220
rect 20496 25208 20508 25217
rect 21652 25208 21680 25239
rect 22738 25236 22744 25248
rect 22796 25236 22802 25288
rect 22833 25279 22891 25285
rect 22833 25245 22845 25279
rect 22879 25245 22891 25279
rect 22833 25239 22891 25245
rect 22925 25279 22983 25285
rect 22925 25245 22937 25279
rect 22971 25276 22983 25279
rect 23032 25276 23060 25384
rect 26145 25381 26157 25384
rect 26191 25381 26203 25415
rect 26145 25375 26203 25381
rect 24765 25347 24823 25353
rect 24765 25344 24777 25347
rect 23860 25316 24777 25344
rect 22971 25248 23060 25276
rect 22971 25245 22983 25248
rect 22925 25239 22983 25245
rect 22186 25208 22192 25220
rect 20496 25180 20541 25208
rect 21652 25180 22192 25208
rect 20496 25171 20508 25180
rect 20496 25168 20502 25171
rect 22186 25168 22192 25180
rect 22244 25168 22250 25220
rect 22848 25208 22876 25239
rect 23106 25236 23112 25288
rect 23164 25276 23170 25288
rect 23860 25285 23888 25316
rect 24765 25313 24777 25316
rect 24811 25313 24823 25347
rect 24765 25307 24823 25313
rect 23845 25279 23903 25285
rect 23164 25248 23209 25276
rect 23164 25236 23170 25248
rect 23845 25245 23857 25279
rect 23891 25245 23903 25279
rect 24394 25276 24400 25288
rect 24355 25248 24400 25276
rect 23845 25239 23903 25245
rect 24394 25236 24400 25248
rect 24452 25236 24458 25288
rect 24578 25276 24584 25288
rect 24539 25248 24584 25276
rect 24578 25236 24584 25248
rect 24636 25236 24642 25288
rect 25777 25279 25835 25285
rect 25777 25245 25789 25279
rect 25823 25276 25835 25279
rect 26878 25276 26884 25288
rect 25823 25248 26884 25276
rect 25823 25245 25835 25248
rect 25777 25239 25835 25245
rect 26878 25236 26884 25248
rect 26936 25236 26942 25288
rect 27062 25276 27068 25288
rect 27023 25248 27068 25276
rect 27062 25236 27068 25248
rect 27120 25236 27126 25288
rect 25682 25208 25688 25220
rect 22848 25180 25688 25208
rect 25682 25168 25688 25180
rect 25740 25168 25746 25220
rect 25961 25211 26019 25217
rect 25961 25177 25973 25211
rect 26007 25208 26019 25211
rect 26142 25208 26148 25220
rect 26007 25180 26148 25208
rect 26007 25177 26019 25180
rect 25961 25171 26019 25177
rect 26142 25168 26148 25180
rect 26200 25168 26206 25220
rect 17431 25143 17489 25149
rect 17431 25140 17443 25143
rect 16776 25112 17443 25140
rect 16669 25103 16727 25109
rect 17431 25109 17443 25112
rect 17477 25140 17489 25143
rect 18966 25140 18972 25152
rect 17477 25112 18972 25140
rect 17477 25109 17489 25112
rect 17431 25103 17489 25109
rect 18966 25100 18972 25112
rect 19024 25100 19030 25152
rect 19613 25143 19671 25149
rect 19613 25109 19625 25143
rect 19659 25140 19671 25143
rect 20806 25140 20812 25152
rect 19659 25112 20812 25140
rect 19659 25109 19671 25112
rect 19613 25103 19671 25109
rect 20806 25100 20812 25112
rect 20864 25100 20870 25152
rect 23658 25140 23664 25152
rect 23619 25112 23664 25140
rect 23658 25100 23664 25112
rect 23716 25100 23722 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 7926 24896 7932 24948
rect 7984 24936 7990 24948
rect 8113 24939 8171 24945
rect 8113 24936 8125 24939
rect 7984 24908 8125 24936
rect 7984 24896 7990 24908
rect 8113 24905 8125 24908
rect 8159 24905 8171 24939
rect 8113 24899 8171 24905
rect 8662 24896 8668 24948
rect 8720 24936 8726 24948
rect 8757 24939 8815 24945
rect 8757 24936 8769 24939
rect 8720 24908 8769 24936
rect 8720 24896 8726 24908
rect 8757 24905 8769 24908
rect 8803 24905 8815 24939
rect 9122 24936 9128 24948
rect 9083 24908 9128 24936
rect 8757 24899 8815 24905
rect 9122 24896 9128 24908
rect 9180 24896 9186 24948
rect 14458 24896 14464 24948
rect 14516 24936 14522 24948
rect 17954 24936 17960 24948
rect 14516 24908 17960 24936
rect 14516 24896 14522 24908
rect 17954 24896 17960 24908
rect 18012 24896 18018 24948
rect 22554 24896 22560 24948
rect 22612 24896 22618 24948
rect 25498 24936 25504 24948
rect 25459 24908 25504 24936
rect 25498 24896 25504 24908
rect 25556 24896 25562 24948
rect 8680 24868 8708 24896
rect 8128 24840 8708 24868
rect 9140 24868 9168 24896
rect 9140 24840 9720 24868
rect 8021 24803 8079 24809
rect 8021 24769 8033 24803
rect 8067 24800 8079 24803
rect 8128 24800 8156 24840
rect 8067 24772 8156 24800
rect 8205 24803 8263 24809
rect 8067 24769 8079 24772
rect 8021 24763 8079 24769
rect 8205 24769 8217 24803
rect 8251 24800 8263 24803
rect 8386 24800 8392 24812
rect 8251 24772 8392 24800
rect 8251 24769 8263 24772
rect 8205 24763 8263 24769
rect 8386 24760 8392 24772
rect 8444 24760 8450 24812
rect 9692 24800 9720 24840
rect 9950 24828 9956 24880
rect 10008 24868 10014 24880
rect 10321 24871 10379 24877
rect 10321 24868 10333 24871
rect 10008 24840 10333 24868
rect 10008 24828 10014 24840
rect 10321 24837 10333 24840
rect 10367 24837 10379 24871
rect 10321 24831 10379 24837
rect 10410 24828 10416 24880
rect 10468 24868 10474 24880
rect 14826 24868 14832 24880
rect 10468 24840 10513 24868
rect 13372 24840 14832 24868
rect 10468 24828 10474 24840
rect 10134 24800 10140 24812
rect 9692 24772 10140 24800
rect 10134 24760 10140 24772
rect 10192 24760 10198 24812
rect 10505 24803 10563 24809
rect 10505 24769 10517 24803
rect 10551 24800 10563 24803
rect 10594 24800 10600 24812
rect 10551 24772 10600 24800
rect 10551 24769 10563 24772
rect 10505 24763 10563 24769
rect 10594 24760 10600 24772
rect 10652 24760 10658 24812
rect 10686 24760 10692 24812
rect 10744 24800 10750 24812
rect 13372 24809 13400 24840
rect 14826 24828 14832 24840
rect 14884 24868 14890 24880
rect 15746 24868 15752 24880
rect 14884 24840 15752 24868
rect 14884 24828 14890 24840
rect 15746 24828 15752 24840
rect 15804 24868 15810 24880
rect 21266 24868 21272 24880
rect 15804 24840 15976 24868
rect 15804 24828 15810 24840
rect 11517 24803 11575 24809
rect 11517 24800 11529 24803
rect 10744 24772 11529 24800
rect 10744 24760 10750 24772
rect 11517 24769 11529 24772
rect 11563 24769 11575 24803
rect 11517 24763 11575 24769
rect 11701 24803 11759 24809
rect 11701 24769 11713 24803
rect 11747 24769 11759 24803
rect 11701 24763 11759 24769
rect 13081 24803 13139 24809
rect 13081 24769 13093 24803
rect 13127 24769 13139 24803
rect 13081 24763 13139 24769
rect 13357 24803 13415 24809
rect 13357 24769 13369 24803
rect 13403 24769 13415 24803
rect 13357 24763 13415 24769
rect 9214 24732 9220 24744
rect 9175 24704 9220 24732
rect 9214 24692 9220 24704
rect 9272 24692 9278 24744
rect 9398 24732 9404 24744
rect 9359 24704 9404 24732
rect 9398 24692 9404 24704
rect 9456 24692 9462 24744
rect 10042 24692 10048 24744
rect 10100 24732 10106 24744
rect 11716 24732 11744 24763
rect 10100 24704 11744 24732
rect 13096 24732 13124 24763
rect 13446 24760 13452 24812
rect 13504 24800 13510 24812
rect 13541 24803 13599 24809
rect 13541 24800 13553 24803
rect 13504 24772 13553 24800
rect 13504 24760 13510 24772
rect 13541 24769 13553 24772
rect 13587 24769 13599 24803
rect 13541 24763 13599 24769
rect 14185 24803 14243 24809
rect 14185 24769 14197 24803
rect 14231 24800 14243 24803
rect 14550 24800 14556 24812
rect 14231 24772 14556 24800
rect 14231 24769 14243 24772
rect 14185 24763 14243 24769
rect 14550 24760 14556 24772
rect 14608 24760 14614 24812
rect 15194 24760 15200 24812
rect 15252 24800 15258 24812
rect 15565 24803 15623 24809
rect 15252 24798 15424 24800
rect 15565 24798 15577 24803
rect 15252 24772 15577 24798
rect 15252 24760 15258 24772
rect 15396 24770 15577 24772
rect 15565 24769 15577 24770
rect 15611 24769 15623 24803
rect 15565 24763 15623 24769
rect 15657 24803 15715 24809
rect 15657 24769 15669 24803
rect 15703 24798 15715 24803
rect 15838 24800 15844 24812
rect 15764 24798 15844 24800
rect 15703 24772 15844 24798
rect 15703 24770 15792 24772
rect 15703 24769 15715 24770
rect 15657 24763 15715 24769
rect 15838 24760 15844 24772
rect 15896 24760 15902 24812
rect 13722 24732 13728 24744
rect 13096 24704 13728 24732
rect 10100 24692 10106 24704
rect 13722 24692 13728 24704
rect 13780 24692 13786 24744
rect 13998 24732 14004 24744
rect 13959 24704 14004 24732
rect 13998 24692 14004 24704
rect 14056 24692 14062 24744
rect 14642 24692 14648 24744
rect 14700 24732 14706 24744
rect 15289 24735 15347 24741
rect 15289 24732 15301 24735
rect 14700 24704 15301 24732
rect 14700 24692 14706 24704
rect 15289 24701 15301 24704
rect 15335 24701 15347 24735
rect 15289 24695 15347 24701
rect 15473 24735 15531 24741
rect 15473 24701 15485 24735
rect 15519 24701 15531 24735
rect 15473 24695 15531 24701
rect 15749 24735 15807 24741
rect 15749 24701 15761 24735
rect 15795 24732 15807 24735
rect 15948 24732 15976 24840
rect 21192 24840 21272 24868
rect 16206 24760 16212 24812
rect 16264 24800 16270 24812
rect 16669 24803 16727 24809
rect 16669 24800 16681 24803
rect 16264 24772 16681 24800
rect 16264 24760 16270 24772
rect 16669 24769 16681 24772
rect 16715 24769 16727 24803
rect 16942 24800 16948 24812
rect 16903 24772 16948 24800
rect 16669 24763 16727 24769
rect 16942 24760 16948 24772
rect 17000 24760 17006 24812
rect 17037 24803 17095 24809
rect 17037 24769 17049 24803
rect 17083 24800 17095 24803
rect 17678 24800 17684 24812
rect 17083 24772 17684 24800
rect 17083 24769 17095 24772
rect 17037 24763 17095 24769
rect 17678 24760 17684 24772
rect 17736 24760 17742 24812
rect 18049 24803 18107 24809
rect 18049 24769 18061 24803
rect 18095 24769 18107 24803
rect 18782 24800 18788 24812
rect 18743 24772 18788 24800
rect 18049 24763 18107 24769
rect 15795 24704 15976 24732
rect 15795 24701 15807 24704
rect 15749 24695 15807 24701
rect 13740 24664 13768 24692
rect 14369 24667 14427 24673
rect 14369 24664 14381 24667
rect 13740 24636 14381 24664
rect 14369 24633 14381 24636
rect 14415 24633 14427 24667
rect 14369 24627 14427 24633
rect 15102 24624 15108 24676
rect 15160 24664 15166 24676
rect 15488 24664 15516 24695
rect 17770 24692 17776 24744
rect 17828 24732 17834 24744
rect 18064 24732 18092 24763
rect 18782 24760 18788 24772
rect 18840 24760 18846 24812
rect 18966 24800 18972 24812
rect 18927 24772 18972 24800
rect 18966 24760 18972 24772
rect 19024 24760 19030 24812
rect 20898 24800 20904 24812
rect 20859 24772 20904 24800
rect 20898 24760 20904 24772
rect 20956 24760 20962 24812
rect 21192 24809 21220 24840
rect 21266 24828 21272 24840
rect 21324 24828 21330 24880
rect 21177 24803 21235 24809
rect 21177 24769 21189 24803
rect 21223 24769 21235 24803
rect 21177 24763 21235 24769
rect 21450 24760 21456 24812
rect 21508 24800 21514 24812
rect 22462 24800 22468 24812
rect 21508 24772 22468 24800
rect 21508 24760 21514 24772
rect 22462 24760 22468 24772
rect 22520 24760 22526 24812
rect 22572 24809 22600 24896
rect 23658 24828 23664 24880
rect 23716 24868 23722 24880
rect 23906 24871 23964 24877
rect 23906 24868 23918 24871
rect 23716 24840 23918 24868
rect 23716 24828 23722 24840
rect 23906 24837 23918 24840
rect 23952 24837 23964 24871
rect 23906 24831 23964 24837
rect 25869 24871 25927 24877
rect 25869 24837 25881 24871
rect 25915 24868 25927 24871
rect 26510 24868 26516 24880
rect 25915 24840 26516 24868
rect 25915 24837 25927 24840
rect 25869 24831 25927 24837
rect 26510 24828 26516 24840
rect 26568 24828 26574 24880
rect 22557 24803 22615 24809
rect 22557 24769 22569 24803
rect 22603 24769 22615 24803
rect 22557 24763 22615 24769
rect 22649 24803 22707 24809
rect 22649 24769 22661 24803
rect 22695 24800 22707 24803
rect 22738 24800 22744 24812
rect 22695 24772 22744 24800
rect 22695 24769 22707 24772
rect 22649 24763 22707 24769
rect 22738 24760 22744 24772
rect 22796 24760 22802 24812
rect 22833 24803 22891 24809
rect 22833 24769 22845 24803
rect 22879 24769 22891 24803
rect 22833 24763 22891 24769
rect 27792 24803 27850 24809
rect 27792 24769 27804 24803
rect 27838 24800 27850 24803
rect 28350 24800 28356 24812
rect 27838 24772 28356 24800
rect 27838 24769 27850 24772
rect 27792 24763 27850 24769
rect 19426 24732 19432 24744
rect 17828 24704 19432 24732
rect 17828 24692 17834 24704
rect 19426 24692 19432 24704
rect 19484 24692 19490 24744
rect 19797 24735 19855 24741
rect 19797 24701 19809 24735
rect 19843 24732 19855 24735
rect 21269 24735 21327 24741
rect 19843 24704 21128 24732
rect 19843 24701 19855 24704
rect 19797 24695 19855 24701
rect 15160 24636 15516 24664
rect 18233 24667 18291 24673
rect 15160 24624 15166 24636
rect 18233 24633 18245 24667
rect 18279 24664 18291 24667
rect 18414 24664 18420 24676
rect 18279 24636 18420 24664
rect 18279 24633 18291 24636
rect 18233 24627 18291 24633
rect 18414 24624 18420 24636
rect 18472 24624 18478 24676
rect 10689 24599 10747 24605
rect 10689 24565 10701 24599
rect 10735 24596 10747 24599
rect 11514 24596 11520 24608
rect 10735 24568 11520 24596
rect 10735 24565 10747 24568
rect 10689 24559 10747 24565
rect 11514 24556 11520 24568
rect 11572 24556 11578 24608
rect 11606 24556 11612 24608
rect 11664 24596 11670 24608
rect 11885 24599 11943 24605
rect 11885 24596 11897 24599
rect 11664 24568 11897 24596
rect 11664 24556 11670 24568
rect 11885 24565 11897 24568
rect 11931 24565 11943 24599
rect 11885 24559 11943 24565
rect 12802 24556 12808 24608
rect 12860 24596 12866 24608
rect 12897 24599 12955 24605
rect 12897 24596 12909 24599
rect 12860 24568 12909 24596
rect 12860 24556 12866 24568
rect 12897 24565 12909 24568
rect 12943 24565 12955 24599
rect 12897 24559 12955 24565
rect 14550 24556 14556 24608
rect 14608 24596 14614 24608
rect 17126 24596 17132 24608
rect 14608 24568 17132 24596
rect 14608 24556 14614 24568
rect 17126 24556 17132 24568
rect 17184 24556 17190 24608
rect 21100 24596 21128 24704
rect 21269 24701 21281 24735
rect 21315 24701 21327 24735
rect 22186 24732 22192 24744
rect 22147 24704 22192 24732
rect 21269 24695 21327 24701
rect 21284 24664 21312 24695
rect 22186 24692 22192 24704
rect 22244 24692 22250 24744
rect 22278 24692 22284 24744
rect 22336 24732 22342 24744
rect 22848 24732 22876 24763
rect 28350 24760 28356 24772
rect 28408 24760 28414 24812
rect 22336 24704 22876 24732
rect 23661 24735 23719 24741
rect 22336 24692 22342 24704
rect 23661 24701 23673 24735
rect 23707 24701 23719 24735
rect 25958 24732 25964 24744
rect 25919 24704 25964 24732
rect 23661 24695 23719 24701
rect 22646 24664 22652 24676
rect 21284 24636 22652 24664
rect 22646 24624 22652 24636
rect 22704 24624 22710 24676
rect 21542 24596 21548 24608
rect 21100 24568 21548 24596
rect 21542 24556 21548 24568
rect 21600 24556 21606 24608
rect 23676 24596 23704 24695
rect 25958 24692 25964 24704
rect 26016 24692 26022 24744
rect 26142 24732 26148 24744
rect 26103 24704 26148 24732
rect 26142 24692 26148 24704
rect 26200 24692 26206 24744
rect 27525 24735 27583 24741
rect 27525 24701 27537 24735
rect 27571 24701 27583 24735
rect 27525 24695 27583 24701
rect 26234 24664 26240 24676
rect 24596 24636 26240 24664
rect 24596 24596 24624 24636
rect 26234 24624 26240 24636
rect 26292 24664 26298 24676
rect 27430 24664 27436 24676
rect 26292 24636 27436 24664
rect 26292 24624 26298 24636
rect 27430 24624 27436 24636
rect 27488 24664 27494 24676
rect 27540 24664 27568 24695
rect 27488 24636 27568 24664
rect 27488 24624 27494 24636
rect 24670 24596 24676 24608
rect 23676 24568 24676 24596
rect 24670 24556 24676 24568
rect 24728 24556 24734 24608
rect 25038 24596 25044 24608
rect 24999 24568 25044 24596
rect 25038 24556 25044 24568
rect 25096 24556 25102 24608
rect 26970 24556 26976 24608
rect 27028 24596 27034 24608
rect 28905 24599 28963 24605
rect 28905 24596 28917 24599
rect 27028 24568 28917 24596
rect 27028 24556 27034 24568
rect 28905 24565 28917 24568
rect 28951 24565 28963 24599
rect 28905 24559 28963 24565
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 9214 24352 9220 24404
rect 9272 24392 9278 24404
rect 9585 24395 9643 24401
rect 9585 24392 9597 24395
rect 9272 24364 9597 24392
rect 9272 24352 9278 24364
rect 9585 24361 9597 24364
rect 9631 24361 9643 24395
rect 9585 24355 9643 24361
rect 10594 24352 10600 24404
rect 10652 24392 10658 24404
rect 10781 24395 10839 24401
rect 10781 24392 10793 24395
rect 10652 24364 10793 24392
rect 10652 24352 10658 24364
rect 10781 24361 10793 24364
rect 10827 24392 10839 24395
rect 10962 24392 10968 24404
rect 10827 24364 10968 24392
rect 10827 24361 10839 24364
rect 10781 24355 10839 24361
rect 10962 24352 10968 24364
rect 11020 24352 11026 24404
rect 12897 24395 12955 24401
rect 12897 24392 12909 24395
rect 12406 24364 12909 24392
rect 10226 24284 10232 24336
rect 10284 24324 10290 24336
rect 11790 24324 11796 24336
rect 10284 24296 11796 24324
rect 10284 24284 10290 24296
rect 11790 24284 11796 24296
rect 11848 24324 11854 24336
rect 12406 24324 12434 24364
rect 12897 24361 12909 24364
rect 12943 24361 12955 24395
rect 14274 24392 14280 24404
rect 14235 24364 14280 24392
rect 12897 24355 12955 24361
rect 14274 24352 14280 24364
rect 14332 24392 14338 24404
rect 15289 24395 15347 24401
rect 14332 24364 15240 24392
rect 14332 24352 14338 24364
rect 11848 24296 12434 24324
rect 11848 24284 11854 24296
rect 13170 24284 13176 24336
rect 13228 24324 13234 24336
rect 13630 24324 13636 24336
rect 13228 24296 13636 24324
rect 13228 24284 13234 24296
rect 13630 24284 13636 24296
rect 13688 24284 13694 24336
rect 15102 24324 15108 24336
rect 15063 24296 15108 24324
rect 15102 24284 15108 24296
rect 15160 24284 15166 24336
rect 15212 24324 15240 24364
rect 15289 24361 15301 24395
rect 15335 24392 15347 24395
rect 15378 24392 15384 24404
rect 15335 24364 15384 24392
rect 15335 24361 15347 24364
rect 15289 24355 15347 24361
rect 15378 24352 15384 24364
rect 15436 24352 15442 24404
rect 16114 24392 16120 24404
rect 15764 24364 16120 24392
rect 15764 24324 15792 24364
rect 16114 24352 16120 24364
rect 16172 24352 16178 24404
rect 16298 24352 16304 24404
rect 16356 24392 16362 24404
rect 16942 24392 16948 24404
rect 16356 24364 16948 24392
rect 16356 24352 16362 24364
rect 16942 24352 16948 24364
rect 17000 24352 17006 24404
rect 18046 24352 18052 24404
rect 18104 24392 18110 24404
rect 18506 24392 18512 24404
rect 18104 24364 18512 24392
rect 18104 24352 18110 24364
rect 18506 24352 18512 24364
rect 18564 24352 18570 24404
rect 18690 24352 18696 24404
rect 18748 24392 18754 24404
rect 19242 24392 19248 24404
rect 18748 24364 19248 24392
rect 18748 24352 18754 24364
rect 19242 24352 19248 24364
rect 19300 24392 19306 24404
rect 19705 24395 19763 24401
rect 19705 24392 19717 24395
rect 19300 24364 19717 24392
rect 19300 24352 19306 24364
rect 19705 24361 19717 24364
rect 19751 24361 19763 24395
rect 19705 24355 19763 24361
rect 19889 24395 19947 24401
rect 19889 24361 19901 24395
rect 19935 24392 19947 24395
rect 21082 24392 21088 24404
rect 19935 24364 21088 24392
rect 19935 24361 19947 24364
rect 19889 24355 19947 24361
rect 21082 24352 21088 24364
rect 21140 24352 21146 24404
rect 21266 24352 21272 24404
rect 21324 24392 21330 24404
rect 21453 24395 21511 24401
rect 21453 24392 21465 24395
rect 21324 24364 21465 24392
rect 21324 24352 21330 24364
rect 21453 24361 21465 24364
rect 21499 24361 21511 24395
rect 21453 24355 21511 24361
rect 22097 24395 22155 24401
rect 22097 24361 22109 24395
rect 22143 24392 22155 24395
rect 22278 24392 22284 24404
rect 22143 24364 22284 24392
rect 22143 24361 22155 24364
rect 22097 24355 22155 24361
rect 22278 24352 22284 24364
rect 22336 24352 22342 24404
rect 22554 24352 22560 24404
rect 22612 24392 22618 24404
rect 23109 24395 23167 24401
rect 23109 24392 23121 24395
rect 22612 24364 23121 24392
rect 22612 24352 22618 24364
rect 23109 24361 23121 24364
rect 23155 24361 23167 24395
rect 24486 24392 24492 24404
rect 23109 24355 23167 24361
rect 23584 24364 24492 24392
rect 15212 24296 15792 24324
rect 21637 24327 21695 24333
rect 21637 24293 21649 24327
rect 21683 24324 21695 24327
rect 21683 24296 22600 24324
rect 21683 24293 21695 24296
rect 21637 24287 21695 24293
rect 10410 24216 10416 24268
rect 10468 24256 10474 24268
rect 11514 24256 11520 24268
rect 10468 24228 10916 24256
rect 11475 24228 11520 24256
rect 10468 24216 10474 24228
rect 9493 24191 9551 24197
rect 9493 24157 9505 24191
rect 9539 24188 9551 24191
rect 9674 24188 9680 24200
rect 9539 24160 9680 24188
rect 9539 24157 9551 24160
rect 9493 24151 9551 24157
rect 9674 24148 9680 24160
rect 9732 24148 9738 24200
rect 10042 24148 10048 24200
rect 10100 24188 10106 24200
rect 10505 24191 10563 24197
rect 10505 24188 10517 24191
rect 10100 24160 10517 24188
rect 10100 24148 10106 24160
rect 10244 24052 10272 24160
rect 10505 24157 10517 24160
rect 10551 24157 10563 24191
rect 10505 24151 10563 24157
rect 10594 24148 10600 24200
rect 10652 24188 10658 24200
rect 10888 24197 10916 24228
rect 11514 24216 11520 24228
rect 11572 24216 11578 24268
rect 11606 24216 11612 24268
rect 11664 24256 11670 24268
rect 13081 24259 13139 24265
rect 11664 24228 11709 24256
rect 11664 24216 11670 24228
rect 13081 24225 13093 24259
rect 13127 24256 13139 24259
rect 13998 24256 14004 24268
rect 13127 24228 14004 24256
rect 13127 24225 13139 24228
rect 13081 24219 13139 24225
rect 13998 24216 14004 24228
rect 14056 24216 14062 24268
rect 17034 24256 17040 24268
rect 15948 24228 17040 24256
rect 10873 24191 10931 24197
rect 10652 24160 10697 24188
rect 10652 24148 10658 24160
rect 10873 24157 10885 24191
rect 10919 24157 10931 24191
rect 11698 24188 11704 24200
rect 10873 24151 10931 24157
rect 11256 24160 11704 24188
rect 10321 24123 10379 24129
rect 10321 24089 10333 24123
rect 10367 24120 10379 24123
rect 11256 24120 11284 24160
rect 11698 24148 11704 24160
rect 11756 24148 11762 24200
rect 12250 24188 12256 24200
rect 12211 24160 12256 24188
rect 12250 24148 12256 24160
rect 12308 24148 12314 24200
rect 12894 24188 12900 24200
rect 12855 24160 12900 24188
rect 12894 24148 12900 24160
rect 12952 24148 12958 24200
rect 13173 24191 13231 24197
rect 13173 24157 13185 24191
rect 13219 24188 13231 24191
rect 13219 24160 15700 24188
rect 13219 24157 13231 24160
rect 13173 24151 13231 24157
rect 14182 24120 14188 24132
rect 10367 24092 11284 24120
rect 14143 24092 14188 24120
rect 10367 24089 10379 24092
rect 10321 24083 10379 24089
rect 14182 24080 14188 24092
rect 14240 24080 14246 24132
rect 14826 24120 14832 24132
rect 14787 24092 14832 24120
rect 14826 24080 14832 24092
rect 14884 24080 14890 24132
rect 14918 24080 14924 24132
rect 14976 24120 14982 24132
rect 15378 24120 15384 24132
rect 14976 24092 15384 24120
rect 14976 24080 14982 24092
rect 15378 24080 15384 24092
rect 15436 24080 15442 24132
rect 10594 24052 10600 24064
rect 10244 24024 10600 24052
rect 10594 24012 10600 24024
rect 10652 24012 10658 24064
rect 11333 24055 11391 24061
rect 11333 24021 11345 24055
rect 11379 24052 11391 24055
rect 11882 24052 11888 24064
rect 11379 24024 11888 24052
rect 11379 24021 11391 24024
rect 11333 24015 11391 24021
rect 11882 24012 11888 24024
rect 11940 24012 11946 24064
rect 12342 24052 12348 24064
rect 12303 24024 12348 24052
rect 12342 24012 12348 24024
rect 12400 24012 12406 24064
rect 13354 24052 13360 24064
rect 13315 24024 13360 24052
rect 13354 24012 13360 24024
rect 13412 24012 13418 24064
rect 15672 24052 15700 24160
rect 15746 24148 15752 24200
rect 15804 24188 15810 24200
rect 15948 24197 15976 24228
rect 17034 24216 17040 24228
rect 17092 24216 17098 24268
rect 17218 24216 17224 24268
rect 17276 24256 17282 24268
rect 17497 24259 17555 24265
rect 17497 24256 17509 24259
rect 17276 24228 17509 24256
rect 17276 24216 17282 24228
rect 17497 24225 17509 24228
rect 17543 24225 17555 24259
rect 17770 24256 17776 24268
rect 17731 24228 17776 24256
rect 17497 24219 17555 24225
rect 17770 24216 17776 24228
rect 17828 24216 17834 24268
rect 20070 24256 20076 24268
rect 17880 24228 20076 24256
rect 15933 24191 15991 24197
rect 15804 24160 15849 24188
rect 15804 24148 15810 24160
rect 15933 24157 15945 24191
rect 15979 24157 15991 24191
rect 16114 24188 16120 24200
rect 16075 24160 16120 24188
rect 15933 24151 15991 24157
rect 16114 24148 16120 24160
rect 16172 24148 16178 24200
rect 16761 24191 16819 24197
rect 16761 24157 16773 24191
rect 16807 24188 16819 24191
rect 16942 24188 16948 24200
rect 16807 24160 16948 24188
rect 16807 24157 16819 24160
rect 16761 24151 16819 24157
rect 16942 24148 16948 24160
rect 17000 24148 17006 24200
rect 16022 24120 16028 24132
rect 15983 24092 16028 24120
rect 16022 24080 16028 24092
rect 16080 24080 16086 24132
rect 17880 24120 17908 24228
rect 20070 24216 20076 24228
rect 20128 24216 20134 24268
rect 21284 24228 21588 24256
rect 18782 24148 18788 24200
rect 18840 24188 18846 24200
rect 20349 24191 20407 24197
rect 20349 24188 20361 24191
rect 18840 24160 20361 24188
rect 18840 24148 18846 24160
rect 20349 24157 20361 24160
rect 20395 24157 20407 24191
rect 20349 24151 20407 24157
rect 16132 24092 17908 24120
rect 16132 24052 16160 24092
rect 19426 24080 19432 24132
rect 19484 24120 19490 24132
rect 21284 24129 21312 24228
rect 21560 24188 21588 24228
rect 22278 24188 22284 24200
rect 21560 24160 22094 24188
rect 22239 24160 22284 24188
rect 19521 24123 19579 24129
rect 19521 24120 19533 24123
rect 19484 24092 19533 24120
rect 19484 24080 19490 24092
rect 19521 24089 19533 24092
rect 19567 24089 19579 24123
rect 19521 24083 19579 24089
rect 19737 24123 19795 24129
rect 19737 24089 19749 24123
rect 19783 24120 19795 24123
rect 21269 24123 21327 24129
rect 19783 24092 21128 24120
rect 19783 24089 19795 24092
rect 19737 24083 19795 24089
rect 15672 24024 16160 24052
rect 16301 24055 16359 24061
rect 16301 24021 16313 24055
rect 16347 24052 16359 24055
rect 16390 24052 16396 24064
rect 16347 24024 16396 24052
rect 16347 24021 16359 24024
rect 16301 24015 16359 24021
rect 16390 24012 16396 24024
rect 16448 24012 16454 24064
rect 16850 24012 16856 24064
rect 16908 24052 16914 24064
rect 17126 24052 17132 24064
rect 16908 24024 17132 24052
rect 16908 24012 16914 24024
rect 17126 24012 17132 24024
rect 17184 24012 17190 24064
rect 19978 24012 19984 24064
rect 20036 24052 20042 24064
rect 20533 24055 20591 24061
rect 20533 24052 20545 24055
rect 20036 24024 20545 24052
rect 20036 24012 20042 24024
rect 20533 24021 20545 24024
rect 20579 24052 20591 24055
rect 20622 24052 20628 24064
rect 20579 24024 20628 24052
rect 20579 24021 20591 24024
rect 20533 24015 20591 24021
rect 20622 24012 20628 24024
rect 20680 24012 20686 24064
rect 21100 24052 21128 24092
rect 21269 24089 21281 24123
rect 21315 24089 21327 24123
rect 22066 24120 22094 24160
rect 22278 24148 22284 24160
rect 22336 24148 22342 24200
rect 22373 24191 22431 24197
rect 22373 24157 22385 24191
rect 22419 24188 22431 24191
rect 22462 24188 22468 24200
rect 22419 24160 22468 24188
rect 22419 24157 22431 24160
rect 22373 24151 22431 24157
rect 22462 24148 22468 24160
rect 22520 24148 22526 24200
rect 22572 24197 22600 24296
rect 23584 24265 23612 24364
rect 24486 24352 24492 24364
rect 24544 24392 24550 24404
rect 26053 24395 26111 24401
rect 26053 24392 26065 24395
rect 24544 24364 26065 24392
rect 24544 24352 24550 24364
rect 26053 24361 26065 24364
rect 26099 24361 26111 24395
rect 26510 24392 26516 24404
rect 26471 24364 26516 24392
rect 26053 24355 26111 24361
rect 26510 24352 26516 24364
rect 26568 24352 26574 24404
rect 28350 24352 28356 24404
rect 28408 24392 28414 24404
rect 28445 24395 28503 24401
rect 28445 24392 28457 24395
rect 28408 24364 28457 24392
rect 28408 24352 28414 24364
rect 28445 24361 28457 24364
rect 28491 24361 28503 24395
rect 28445 24355 28503 24361
rect 23569 24259 23627 24265
rect 23569 24225 23581 24259
rect 23615 24225 23627 24259
rect 23569 24219 23627 24225
rect 23753 24259 23811 24265
rect 23753 24225 23765 24259
rect 23799 24225 23811 24259
rect 24670 24256 24676 24268
rect 24631 24228 24676 24256
rect 23753 24219 23811 24225
rect 22557 24191 22615 24197
rect 22557 24157 22569 24191
rect 22603 24157 22615 24191
rect 22557 24151 22615 24157
rect 22646 24148 22652 24200
rect 22704 24188 22710 24200
rect 22704 24160 22749 24188
rect 22704 24148 22710 24160
rect 23106 24148 23112 24200
rect 23164 24188 23170 24200
rect 23768 24188 23796 24219
rect 24670 24216 24676 24228
rect 24728 24216 24734 24268
rect 26970 24256 26976 24268
rect 26931 24228 26976 24256
rect 26970 24216 26976 24228
rect 27028 24216 27034 24268
rect 27154 24216 27160 24268
rect 27212 24256 27218 24268
rect 27985 24259 28043 24265
rect 27985 24256 27997 24259
rect 27212 24228 27997 24256
rect 27212 24216 27218 24228
rect 27985 24225 27997 24228
rect 28031 24225 28043 24259
rect 27985 24219 28043 24225
rect 27172 24188 27200 24216
rect 23164 24160 27200 24188
rect 23164 24148 23170 24160
rect 28534 24148 28540 24200
rect 28592 24188 28598 24200
rect 28629 24191 28687 24197
rect 28629 24188 28641 24191
rect 28592 24160 28641 24188
rect 28592 24148 28598 24160
rect 28629 24157 28641 24160
rect 28675 24157 28687 24191
rect 28629 24151 28687 24157
rect 22738 24120 22744 24132
rect 22066 24092 22744 24120
rect 21269 24083 21327 24089
rect 22738 24080 22744 24092
rect 22796 24080 22802 24132
rect 24946 24129 24952 24132
rect 24940 24083 24952 24129
rect 25004 24120 25010 24132
rect 25004 24092 25040 24120
rect 24946 24080 24952 24083
rect 25004 24080 25010 24092
rect 27338 24080 27344 24132
rect 27396 24120 27402 24132
rect 27801 24123 27859 24129
rect 27801 24120 27813 24123
rect 27396 24092 27813 24120
rect 27396 24080 27402 24092
rect 27801 24089 27813 24092
rect 27847 24089 27859 24123
rect 27801 24083 27859 24089
rect 21450 24052 21456 24064
rect 21508 24061 21514 24064
rect 21508 24055 21527 24061
rect 21100 24024 21456 24052
rect 21450 24012 21456 24024
rect 21515 24021 21527 24055
rect 21508 24015 21527 24021
rect 21508 24012 21514 24015
rect 22278 24012 22284 24064
rect 22336 24052 22342 24064
rect 23106 24052 23112 24064
rect 22336 24024 23112 24052
rect 22336 24012 22342 24024
rect 23106 24012 23112 24024
rect 23164 24012 23170 24064
rect 23474 24052 23480 24064
rect 23435 24024 23480 24052
rect 23474 24012 23480 24024
rect 23532 24012 23538 24064
rect 26050 24012 26056 24064
rect 26108 24052 26114 24064
rect 26881 24055 26939 24061
rect 26881 24052 26893 24055
rect 26108 24024 26893 24052
rect 26108 24012 26114 24024
rect 26881 24021 26893 24024
rect 26927 24021 26939 24055
rect 26881 24015 26939 24021
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 11882 23848 11888 23860
rect 10796 23820 11888 23848
rect 10502 23780 10508 23792
rect 7300 23752 10508 23780
rect 7006 23672 7012 23724
rect 7064 23712 7070 23724
rect 7300 23721 7328 23752
rect 10502 23740 10508 23752
rect 10560 23740 10566 23792
rect 7285 23715 7343 23721
rect 7285 23712 7297 23715
rect 7064 23684 7297 23712
rect 7064 23672 7070 23684
rect 7285 23681 7297 23684
rect 7331 23681 7343 23715
rect 7285 23675 7343 23681
rect 7552 23715 7610 23721
rect 7552 23681 7564 23715
rect 7598 23712 7610 23715
rect 8938 23712 8944 23724
rect 7598 23684 8944 23712
rect 7598 23681 7610 23684
rect 7552 23675 7610 23681
rect 8938 23672 8944 23684
rect 8996 23672 9002 23724
rect 9953 23715 10011 23721
rect 9953 23681 9965 23715
rect 9999 23712 10011 23715
rect 10134 23712 10140 23724
rect 9999 23684 10140 23712
rect 9999 23681 10011 23684
rect 9953 23675 10011 23681
rect 10134 23672 10140 23684
rect 10192 23672 10198 23724
rect 10597 23715 10655 23721
rect 10597 23681 10609 23715
rect 10643 23681 10655 23715
rect 10597 23675 10655 23681
rect 10689 23715 10747 23721
rect 10689 23681 10701 23715
rect 10735 23712 10747 23715
rect 10796 23712 10824 23820
rect 11882 23808 11888 23820
rect 11940 23808 11946 23860
rect 12526 23848 12532 23860
rect 12452 23820 12532 23848
rect 11609 23783 11667 23789
rect 11609 23780 11621 23783
rect 10980 23752 11621 23780
rect 10980 23721 11008 23752
rect 11609 23749 11621 23752
rect 11655 23749 11667 23783
rect 11609 23743 11667 23749
rect 10735 23684 10824 23712
rect 10873 23715 10931 23721
rect 10735 23681 10747 23684
rect 10689 23675 10747 23681
rect 10873 23681 10885 23715
rect 10919 23681 10931 23715
rect 10873 23675 10931 23681
rect 10965 23715 11023 23721
rect 10965 23681 10977 23715
rect 11011 23681 11023 23715
rect 11514 23712 11520 23724
rect 11475 23684 11520 23712
rect 10965 23675 11023 23681
rect 9490 23644 9496 23656
rect 8680 23616 9496 23644
rect 8680 23520 8708 23616
rect 9490 23604 9496 23616
rect 9548 23644 9554 23656
rect 9769 23647 9827 23653
rect 9769 23644 9781 23647
rect 9548 23616 9781 23644
rect 9548 23604 9554 23616
rect 9769 23613 9781 23616
rect 9815 23613 9827 23647
rect 9769 23607 9827 23613
rect 9585 23579 9643 23585
rect 9585 23545 9597 23579
rect 9631 23576 9643 23579
rect 9674 23576 9680 23588
rect 9631 23548 9680 23576
rect 9631 23545 9643 23548
rect 9585 23539 9643 23545
rect 9674 23536 9680 23548
rect 9732 23536 9738 23588
rect 10612 23576 10640 23675
rect 10888 23644 10916 23675
rect 11514 23672 11520 23684
rect 11572 23672 11578 23724
rect 11698 23712 11704 23724
rect 11659 23684 11704 23712
rect 11698 23672 11704 23684
rect 11756 23672 11762 23724
rect 12452 23721 12480 23820
rect 12526 23808 12532 23820
rect 12584 23808 12590 23860
rect 13170 23808 13176 23860
rect 13228 23848 13234 23860
rect 14829 23851 14887 23857
rect 13228 23820 13676 23848
rect 13228 23808 13234 23820
rect 13446 23780 13452 23792
rect 13407 23752 13452 23780
rect 13446 23740 13452 23752
rect 13504 23740 13510 23792
rect 13648 23743 13676 23820
rect 14829 23817 14841 23851
rect 14875 23848 14887 23851
rect 15102 23848 15108 23860
rect 14875 23820 15108 23848
rect 14875 23817 14887 23820
rect 14829 23811 14887 23817
rect 15102 23808 15108 23820
rect 15160 23808 15166 23860
rect 16850 23808 16856 23860
rect 16908 23848 16914 23860
rect 17037 23851 17095 23857
rect 17037 23848 17049 23851
rect 16908 23820 17049 23848
rect 16908 23808 16914 23820
rect 17037 23817 17049 23820
rect 17083 23817 17095 23851
rect 18322 23848 18328 23860
rect 17037 23811 17095 23817
rect 17135 23820 18328 23848
rect 13638 23737 13696 23743
rect 15194 23740 15200 23792
rect 15252 23780 15258 23792
rect 15470 23780 15476 23792
rect 15252 23752 15476 23780
rect 15252 23740 15258 23752
rect 15470 23740 15476 23752
rect 15528 23740 15534 23792
rect 15562 23740 15568 23792
rect 15620 23780 15626 23792
rect 15838 23780 15844 23792
rect 15620 23752 15844 23780
rect 15620 23740 15626 23752
rect 15838 23740 15844 23752
rect 15896 23780 15902 23792
rect 15933 23783 15991 23789
rect 15933 23780 15945 23783
rect 15896 23752 15945 23780
rect 15896 23740 15902 23752
rect 15933 23749 15945 23752
rect 15979 23780 15991 23783
rect 17135 23780 17163 23820
rect 18322 23808 18328 23820
rect 18380 23808 18386 23860
rect 18782 23808 18788 23860
rect 18840 23848 18846 23860
rect 19613 23851 19671 23857
rect 19613 23848 19625 23851
rect 18840 23820 19625 23848
rect 18840 23808 18846 23820
rect 19613 23817 19625 23820
rect 19659 23817 19671 23851
rect 21174 23848 21180 23860
rect 21135 23820 21180 23848
rect 19613 23811 19671 23817
rect 21174 23808 21180 23820
rect 21232 23808 21238 23860
rect 21358 23808 21364 23860
rect 21416 23848 21422 23860
rect 21821 23851 21879 23857
rect 21821 23848 21833 23851
rect 21416 23820 21833 23848
rect 21416 23808 21422 23820
rect 21821 23817 21833 23820
rect 21867 23817 21879 23851
rect 21821 23811 21879 23817
rect 23937 23851 23995 23857
rect 23937 23817 23949 23851
rect 23983 23848 23995 23851
rect 24578 23848 24584 23860
rect 23983 23820 24584 23848
rect 23983 23817 23995 23820
rect 23937 23811 23995 23817
rect 24578 23808 24584 23820
rect 24636 23808 24642 23860
rect 25682 23848 25688 23860
rect 25643 23820 25688 23848
rect 25682 23808 25688 23820
rect 25740 23808 25746 23860
rect 25958 23808 25964 23860
rect 26016 23848 26022 23860
rect 26973 23851 27031 23857
rect 26973 23848 26985 23851
rect 26016 23820 26985 23848
rect 26016 23808 26022 23820
rect 26973 23817 26985 23820
rect 27019 23817 27031 23851
rect 28534 23848 28540 23860
rect 28495 23820 28540 23848
rect 26973 23811 27031 23817
rect 28534 23808 28540 23820
rect 28592 23808 28598 23860
rect 15979 23752 17163 23780
rect 15979 23749 15991 23752
rect 15933 23743 15991 23749
rect 17678 23740 17684 23792
rect 17736 23780 17742 23792
rect 18478 23783 18536 23789
rect 18478 23780 18490 23783
rect 17736 23752 18490 23780
rect 17736 23740 17742 23752
rect 18478 23749 18490 23752
rect 18524 23749 18536 23783
rect 18478 23743 18536 23749
rect 23661 23783 23719 23789
rect 23661 23749 23673 23783
rect 23707 23780 23719 23783
rect 24302 23780 24308 23792
rect 23707 23752 24308 23780
rect 23707 23749 23719 23752
rect 23661 23743 23719 23749
rect 24302 23740 24308 23752
rect 24360 23740 24366 23792
rect 25038 23780 25044 23792
rect 24412 23752 25044 23780
rect 12437 23715 12495 23721
rect 12437 23681 12449 23715
rect 12483 23681 12495 23715
rect 12437 23675 12495 23681
rect 12529 23715 12587 23721
rect 12529 23681 12541 23715
rect 12575 23681 12587 23715
rect 12529 23675 12587 23681
rect 12621 23715 12679 23721
rect 12621 23681 12633 23715
rect 12667 23681 12679 23715
rect 12621 23675 12679 23681
rect 12781 23718 12839 23721
rect 12781 23715 12940 23718
rect 12781 23681 12793 23715
rect 12827 23712 12940 23715
rect 12986 23712 12992 23724
rect 12827 23690 12992 23712
rect 12827 23684 12848 23690
rect 12912 23684 12992 23690
rect 12827 23681 12839 23684
rect 12781 23675 12839 23681
rect 11330 23644 11336 23656
rect 10888 23616 11336 23644
rect 11330 23604 11336 23616
rect 11388 23604 11394 23656
rect 9784 23548 10640 23576
rect 9784 23520 9812 23548
rect 8662 23508 8668 23520
rect 8623 23480 8668 23508
rect 8662 23468 8668 23480
rect 8720 23468 8726 23520
rect 9766 23508 9772 23520
rect 9727 23480 9772 23508
rect 9766 23468 9772 23480
rect 9824 23468 9830 23520
rect 9861 23511 9919 23517
rect 9861 23477 9873 23511
rect 9907 23508 9919 23511
rect 9950 23508 9956 23520
rect 9907 23480 9956 23508
rect 9907 23477 9919 23480
rect 9861 23471 9919 23477
rect 9950 23468 9956 23480
rect 10008 23468 10014 23520
rect 10410 23508 10416 23520
rect 10371 23480 10416 23508
rect 10410 23468 10416 23480
rect 10468 23468 10474 23520
rect 11606 23468 11612 23520
rect 11664 23508 11670 23520
rect 12161 23511 12219 23517
rect 12161 23508 12173 23511
rect 11664 23480 12173 23508
rect 11664 23468 11670 23480
rect 12161 23477 12173 23480
rect 12207 23477 12219 23511
rect 12161 23471 12219 23477
rect 12434 23468 12440 23520
rect 12492 23508 12498 23520
rect 12544 23508 12572 23675
rect 12636 23644 12664 23675
rect 12986 23672 12992 23684
rect 13044 23672 13050 23724
rect 13078 23672 13084 23724
rect 13136 23712 13142 23724
rect 13265 23715 13323 23721
rect 13265 23712 13277 23715
rect 13136 23684 13277 23712
rect 13136 23672 13142 23684
rect 13265 23681 13277 23684
rect 13311 23681 13323 23715
rect 13538 23712 13544 23724
rect 13451 23684 13544 23712
rect 13265 23675 13323 23681
rect 13538 23672 13544 23684
rect 13596 23672 13602 23724
rect 13638 23703 13650 23737
rect 13684 23703 13696 23737
rect 14182 23712 14188 23724
rect 13638 23697 13696 23703
rect 14143 23684 14188 23712
rect 14182 23672 14188 23684
rect 14240 23672 14246 23724
rect 14369 23715 14427 23721
rect 14369 23681 14381 23715
rect 14415 23681 14427 23715
rect 14369 23675 14427 23681
rect 13357 23647 13415 23653
rect 13357 23644 13369 23647
rect 12636 23616 12756 23644
rect 12728 23588 12756 23616
rect 12820 23616 13369 23644
rect 12710 23536 12716 23588
rect 12768 23536 12774 23588
rect 12820 23508 12848 23616
rect 13357 23613 13369 23616
rect 13403 23613 13415 23647
rect 13357 23607 13415 23613
rect 13262 23536 13268 23588
rect 13320 23576 13326 23588
rect 13556 23576 13584 23672
rect 13320 23548 13584 23576
rect 13320 23536 13326 23548
rect 13814 23536 13820 23588
rect 13872 23576 13878 23588
rect 14384 23576 14412 23675
rect 14918 23672 14924 23724
rect 14976 23712 14982 23724
rect 15289 23715 15347 23721
rect 15289 23712 15301 23715
rect 14976 23684 15301 23712
rect 14976 23672 14982 23684
rect 15289 23681 15301 23684
rect 15335 23681 15347 23715
rect 15289 23675 15347 23681
rect 16114 23672 16120 23724
rect 16172 23712 16178 23724
rect 16482 23712 16488 23724
rect 16172 23684 16488 23712
rect 16172 23672 16178 23684
rect 16482 23672 16488 23684
rect 16540 23712 16546 23724
rect 18233 23715 18291 23721
rect 18233 23712 18245 23715
rect 16540 23684 18245 23712
rect 16540 23672 16546 23684
rect 18233 23681 18245 23684
rect 18279 23681 18291 23715
rect 18233 23675 18291 23681
rect 21085 23715 21143 23721
rect 21085 23681 21097 23715
rect 21131 23712 21143 23715
rect 21542 23712 21548 23724
rect 21131 23684 21548 23712
rect 21131 23681 21143 23684
rect 21085 23675 21143 23681
rect 21542 23672 21548 23684
rect 21600 23672 21606 23724
rect 22186 23712 22192 23724
rect 22147 23684 22192 23712
rect 22186 23672 22192 23684
rect 22244 23672 22250 23724
rect 22462 23672 22468 23724
rect 22520 23712 22526 23724
rect 23385 23715 23443 23721
rect 23385 23712 23397 23715
rect 22520 23684 23397 23712
rect 22520 23672 22526 23684
rect 23385 23681 23397 23684
rect 23431 23681 23443 23715
rect 23566 23712 23572 23724
rect 23527 23684 23572 23712
rect 23385 23675 23443 23681
rect 15010 23644 15016 23656
rect 14971 23616 15016 23644
rect 15010 23604 15016 23616
rect 15068 23604 15074 23656
rect 15105 23647 15163 23653
rect 15105 23613 15117 23647
rect 15151 23613 15163 23647
rect 15105 23607 15163 23613
rect 15197 23647 15255 23653
rect 15197 23613 15209 23647
rect 15243 23644 15255 23647
rect 15378 23644 15384 23656
rect 15243 23616 15384 23644
rect 15243 23613 15255 23616
rect 15197 23607 15255 23613
rect 13872 23548 14412 23576
rect 13872 23536 13878 23548
rect 12492 23480 12848 23508
rect 12492 23468 12498 23480
rect 13538 23468 13544 23520
rect 13596 23508 13602 23520
rect 14185 23511 14243 23517
rect 14185 23508 14197 23511
rect 13596 23480 14197 23508
rect 13596 23468 13602 23480
rect 14185 23477 14197 23480
rect 14231 23477 14243 23511
rect 14185 23471 14243 23477
rect 14274 23468 14280 23520
rect 14332 23508 14338 23520
rect 15120 23508 15148 23607
rect 15378 23604 15384 23616
rect 15436 23644 15442 23656
rect 15746 23644 15752 23656
rect 15436 23616 15752 23644
rect 15436 23604 15442 23616
rect 15746 23604 15752 23616
rect 15804 23644 15810 23656
rect 16853 23647 16911 23653
rect 15804 23616 16160 23644
rect 15804 23604 15810 23616
rect 16132 23585 16160 23616
rect 16853 23613 16865 23647
rect 16899 23644 16911 23647
rect 17126 23644 17132 23656
rect 16899 23616 17132 23644
rect 16899 23613 16911 23616
rect 16853 23607 16911 23613
rect 17126 23604 17132 23616
rect 17184 23604 17190 23656
rect 17221 23647 17279 23653
rect 17221 23613 17233 23647
rect 17267 23644 17279 23647
rect 17770 23644 17776 23656
rect 17267 23616 17776 23644
rect 17267 23613 17279 23616
rect 17221 23607 17279 23613
rect 17770 23604 17776 23616
rect 17828 23604 17834 23656
rect 22278 23644 22284 23656
rect 22239 23616 22284 23644
rect 22278 23604 22284 23616
rect 22336 23604 22342 23656
rect 22373 23647 22431 23653
rect 22373 23613 22385 23647
rect 22419 23644 22431 23647
rect 22646 23644 22652 23656
rect 22419 23616 22652 23644
rect 22419 23613 22431 23616
rect 22373 23607 22431 23613
rect 22646 23604 22652 23616
rect 22704 23604 22710 23656
rect 23400 23644 23428 23675
rect 23566 23672 23572 23684
rect 23624 23672 23630 23724
rect 23750 23712 23756 23724
rect 23711 23684 23756 23712
rect 23750 23672 23756 23684
rect 23808 23672 23814 23724
rect 24412 23712 24440 23752
rect 25038 23740 25044 23752
rect 25096 23740 25102 23792
rect 26145 23783 26203 23789
rect 26145 23749 26157 23783
rect 26191 23780 26203 23783
rect 26694 23780 26700 23792
rect 26191 23752 26700 23780
rect 26191 23749 26203 23752
rect 26145 23743 26203 23749
rect 26694 23740 26700 23752
rect 26752 23740 26758 23792
rect 27433 23783 27491 23789
rect 27433 23749 27445 23783
rect 27479 23780 27491 23783
rect 27522 23780 27528 23792
rect 27479 23752 27528 23780
rect 27479 23749 27491 23752
rect 27433 23743 27491 23749
rect 27522 23740 27528 23752
rect 27580 23740 27586 23792
rect 23860 23684 24440 23712
rect 24581 23715 24639 23721
rect 23860 23644 23888 23684
rect 24581 23681 24593 23715
rect 24627 23712 24639 23715
rect 24946 23712 24952 23724
rect 24627 23684 24952 23712
rect 24627 23681 24639 23684
rect 24581 23675 24639 23681
rect 24946 23672 24952 23684
rect 25004 23672 25010 23724
rect 26053 23715 26111 23721
rect 26053 23681 26065 23715
rect 26099 23712 26111 23715
rect 27062 23712 27068 23724
rect 26099 23684 27068 23712
rect 26099 23681 26111 23684
rect 26053 23675 26111 23681
rect 27062 23672 27068 23684
rect 27120 23672 27126 23724
rect 27246 23672 27252 23724
rect 27304 23712 27310 23724
rect 27341 23715 27399 23721
rect 27341 23712 27353 23715
rect 27304 23684 27353 23712
rect 27304 23672 27310 23684
rect 27341 23681 27353 23684
rect 27387 23681 27399 23715
rect 28350 23712 28356 23724
rect 28311 23684 28356 23712
rect 27341 23675 27399 23681
rect 28350 23672 28356 23684
rect 28408 23672 28414 23724
rect 29178 23712 29184 23724
rect 29139 23684 29184 23712
rect 29178 23672 29184 23684
rect 29236 23672 29242 23724
rect 29825 23715 29883 23721
rect 29825 23681 29837 23715
rect 29871 23712 29883 23715
rect 29914 23712 29920 23724
rect 29871 23684 29920 23712
rect 29871 23681 29883 23684
rect 29825 23675 29883 23681
rect 29914 23672 29920 23684
rect 29972 23672 29978 23724
rect 23400 23616 23888 23644
rect 23934 23604 23940 23656
rect 23992 23644 23998 23656
rect 24394 23644 24400 23656
rect 23992 23616 24400 23644
rect 23992 23604 23998 23616
rect 24394 23604 24400 23616
rect 24452 23604 24458 23656
rect 26329 23647 26387 23653
rect 26329 23613 26341 23647
rect 26375 23644 26387 23647
rect 27154 23644 27160 23656
rect 26375 23616 27160 23644
rect 26375 23613 26387 23616
rect 26329 23607 26387 23613
rect 27154 23604 27160 23616
rect 27212 23604 27218 23656
rect 27525 23647 27583 23653
rect 27525 23613 27537 23647
rect 27571 23613 27583 23647
rect 27525 23607 27583 23613
rect 28169 23647 28227 23653
rect 28169 23613 28181 23647
rect 28215 23644 28227 23647
rect 28258 23644 28264 23656
rect 28215 23616 28264 23644
rect 28215 23613 28227 23616
rect 28169 23607 28227 23613
rect 16117 23579 16175 23585
rect 16117 23545 16129 23579
rect 16163 23545 16175 23579
rect 16117 23539 16175 23545
rect 26418 23536 26424 23588
rect 26476 23576 26482 23588
rect 27338 23576 27344 23588
rect 26476 23548 27344 23576
rect 26476 23536 26482 23548
rect 27338 23536 27344 23548
rect 27396 23576 27402 23588
rect 27540 23576 27568 23607
rect 28258 23604 28264 23616
rect 28316 23604 28322 23656
rect 27396 23548 27568 23576
rect 27396 23536 27402 23548
rect 15470 23508 15476 23520
rect 14332 23480 15476 23508
rect 14332 23468 14338 23480
rect 15470 23468 15476 23480
rect 15528 23468 15534 23520
rect 16942 23468 16948 23520
rect 17000 23508 17006 23520
rect 17221 23511 17279 23517
rect 17221 23508 17233 23511
rect 17000 23480 17233 23508
rect 17000 23468 17006 23480
rect 17221 23477 17233 23480
rect 17267 23477 17279 23511
rect 17221 23471 17279 23477
rect 24026 23468 24032 23520
rect 24084 23508 24090 23520
rect 24765 23511 24823 23517
rect 24765 23508 24777 23511
rect 24084 23480 24777 23508
rect 24084 23468 24090 23480
rect 24765 23477 24777 23480
rect 24811 23477 24823 23511
rect 28994 23508 29000 23520
rect 28955 23480 29000 23508
rect 24765 23471 24823 23477
rect 28994 23468 29000 23480
rect 29052 23468 29058 23520
rect 29638 23508 29644 23520
rect 29599 23480 29644 23508
rect 29638 23468 29644 23480
rect 29696 23468 29702 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 8110 23264 8116 23316
rect 8168 23304 8174 23316
rect 8297 23307 8355 23313
rect 8297 23304 8309 23307
rect 8168 23276 8309 23304
rect 8168 23264 8174 23276
rect 8297 23273 8309 23276
rect 8343 23273 8355 23307
rect 8938 23304 8944 23316
rect 8899 23276 8944 23304
rect 8297 23267 8355 23273
rect 8312 23236 8340 23267
rect 8938 23264 8944 23276
rect 8996 23264 9002 23316
rect 9398 23264 9404 23316
rect 9456 23304 9462 23316
rect 11146 23304 11152 23316
rect 9456 23276 11152 23304
rect 9456 23264 9462 23276
rect 11146 23264 11152 23276
rect 11204 23264 11210 23316
rect 11330 23304 11336 23316
rect 11291 23276 11336 23304
rect 11330 23264 11336 23276
rect 11388 23264 11394 23316
rect 12526 23264 12532 23316
rect 12584 23304 12590 23316
rect 12989 23307 13047 23313
rect 12989 23304 13001 23307
rect 12584 23276 13001 23304
rect 12584 23264 12590 23276
rect 12989 23273 13001 23276
rect 13035 23304 13047 23307
rect 14093 23307 14151 23313
rect 14093 23304 14105 23307
rect 13035 23276 14105 23304
rect 13035 23273 13047 23276
rect 12989 23267 13047 23273
rect 14093 23273 14105 23276
rect 14139 23273 14151 23307
rect 14093 23267 14151 23273
rect 14737 23307 14795 23313
rect 14737 23273 14749 23307
rect 14783 23304 14795 23307
rect 14826 23304 14832 23316
rect 14783 23276 14832 23304
rect 14783 23273 14795 23276
rect 14737 23267 14795 23273
rect 14826 23264 14832 23276
rect 14884 23264 14890 23316
rect 15654 23304 15660 23316
rect 15028 23276 15660 23304
rect 9214 23236 9220 23248
rect 8312 23208 9220 23236
rect 9214 23196 9220 23208
rect 9272 23196 9278 23248
rect 10045 23239 10103 23245
rect 10045 23205 10057 23239
rect 10091 23236 10103 23239
rect 11514 23236 11520 23248
rect 10091 23208 11520 23236
rect 10091 23205 10103 23208
rect 10045 23199 10103 23205
rect 11514 23196 11520 23208
rect 11572 23236 11578 23248
rect 11572 23208 12020 23236
rect 11572 23196 11578 23208
rect 8938 23128 8944 23180
rect 8996 23168 9002 23180
rect 9122 23168 9128 23180
rect 8996 23140 9128 23168
rect 8996 23128 9002 23140
rect 9122 23128 9128 23140
rect 9180 23168 9186 23180
rect 9180 23140 9352 23168
rect 9180 23128 9186 23140
rect 8662 23060 8668 23112
rect 8720 23100 8726 23112
rect 9324 23109 9352 23140
rect 9490 23128 9496 23180
rect 9548 23168 9554 23180
rect 9548 23140 10272 23168
rect 9548 23128 9554 23140
rect 9217 23103 9275 23109
rect 9217 23100 9229 23103
rect 8720 23072 9229 23100
rect 8720 23060 8726 23072
rect 9217 23069 9229 23072
rect 9263 23069 9275 23103
rect 9217 23063 9275 23069
rect 9309 23103 9367 23109
rect 9309 23069 9321 23103
rect 9355 23069 9367 23103
rect 9309 23063 9367 23069
rect 9398 23060 9404 23112
rect 9456 23100 9462 23112
rect 9456 23072 9501 23100
rect 9456 23060 9462 23072
rect 9582 23060 9588 23112
rect 9640 23100 9646 23112
rect 9640 23072 9685 23100
rect 9640 23060 9646 23072
rect 9766 23060 9772 23112
rect 9824 23100 9830 23112
rect 10244 23109 10272 23140
rect 10045 23103 10103 23109
rect 10045 23100 10057 23103
rect 9824 23072 10057 23100
rect 9824 23060 9830 23072
rect 10045 23069 10057 23072
rect 10091 23069 10103 23103
rect 10045 23063 10103 23069
rect 10229 23103 10287 23109
rect 10229 23069 10241 23103
rect 10275 23069 10287 23103
rect 10229 23063 10287 23069
rect 10321 23103 10379 23109
rect 10321 23069 10333 23103
rect 10367 23069 10379 23103
rect 11606 23100 11612 23112
rect 11567 23072 11612 23100
rect 10321 23063 10379 23069
rect 8205 23035 8263 23041
rect 8205 23001 8217 23035
rect 8251 23032 8263 23035
rect 8846 23032 8852 23044
rect 8251 23004 8852 23032
rect 8251 23001 8263 23004
rect 8205 22995 8263 23001
rect 8680 22976 8708 23004
rect 8846 22992 8852 23004
rect 8904 22992 8910 23044
rect 9030 22992 9036 23044
rect 9088 23032 9094 23044
rect 9600 23032 9628 23060
rect 10336 23032 10364 23063
rect 11606 23060 11612 23072
rect 11664 23060 11670 23112
rect 11701 23103 11759 23109
rect 11701 23069 11713 23103
rect 11747 23069 11759 23103
rect 11701 23063 11759 23069
rect 11793 23103 11851 23109
rect 11793 23069 11805 23103
rect 11839 23100 11851 23103
rect 11882 23100 11888 23112
rect 11839 23072 11888 23100
rect 11839 23069 11851 23072
rect 11793 23063 11851 23069
rect 9088 23004 9628 23032
rect 9784 23004 10364 23032
rect 9088 22992 9094 23004
rect 9784 22976 9812 23004
rect 8662 22924 8668 22976
rect 8720 22924 8726 22976
rect 9306 22924 9312 22976
rect 9364 22964 9370 22976
rect 9582 22964 9588 22976
rect 9364 22936 9588 22964
rect 9364 22924 9370 22936
rect 9582 22924 9588 22936
rect 9640 22924 9646 22976
rect 9766 22924 9772 22976
rect 9824 22924 9830 22976
rect 11716 22964 11744 23063
rect 11882 23060 11888 23072
rect 11940 23060 11946 23112
rect 11992 23109 12020 23208
rect 12250 23196 12256 23248
rect 12308 23236 12314 23248
rect 12618 23236 12624 23248
rect 12308 23208 12624 23236
rect 12308 23196 12314 23208
rect 12618 23196 12624 23208
rect 12676 23196 12682 23248
rect 13173 23239 13231 23245
rect 13173 23205 13185 23239
rect 13219 23236 13231 23239
rect 13906 23236 13912 23248
rect 13219 23208 13912 23236
rect 13219 23205 13231 23208
rect 13173 23199 13231 23205
rect 13906 23196 13912 23208
rect 13964 23196 13970 23248
rect 15028 23236 15056 23276
rect 15654 23264 15660 23276
rect 15712 23304 15718 23316
rect 16298 23304 16304 23316
rect 15712 23276 16304 23304
rect 15712 23264 15718 23276
rect 16298 23264 16304 23276
rect 16356 23264 16362 23316
rect 17218 23264 17224 23316
rect 17276 23304 17282 23316
rect 17497 23307 17555 23313
rect 17497 23304 17509 23307
rect 17276 23276 17509 23304
rect 17276 23264 17282 23276
rect 17497 23273 17509 23276
rect 17543 23273 17555 23307
rect 17497 23267 17555 23273
rect 18233 23307 18291 23313
rect 18233 23273 18245 23307
rect 18279 23304 18291 23307
rect 20070 23304 20076 23316
rect 18279 23276 20076 23304
rect 18279 23273 18291 23276
rect 18233 23267 18291 23273
rect 14936 23208 15056 23236
rect 12434 23128 12440 23180
rect 12492 23168 12498 23180
rect 14936 23177 14964 23208
rect 12529 23171 12587 23177
rect 12529 23168 12541 23171
rect 12492 23140 12541 23168
rect 12492 23128 12498 23140
rect 12529 23137 12541 23140
rect 12575 23137 12587 23171
rect 12529 23131 12587 23137
rect 14921 23171 14979 23177
rect 14921 23137 14933 23171
rect 14967 23137 14979 23171
rect 14921 23131 14979 23137
rect 15013 23171 15071 23177
rect 15013 23137 15025 23171
rect 15059 23168 15071 23171
rect 15562 23168 15568 23180
rect 15059 23140 15568 23168
rect 15059 23137 15071 23140
rect 15013 23131 15071 23137
rect 15562 23128 15568 23140
rect 15620 23128 15626 23180
rect 16114 23168 16120 23180
rect 16075 23140 16120 23168
rect 16114 23128 16120 23140
rect 16172 23128 16178 23180
rect 17512 23168 17540 23267
rect 20070 23264 20076 23276
rect 20128 23264 20134 23316
rect 22186 23264 22192 23316
rect 22244 23304 22250 23316
rect 22465 23307 22523 23313
rect 22465 23304 22477 23307
rect 22244 23276 22477 23304
rect 22244 23264 22250 23276
rect 22465 23273 22477 23276
rect 22511 23273 22523 23307
rect 22465 23267 22523 23273
rect 23290 23264 23296 23316
rect 23348 23304 23354 23316
rect 23348 23276 24900 23304
rect 23348 23264 23354 23276
rect 23661 23239 23719 23245
rect 23661 23205 23673 23239
rect 23707 23236 23719 23239
rect 24762 23236 24768 23248
rect 23707 23208 24768 23236
rect 23707 23205 23719 23208
rect 23661 23199 23719 23205
rect 24762 23196 24768 23208
rect 24820 23196 24826 23248
rect 23106 23168 23112 23180
rect 17512 23140 18092 23168
rect 23067 23140 23112 23168
rect 11977 23103 12035 23109
rect 11977 23069 11989 23103
rect 12023 23069 12035 23103
rect 11977 23063 12035 23069
rect 12618 23060 12624 23112
rect 12676 23100 12682 23112
rect 12676 23072 12721 23100
rect 12676 23060 12682 23072
rect 12894 23060 12900 23112
rect 12952 23100 12958 23112
rect 12989 23103 13047 23109
rect 12989 23100 13001 23103
rect 12952 23072 13001 23100
rect 12952 23060 12958 23072
rect 12989 23069 13001 23072
rect 13035 23069 13047 23103
rect 12989 23063 13047 23069
rect 13170 23060 13176 23112
rect 13228 23100 13234 23112
rect 14093 23103 14151 23109
rect 14093 23100 14105 23103
rect 13228 23072 14105 23100
rect 13228 23060 13234 23072
rect 14093 23069 14105 23072
rect 14139 23069 14151 23103
rect 14093 23063 14151 23069
rect 14277 23103 14335 23109
rect 14277 23069 14289 23103
rect 14323 23069 14335 23103
rect 14277 23063 14335 23069
rect 12526 22992 12532 23044
rect 12584 23032 12590 23044
rect 13188 23032 13216 23060
rect 12584 23004 13216 23032
rect 12584 22992 12590 23004
rect 13262 22992 13268 23044
rect 13320 23032 13326 23044
rect 14292 23032 14320 23063
rect 15102 23060 15108 23112
rect 15160 23100 15166 23112
rect 16390 23109 16396 23112
rect 15381 23103 15439 23109
rect 15381 23100 15393 23103
rect 15160 23072 15393 23100
rect 15160 23060 15166 23072
rect 15381 23069 15393 23072
rect 15427 23069 15439 23103
rect 16384 23100 16396 23109
rect 16351 23072 16396 23100
rect 15381 23063 15439 23069
rect 16384 23063 16396 23072
rect 16390 23060 16396 23063
rect 16448 23060 16454 23112
rect 16850 23060 16856 23112
rect 16908 23100 16914 23112
rect 17770 23100 17776 23112
rect 16908 23072 17776 23100
rect 16908 23060 16914 23072
rect 17770 23060 17776 23072
rect 17828 23100 17834 23112
rect 18064 23109 18092 23140
rect 23106 23128 23112 23140
rect 23164 23128 23170 23180
rect 23750 23128 23756 23180
rect 23808 23168 23814 23180
rect 24872 23168 24900 23276
rect 24946 23264 24952 23316
rect 25004 23304 25010 23316
rect 27341 23307 27399 23313
rect 25004 23276 25049 23304
rect 25004 23264 25010 23276
rect 27341 23273 27353 23307
rect 27387 23304 27399 23307
rect 28350 23304 28356 23316
rect 27387 23276 28356 23304
rect 27387 23273 27399 23276
rect 27341 23267 27399 23273
rect 28350 23264 28356 23276
rect 28408 23264 28414 23316
rect 28629 23307 28687 23313
rect 28629 23273 28641 23307
rect 28675 23304 28687 23307
rect 29178 23304 29184 23316
rect 28675 23276 29184 23304
rect 28675 23273 28687 23276
rect 28629 23267 28687 23273
rect 29178 23264 29184 23276
rect 29236 23264 29242 23316
rect 26418 23168 26424 23180
rect 23808 23140 24808 23168
rect 24872 23140 26424 23168
rect 23808 23128 23814 23140
rect 17957 23103 18015 23109
rect 17957 23100 17969 23103
rect 17828 23072 17969 23100
rect 17828 23060 17834 23072
rect 17957 23069 17969 23072
rect 18003 23069 18015 23103
rect 17957 23063 18015 23069
rect 18049 23103 18107 23109
rect 18049 23069 18061 23103
rect 18095 23069 18107 23103
rect 18322 23100 18328 23112
rect 18283 23072 18328 23100
rect 18049 23063 18107 23069
rect 18322 23060 18328 23072
rect 18380 23060 18386 23112
rect 20625 23103 20683 23109
rect 20625 23069 20637 23103
rect 20671 23100 20683 23103
rect 21174 23100 21180 23112
rect 20671 23072 21180 23100
rect 20671 23069 20683 23072
rect 20625 23063 20683 23069
rect 21174 23060 21180 23072
rect 21232 23060 21238 23112
rect 23845 23103 23903 23109
rect 23845 23069 23857 23103
rect 23891 23100 23903 23103
rect 24026 23100 24032 23112
rect 23891 23072 24032 23100
rect 23891 23069 23903 23072
rect 23845 23063 23903 23069
rect 24026 23060 24032 23072
rect 24084 23060 24090 23112
rect 24397 23103 24455 23109
rect 24397 23069 24409 23103
rect 24443 23100 24455 23103
rect 24486 23100 24492 23112
rect 24443 23072 24492 23100
rect 24443 23069 24455 23072
rect 24397 23063 24455 23069
rect 24486 23060 24492 23072
rect 24544 23060 24550 23112
rect 24780 23109 24808 23140
rect 26418 23128 26424 23140
rect 26476 23128 26482 23180
rect 26970 23168 26976 23180
rect 26804 23140 26976 23168
rect 24765 23103 24823 23109
rect 24765 23069 24777 23103
rect 24811 23069 24823 23103
rect 25590 23100 25596 23112
rect 25551 23072 25596 23100
rect 24765 23063 24823 23069
rect 25590 23060 25596 23072
rect 25648 23060 25654 23112
rect 26145 23103 26203 23109
rect 26145 23069 26157 23103
rect 26191 23100 26203 23103
rect 26234 23100 26240 23112
rect 26191 23072 26240 23100
rect 26191 23069 26203 23072
rect 26145 23063 26203 23069
rect 26234 23060 26240 23072
rect 26292 23060 26298 23112
rect 26804 23109 26832 23140
rect 26970 23128 26976 23140
rect 27028 23128 27034 23180
rect 27430 23128 27436 23180
rect 27488 23168 27494 23180
rect 29549 23171 29607 23177
rect 29549 23168 29561 23171
rect 27488 23140 29561 23168
rect 27488 23128 27494 23140
rect 29549 23137 29561 23140
rect 29595 23137 29607 23171
rect 29549 23131 29607 23137
rect 26789 23103 26847 23109
rect 26789 23069 26801 23103
rect 26835 23069 26847 23103
rect 26789 23063 26847 23069
rect 27157 23103 27215 23109
rect 27157 23069 27169 23103
rect 27203 23100 27215 23103
rect 28074 23100 28080 23112
rect 27203 23072 28080 23100
rect 27203 23069 27215 23072
rect 27157 23063 27215 23069
rect 28074 23060 28080 23072
rect 28132 23060 28138 23112
rect 28258 23100 28264 23112
rect 28219 23072 28264 23100
rect 28258 23060 28264 23072
rect 28316 23060 28322 23112
rect 28442 23100 28448 23112
rect 28403 23072 28448 23100
rect 28442 23060 28448 23072
rect 28500 23060 28506 23112
rect 28994 23060 29000 23112
rect 29052 23100 29058 23112
rect 29805 23103 29863 23109
rect 29805 23100 29817 23103
rect 29052 23072 29817 23100
rect 29052 23060 29058 23072
rect 29805 23069 29817 23072
rect 29851 23069 29863 23103
rect 29805 23063 29863 23069
rect 13320 23004 14320 23032
rect 16224 23004 18276 23032
rect 13320 22992 13326 23004
rect 11790 22964 11796 22976
rect 11716 22936 11796 22964
rect 11790 22924 11796 22936
rect 11848 22924 11854 22976
rect 12342 22924 12348 22976
rect 12400 22964 12406 22976
rect 12802 22964 12808 22976
rect 12400 22936 12808 22964
rect 12400 22924 12406 22936
rect 12802 22924 12808 22936
rect 12860 22964 12866 22976
rect 13998 22964 14004 22976
rect 12860 22936 14004 22964
rect 12860 22924 12866 22936
rect 13998 22924 14004 22936
rect 14056 22964 14062 22976
rect 14826 22964 14832 22976
rect 14056 22936 14832 22964
rect 14056 22924 14062 22936
rect 14826 22924 14832 22936
rect 14884 22924 14890 22976
rect 15010 22924 15016 22976
rect 15068 22964 15074 22976
rect 15105 22967 15163 22973
rect 15105 22964 15117 22967
rect 15068 22936 15117 22964
rect 15068 22924 15074 22936
rect 15105 22933 15117 22936
rect 15151 22933 15163 22967
rect 15105 22927 15163 22933
rect 15289 22967 15347 22973
rect 15289 22933 15301 22967
rect 15335 22964 15347 22967
rect 15470 22964 15476 22976
rect 15335 22936 15476 22964
rect 15335 22933 15347 22936
rect 15289 22927 15347 22933
rect 15470 22924 15476 22936
rect 15528 22924 15534 22976
rect 15562 22924 15568 22976
rect 15620 22964 15626 22976
rect 16224 22964 16252 23004
rect 15620 22936 16252 22964
rect 15620 22924 15626 22936
rect 17126 22924 17132 22976
rect 17184 22964 17190 22976
rect 17862 22964 17868 22976
rect 17184 22936 17868 22964
rect 17184 22924 17190 22936
rect 17862 22924 17868 22936
rect 17920 22964 17926 22976
rect 18141 22967 18199 22973
rect 18141 22964 18153 22967
rect 17920 22936 18153 22964
rect 17920 22924 17926 22936
rect 18141 22933 18153 22936
rect 18187 22933 18199 22967
rect 18248 22964 18276 23004
rect 20714 22992 20720 23044
rect 20772 23032 20778 23044
rect 20870 23035 20928 23041
rect 20870 23032 20882 23035
rect 20772 23004 20882 23032
rect 20772 22992 20778 23004
rect 20870 23001 20882 23004
rect 20916 23001 20928 23035
rect 20870 22995 20928 23001
rect 21082 22992 21088 23044
rect 21140 23032 21146 23044
rect 21910 23032 21916 23044
rect 21140 23004 21916 23032
rect 21140 22992 21146 23004
rect 21910 22992 21916 23004
rect 21968 22992 21974 23044
rect 23566 22992 23572 23044
rect 23624 23032 23630 23044
rect 24581 23035 24639 23041
rect 24581 23032 24593 23035
rect 23624 23004 24593 23032
rect 23624 22992 23630 23004
rect 24581 23001 24593 23004
rect 24627 23001 24639 23035
rect 24581 22995 24639 23001
rect 21358 22964 21364 22976
rect 18248 22936 21364 22964
rect 18141 22927 18199 22933
rect 21358 22924 21364 22936
rect 21416 22924 21422 22976
rect 22005 22967 22063 22973
rect 22005 22933 22017 22967
rect 22051 22964 22063 22967
rect 22094 22964 22100 22976
rect 22051 22936 22100 22964
rect 22051 22933 22063 22936
rect 22005 22927 22063 22933
rect 22094 22924 22100 22936
rect 22152 22924 22158 22976
rect 22554 22924 22560 22976
rect 22612 22964 22618 22976
rect 22833 22967 22891 22973
rect 22833 22964 22845 22967
rect 22612 22936 22845 22964
rect 22612 22924 22618 22936
rect 22833 22933 22845 22936
rect 22879 22933 22891 22967
rect 22833 22927 22891 22933
rect 22922 22924 22928 22976
rect 22980 22964 22986 22976
rect 24596 22964 24624 22995
rect 24670 22992 24676 23044
rect 24728 23032 24734 23044
rect 26973 23035 27031 23041
rect 24728 23004 24773 23032
rect 25240 23004 25544 23032
rect 24728 22992 24734 23004
rect 25240 22964 25268 23004
rect 25406 22964 25412 22976
rect 22980 22936 23025 22964
rect 24596 22936 25268 22964
rect 25367 22936 25412 22964
rect 22980 22924 22986 22936
rect 25406 22924 25412 22936
rect 25464 22924 25470 22976
rect 25516 22964 25544 23004
rect 26973 23001 26985 23035
rect 27019 23001 27031 23035
rect 26973 22995 27031 23001
rect 27065 23035 27123 23041
rect 27065 23001 27077 23035
rect 27111 23032 27123 23035
rect 27614 23032 27620 23044
rect 27111 23004 27620 23032
rect 27111 23001 27123 23004
rect 27065 22995 27123 23001
rect 26237 22967 26295 22973
rect 26237 22964 26249 22967
rect 25516 22936 26249 22964
rect 26237 22933 26249 22936
rect 26283 22964 26295 22967
rect 26418 22964 26424 22976
rect 26283 22936 26424 22964
rect 26283 22933 26295 22936
rect 26237 22927 26295 22933
rect 26418 22924 26424 22936
rect 26476 22964 26482 22976
rect 26988 22964 27016 22995
rect 27614 22992 27620 23004
rect 27672 22992 27678 23044
rect 26476 22936 27016 22964
rect 26476 22924 26482 22936
rect 27522 22924 27528 22976
rect 27580 22964 27586 22976
rect 30929 22967 30987 22973
rect 30929 22964 30941 22967
rect 27580 22936 30941 22964
rect 27580 22924 27586 22936
rect 30929 22933 30941 22936
rect 30975 22933 30987 22967
rect 30929 22927 30987 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 7101 22763 7159 22769
rect 7101 22729 7113 22763
rect 7147 22760 7159 22763
rect 9398 22760 9404 22772
rect 7147 22732 9404 22760
rect 7147 22729 7159 22732
rect 7101 22723 7159 22729
rect 9398 22720 9404 22732
rect 9456 22720 9462 22772
rect 10226 22760 10232 22772
rect 10187 22732 10232 22760
rect 10226 22720 10232 22732
rect 10284 22720 10290 22772
rect 10502 22720 10508 22772
rect 10560 22760 10566 22772
rect 10873 22763 10931 22769
rect 10873 22760 10885 22763
rect 10560 22732 10885 22760
rect 10560 22720 10566 22732
rect 10873 22729 10885 22732
rect 10919 22729 10931 22763
rect 10873 22723 10931 22729
rect 11146 22720 11152 22772
rect 11204 22760 11210 22772
rect 11701 22763 11759 22769
rect 11701 22760 11713 22763
rect 11204 22732 11713 22760
rect 11204 22720 11210 22732
rect 11701 22729 11713 22732
rect 11747 22729 11759 22763
rect 11701 22723 11759 22729
rect 12253 22763 12311 22769
rect 12253 22729 12265 22763
rect 12299 22760 12311 22763
rect 12618 22760 12624 22772
rect 12299 22732 12624 22760
rect 12299 22729 12311 22732
rect 12253 22723 12311 22729
rect 12618 22720 12624 22732
rect 12676 22720 12682 22772
rect 12710 22720 12716 22772
rect 12768 22760 12774 22772
rect 13725 22763 13783 22769
rect 12768 22732 12813 22760
rect 12768 22720 12774 22732
rect 13725 22729 13737 22763
rect 13771 22760 13783 22763
rect 13909 22763 13967 22769
rect 13771 22732 13860 22760
rect 13771 22729 13783 22732
rect 13725 22723 13783 22729
rect 8110 22692 8116 22704
rect 7116 22664 8116 22692
rect 6914 22624 6920 22636
rect 6875 22596 6920 22624
rect 6914 22584 6920 22596
rect 6972 22584 6978 22636
rect 7116 22633 7144 22664
rect 8110 22652 8116 22664
rect 8168 22652 8174 22704
rect 8570 22692 8576 22704
rect 8404 22664 8576 22692
rect 7101 22627 7159 22633
rect 7101 22593 7113 22627
rect 7147 22593 7159 22627
rect 7101 22587 7159 22593
rect 7561 22627 7619 22633
rect 7561 22593 7573 22627
rect 7607 22593 7619 22627
rect 8202 22624 8208 22636
rect 8163 22596 8208 22624
rect 7561 22587 7619 22593
rect 7576 22556 7604 22587
rect 8202 22584 8208 22596
rect 8260 22584 8266 22636
rect 8404 22633 8432 22664
rect 8570 22652 8576 22664
rect 8628 22692 8634 22704
rect 9309 22695 9367 22701
rect 9309 22692 9321 22695
rect 8628 22664 9321 22692
rect 8628 22652 8634 22664
rect 9309 22661 9321 22664
rect 9355 22661 9367 22695
rect 9309 22655 9367 22661
rect 10781 22695 10839 22701
rect 10781 22661 10793 22695
rect 10827 22692 10839 22695
rect 13078 22692 13084 22704
rect 10827 22664 13084 22692
rect 10827 22661 10839 22664
rect 10781 22655 10839 22661
rect 13078 22652 13084 22664
rect 13136 22652 13142 22704
rect 13633 22695 13691 22701
rect 13633 22692 13645 22695
rect 13188 22664 13645 22692
rect 8389 22627 8447 22633
rect 8389 22593 8401 22627
rect 8435 22593 8447 22627
rect 9122 22624 9128 22636
rect 9083 22596 9128 22624
rect 8389 22587 8447 22593
rect 9122 22584 9128 22596
rect 9180 22584 9186 22636
rect 9214 22584 9220 22636
rect 9272 22624 9278 22636
rect 9401 22627 9459 22633
rect 9401 22624 9413 22627
rect 9272 22596 9413 22624
rect 9272 22584 9278 22596
rect 9401 22593 9413 22596
rect 9447 22593 9459 22627
rect 9401 22587 9459 22593
rect 9861 22627 9919 22633
rect 9861 22593 9873 22627
rect 9907 22624 9919 22627
rect 10502 22624 10508 22636
rect 9907 22596 10508 22624
rect 9907 22593 9919 22596
rect 9861 22587 9919 22593
rect 10502 22584 10508 22596
rect 10560 22584 10566 22636
rect 11330 22584 11336 22636
rect 11388 22624 11394 22636
rect 11609 22627 11667 22633
rect 11609 22624 11621 22627
rect 11388 22596 11621 22624
rect 11388 22584 11394 22596
rect 11609 22593 11621 22596
rect 11655 22593 11667 22627
rect 11609 22587 11667 22593
rect 11974 22584 11980 22636
rect 12032 22624 12038 22636
rect 12529 22627 12587 22633
rect 12529 22624 12541 22627
rect 12032 22596 12541 22624
rect 12032 22584 12038 22596
rect 12529 22593 12541 22596
rect 12575 22593 12587 22627
rect 12529 22587 12587 22593
rect 12621 22627 12679 22633
rect 12621 22593 12633 22627
rect 12667 22624 12679 22627
rect 12802 22624 12808 22636
rect 12667 22596 12808 22624
rect 12667 22593 12679 22596
rect 12621 22587 12679 22593
rect 12802 22584 12808 22596
rect 12860 22584 12866 22636
rect 13188 22624 13216 22664
rect 13633 22661 13645 22664
rect 13679 22661 13691 22695
rect 13832 22692 13860 22732
rect 13909 22729 13921 22763
rect 13955 22760 13967 22763
rect 14274 22760 14280 22772
rect 13955 22732 14280 22760
rect 13955 22729 13967 22732
rect 13909 22723 13967 22729
rect 14274 22720 14280 22732
rect 14332 22720 14338 22772
rect 14369 22763 14427 22769
rect 14369 22729 14381 22763
rect 14415 22760 14427 22763
rect 15102 22760 15108 22772
rect 14415 22732 15108 22760
rect 14415 22729 14427 22732
rect 14369 22723 14427 22729
rect 15102 22720 15108 22732
rect 15160 22720 15166 22772
rect 15286 22720 15292 22772
rect 15344 22760 15350 22772
rect 15565 22763 15623 22769
rect 15565 22760 15577 22763
rect 15344 22732 15577 22760
rect 15344 22720 15350 22732
rect 15565 22729 15577 22732
rect 15611 22729 15623 22763
rect 16942 22760 16948 22772
rect 16903 22732 16948 22760
rect 15565 22723 15623 22729
rect 16942 22720 16948 22732
rect 17000 22720 17006 22772
rect 21821 22763 21879 22769
rect 21821 22729 21833 22763
rect 21867 22760 21879 22763
rect 22278 22760 22284 22772
rect 21867 22732 22284 22760
rect 21867 22729 21879 22732
rect 21821 22723 21879 22729
rect 22278 22720 22284 22732
rect 22336 22720 22342 22772
rect 22922 22720 22928 22772
rect 22980 22760 22986 22772
rect 25869 22763 25927 22769
rect 25869 22760 25881 22763
rect 22980 22732 25881 22760
rect 22980 22720 22986 22732
rect 14090 22692 14096 22704
rect 13832 22664 14096 22692
rect 13633 22655 13691 22661
rect 12912 22596 13216 22624
rect 13541 22627 13599 22633
rect 7576 22528 9444 22556
rect 7653 22491 7711 22497
rect 7653 22457 7665 22491
rect 7699 22488 7711 22491
rect 9306 22488 9312 22500
rect 7699 22460 9312 22488
rect 7699 22457 7711 22460
rect 7653 22451 7711 22457
rect 9306 22448 9312 22460
rect 9364 22448 9370 22500
rect 9416 22488 9444 22528
rect 9490 22516 9496 22568
rect 9548 22556 9554 22568
rect 9953 22559 10011 22565
rect 9953 22556 9965 22559
rect 9548 22528 9965 22556
rect 9548 22516 9554 22528
rect 9953 22525 9965 22528
rect 9999 22525 10011 22559
rect 9953 22519 10011 22525
rect 10410 22516 10416 22568
rect 10468 22556 10474 22568
rect 12912 22556 12940 22596
rect 13541 22593 13553 22627
rect 13587 22593 13599 22627
rect 13648 22624 13676 22655
rect 14090 22652 14096 22664
rect 14148 22692 14154 22704
rect 18322 22692 18328 22704
rect 14148 22664 14872 22692
rect 14148 22652 14154 22664
rect 14844 22633 14872 22664
rect 16960 22664 18328 22692
rect 14645 22630 14703 22633
rect 14476 22627 14703 22630
rect 14476 22624 14657 22627
rect 13648 22602 14657 22624
rect 13648 22596 14504 22602
rect 13541 22587 13599 22593
rect 14645 22593 14657 22602
rect 14691 22593 14703 22627
rect 14645 22587 14703 22593
rect 14829 22627 14887 22633
rect 14829 22593 14841 22627
rect 14875 22593 14887 22627
rect 14829 22587 14887 22593
rect 10468 22528 12940 22556
rect 12989 22559 13047 22565
rect 10468 22516 10474 22528
rect 12989 22525 13001 22559
rect 13035 22556 13047 22559
rect 13170 22556 13176 22568
rect 13035 22528 13176 22556
rect 13035 22525 13047 22528
rect 12989 22519 13047 22525
rect 13170 22516 13176 22528
rect 13228 22516 13234 22568
rect 13556 22556 13584 22587
rect 15102 22584 15108 22636
rect 15160 22624 15166 22636
rect 15378 22624 15384 22636
rect 15160 22596 15384 22624
rect 15160 22584 15166 22596
rect 15378 22584 15384 22596
rect 15436 22584 15442 22636
rect 15473 22627 15531 22633
rect 15473 22593 15485 22627
rect 15519 22624 15531 22627
rect 15562 22624 15568 22636
rect 15519 22596 15568 22624
rect 15519 22593 15531 22596
rect 15473 22587 15531 22593
rect 15562 22584 15568 22596
rect 15620 22584 15626 22636
rect 16761 22627 16819 22633
rect 16761 22593 16773 22627
rect 16807 22624 16819 22627
rect 16850 22624 16856 22636
rect 16807 22596 16856 22624
rect 16807 22593 16819 22596
rect 16761 22587 16819 22593
rect 16850 22584 16856 22596
rect 16908 22584 16914 22636
rect 16960 22633 16988 22664
rect 18322 22652 18328 22664
rect 18380 22652 18386 22704
rect 22094 22652 22100 22704
rect 22152 22692 22158 22704
rect 22152 22664 22324 22692
rect 22152 22652 22158 22664
rect 16945 22627 17003 22633
rect 16945 22593 16957 22627
rect 16991 22593 17003 22627
rect 16945 22587 17003 22593
rect 17034 22584 17040 22636
rect 17092 22624 17098 22636
rect 17586 22624 17592 22636
rect 17092 22596 17592 22624
rect 17092 22584 17098 22596
rect 17586 22584 17592 22596
rect 17644 22584 17650 22636
rect 17770 22584 17776 22636
rect 17828 22624 17834 22636
rect 18509 22627 18567 22633
rect 18509 22624 18521 22627
rect 17828 22596 18521 22624
rect 17828 22584 17834 22596
rect 18509 22593 18521 22596
rect 18555 22593 18567 22627
rect 18509 22587 18567 22593
rect 19337 22627 19395 22633
rect 19337 22593 19349 22627
rect 19383 22624 19395 22627
rect 22186 22624 22192 22636
rect 19383 22596 20392 22624
rect 22147 22596 22192 22624
rect 19383 22593 19395 22596
rect 19337 22587 19395 22593
rect 13909 22559 13967 22565
rect 13556 22528 13860 22556
rect 11054 22488 11060 22500
rect 9416 22460 11060 22488
rect 11054 22448 11060 22460
rect 11112 22448 11118 22500
rect 8294 22420 8300 22432
rect 8255 22392 8300 22420
rect 8294 22380 8300 22392
rect 8352 22380 8358 22432
rect 8386 22380 8392 22432
rect 8444 22420 8450 22432
rect 8573 22423 8631 22429
rect 8573 22420 8585 22423
rect 8444 22392 8585 22420
rect 8444 22380 8450 22392
rect 8573 22389 8585 22392
rect 8619 22389 8631 22423
rect 8573 22383 8631 22389
rect 8938 22380 8944 22432
rect 8996 22420 9002 22432
rect 9214 22420 9220 22432
rect 8996 22392 9220 22420
rect 8996 22380 9002 22392
rect 9214 22380 9220 22392
rect 9272 22380 9278 22432
rect 9398 22420 9404 22432
rect 9359 22392 9404 22420
rect 9398 22380 9404 22392
rect 9456 22380 9462 22432
rect 9490 22380 9496 22432
rect 9548 22420 9554 22432
rect 9861 22423 9919 22429
rect 9861 22420 9873 22423
rect 9548 22392 9873 22420
rect 9548 22380 9554 22392
rect 9861 22389 9873 22392
rect 9907 22389 9919 22423
rect 9861 22383 9919 22389
rect 12897 22423 12955 22429
rect 12897 22389 12909 22423
rect 12943 22420 12955 22423
rect 13170 22420 13176 22432
rect 12943 22392 13176 22420
rect 12943 22389 12955 22392
rect 12897 22383 12955 22389
rect 13170 22380 13176 22392
rect 13228 22420 13234 22432
rect 13446 22420 13452 22432
rect 13228 22392 13452 22420
rect 13228 22380 13234 22392
rect 13446 22380 13452 22392
rect 13504 22380 13510 22432
rect 13832 22420 13860 22528
rect 13909 22525 13921 22559
rect 13955 22556 13967 22559
rect 13998 22556 14004 22568
rect 13955 22528 14004 22556
rect 13955 22525 13967 22528
rect 13909 22519 13967 22525
rect 13998 22516 14004 22528
rect 14056 22516 14062 22568
rect 14554 22559 14612 22565
rect 14554 22525 14566 22559
rect 14600 22525 14612 22559
rect 14554 22519 14612 22525
rect 14737 22559 14795 22565
rect 14737 22525 14749 22559
rect 14783 22556 14795 22559
rect 17862 22556 17868 22568
rect 14783 22528 14872 22556
rect 17823 22528 17868 22556
rect 14783 22525 14795 22528
rect 14737 22519 14795 22525
rect 14568 22488 14596 22519
rect 14844 22500 14872 22528
rect 17862 22516 17868 22528
rect 17920 22556 17926 22568
rect 18138 22556 18144 22568
rect 17920 22528 18144 22556
rect 17920 22516 17926 22528
rect 18138 22516 18144 22528
rect 18196 22516 18202 22568
rect 18322 22556 18328 22568
rect 18283 22528 18328 22556
rect 18322 22516 18328 22528
rect 18380 22516 18386 22568
rect 20364 22565 20392 22596
rect 22186 22584 22192 22596
rect 22244 22584 22250 22636
rect 22296 22633 22324 22664
rect 22281 22627 22339 22633
rect 22281 22593 22293 22627
rect 22327 22624 22339 22627
rect 22922 22624 22928 22636
rect 22327 22596 22928 22624
rect 22327 22593 22339 22596
rect 22281 22587 22339 22593
rect 22922 22584 22928 22596
rect 22980 22584 22986 22636
rect 23385 22627 23443 22633
rect 23385 22593 23397 22627
rect 23431 22624 23443 22627
rect 23492 22624 23520 22732
rect 25869 22729 25881 22732
rect 25915 22729 25927 22763
rect 25869 22723 25927 22729
rect 27430 22720 27436 22772
rect 27488 22760 27494 22772
rect 28077 22763 28135 22769
rect 27488 22732 28028 22760
rect 27488 22720 27494 22732
rect 23566 22652 23572 22704
rect 23624 22692 23630 22704
rect 24756 22695 24814 22701
rect 23624 22664 23669 22692
rect 23624 22652 23630 22664
rect 24756 22661 24768 22695
rect 24802 22692 24814 22695
rect 25406 22692 25412 22704
rect 24802 22664 25412 22692
rect 24802 22661 24814 22664
rect 24756 22655 24814 22661
rect 25406 22652 25412 22664
rect 25464 22652 25470 22704
rect 26418 22652 26424 22704
rect 26476 22692 26482 22704
rect 26476 22664 27752 22692
rect 26476 22652 26482 22664
rect 23431 22596 23520 22624
rect 23661 22627 23719 22633
rect 23431 22593 23443 22596
rect 23385 22587 23443 22593
rect 23661 22593 23673 22627
rect 23707 22593 23719 22627
rect 23661 22587 23719 22593
rect 20073 22559 20131 22565
rect 20073 22525 20085 22559
rect 20119 22525 20131 22559
rect 20073 22519 20131 22525
rect 20349 22559 20407 22565
rect 20349 22525 20361 22559
rect 20395 22556 20407 22559
rect 21450 22556 21456 22568
rect 20395 22528 21456 22556
rect 20395 22525 20407 22528
rect 20349 22519 20407 22525
rect 14467 22460 14596 22488
rect 13906 22420 13912 22432
rect 13819 22392 13912 22420
rect 13906 22380 13912 22392
rect 13964 22420 13970 22432
rect 14467 22420 14495 22460
rect 14826 22448 14832 22500
rect 14884 22448 14890 22500
rect 15378 22448 15384 22500
rect 15436 22488 15442 22500
rect 18230 22488 18236 22500
rect 15436 22460 18236 22488
rect 15436 22448 15442 22460
rect 18230 22448 18236 22460
rect 18288 22448 18294 22500
rect 17310 22420 17316 22432
rect 13964 22392 17316 22420
rect 13964 22380 13970 22392
rect 17310 22380 17316 22392
rect 17368 22380 17374 22432
rect 17405 22423 17463 22429
rect 17405 22389 17417 22423
rect 17451 22420 17463 22423
rect 17494 22420 17500 22432
rect 17451 22392 17500 22420
rect 17451 22389 17463 22392
rect 17405 22383 17463 22389
rect 17494 22380 17500 22392
rect 17552 22380 17558 22432
rect 17773 22423 17831 22429
rect 17773 22389 17785 22423
rect 17819 22420 17831 22423
rect 18598 22420 18604 22432
rect 17819 22392 18604 22420
rect 17819 22389 17831 22392
rect 17773 22383 17831 22389
rect 18598 22380 18604 22392
rect 18656 22380 18662 22432
rect 18690 22380 18696 22432
rect 18748 22420 18754 22432
rect 18748 22392 18793 22420
rect 18748 22380 18754 22392
rect 19426 22380 19432 22432
rect 19484 22420 19490 22432
rect 19521 22423 19579 22429
rect 19521 22420 19533 22423
rect 19484 22392 19533 22420
rect 19484 22380 19490 22392
rect 19521 22389 19533 22392
rect 19567 22389 19579 22423
rect 20088 22420 20116 22519
rect 21450 22516 21456 22528
rect 21508 22516 21514 22568
rect 22465 22559 22523 22565
rect 22465 22525 22477 22559
rect 22511 22556 22523 22559
rect 23290 22556 23296 22568
rect 22511 22528 23296 22556
rect 22511 22525 22523 22528
rect 22465 22519 22523 22525
rect 23290 22516 23296 22528
rect 23348 22516 23354 22568
rect 20898 22448 20904 22500
rect 20956 22488 20962 22500
rect 23676 22488 23704 22587
rect 23750 22584 23756 22636
rect 23808 22624 23814 22636
rect 27522 22624 27528 22636
rect 23808 22596 23853 22624
rect 27483 22596 27528 22624
rect 23808 22584 23814 22596
rect 27522 22584 27528 22596
rect 27580 22584 27586 22636
rect 27724 22633 27752 22664
rect 27798 22652 27804 22704
rect 27856 22692 27862 22704
rect 27856 22664 27901 22692
rect 27856 22652 27862 22664
rect 27709 22627 27767 22633
rect 27709 22593 27721 22627
rect 27755 22593 27767 22627
rect 27709 22587 27767 22593
rect 27893 22627 27951 22633
rect 27893 22593 27905 22627
rect 27939 22593 27951 22627
rect 27893 22587 27951 22593
rect 24486 22556 24492 22568
rect 24447 22528 24492 22556
rect 24486 22516 24492 22528
rect 24544 22516 24550 22568
rect 20956 22460 23704 22488
rect 27908 22488 27936 22587
rect 28000 22556 28028 22732
rect 28077 22729 28089 22763
rect 28123 22760 28135 22763
rect 28442 22760 28448 22772
rect 28123 22732 28448 22760
rect 28123 22729 28135 22732
rect 28077 22723 28135 22729
rect 28442 22720 28448 22732
rect 28500 22720 28506 22772
rect 28804 22695 28862 22701
rect 28804 22661 28816 22695
rect 28850 22692 28862 22695
rect 29638 22692 29644 22704
rect 28850 22664 29644 22692
rect 28850 22661 28862 22664
rect 28804 22655 28862 22661
rect 29638 22652 29644 22664
rect 29696 22652 29702 22704
rect 28537 22559 28595 22565
rect 28537 22556 28549 22559
rect 28000 22528 28549 22556
rect 28537 22525 28549 22528
rect 28583 22525 28595 22559
rect 28537 22519 28595 22525
rect 28074 22488 28080 22500
rect 27908 22460 28080 22488
rect 20956 22448 20962 22460
rect 28074 22448 28080 22460
rect 28132 22448 28138 22500
rect 21082 22420 21088 22432
rect 20088 22392 21088 22420
rect 19521 22383 19579 22389
rect 21082 22380 21088 22392
rect 21140 22380 21146 22432
rect 23937 22423 23995 22429
rect 23937 22389 23949 22423
rect 23983 22420 23995 22423
rect 24118 22420 24124 22432
rect 23983 22392 24124 22420
rect 23983 22389 23995 22392
rect 23937 22383 23995 22389
rect 24118 22380 24124 22392
rect 24176 22380 24182 22432
rect 26694 22380 26700 22432
rect 26752 22420 26758 22432
rect 29917 22423 29975 22429
rect 29917 22420 29929 22423
rect 26752 22392 29929 22420
rect 26752 22380 26758 22392
rect 29917 22389 29929 22392
rect 29963 22389 29975 22423
rect 29917 22383 29975 22389
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 6914 22176 6920 22228
rect 6972 22216 6978 22228
rect 7653 22219 7711 22225
rect 7653 22216 7665 22219
rect 6972 22188 7665 22216
rect 6972 22176 6978 22188
rect 7653 22185 7665 22188
rect 7699 22185 7711 22219
rect 7653 22179 7711 22185
rect 9122 22176 9128 22228
rect 9180 22216 9186 22228
rect 12253 22219 12311 22225
rect 12253 22216 12265 22219
rect 9180 22188 12265 22216
rect 9180 22176 9186 22188
rect 12253 22185 12265 22188
rect 12299 22185 12311 22219
rect 12253 22179 12311 22185
rect 12802 22176 12808 22228
rect 12860 22216 12866 22228
rect 13538 22216 13544 22228
rect 12860 22188 13544 22216
rect 12860 22176 12866 22188
rect 13538 22176 13544 22188
rect 13596 22176 13602 22228
rect 14826 22216 14832 22228
rect 13832 22188 14832 22216
rect 8202 22148 8208 22160
rect 7300 22120 8208 22148
rect 7300 22080 7328 22120
rect 8202 22108 8208 22120
rect 8260 22108 8266 22160
rect 11054 22108 11060 22160
rect 11112 22148 11118 22160
rect 13357 22151 13415 22157
rect 11112 22120 11192 22148
rect 11112 22108 11118 22120
rect 7469 22083 7527 22089
rect 7469 22080 7481 22083
rect 7300 22052 7481 22080
rect 7469 22049 7481 22052
rect 7515 22049 7527 22083
rect 8294 22080 8300 22092
rect 8207 22052 8300 22080
rect 7469 22043 7527 22049
rect 8220 22021 8248 22052
rect 8294 22040 8300 22052
rect 8352 22080 8358 22092
rect 8352 22052 9076 22080
rect 8352 22040 8358 22052
rect 7377 22015 7435 22021
rect 7377 21981 7389 22015
rect 7423 21981 7435 22015
rect 7377 21975 7435 21981
rect 8205 22015 8263 22021
rect 8205 21981 8217 22015
rect 8251 21981 8263 22015
rect 8205 21975 8263 21981
rect 8389 22015 8447 22021
rect 8389 21981 8401 22015
rect 8435 21981 8447 22015
rect 8389 21975 8447 21981
rect 7392 21944 7420 21975
rect 7926 21944 7932 21956
rect 7392 21916 7932 21944
rect 7926 21904 7932 21916
rect 7984 21944 7990 21956
rect 8297 21947 8355 21953
rect 8297 21944 8309 21947
rect 7984 21916 8309 21944
rect 7984 21904 7990 21916
rect 8297 21913 8309 21916
rect 8343 21913 8355 21947
rect 8404 21944 8432 21975
rect 8570 21944 8576 21956
rect 8404 21916 8576 21944
rect 8297 21907 8355 21913
rect 8570 21904 8576 21916
rect 8628 21904 8634 21956
rect 8202 21836 8208 21888
rect 8260 21876 8266 21888
rect 8941 21879 8999 21885
rect 8941 21876 8953 21879
rect 8260 21848 8953 21876
rect 8260 21836 8266 21848
rect 8941 21845 8953 21848
rect 8987 21845 8999 21879
rect 9048 21876 9076 22052
rect 9306 22040 9312 22092
rect 9364 22080 9370 22092
rect 9401 22083 9459 22089
rect 9401 22080 9413 22083
rect 9364 22052 9413 22080
rect 9364 22040 9370 22052
rect 9401 22049 9413 22052
rect 9447 22049 9459 22083
rect 9401 22043 9459 22049
rect 9490 22040 9496 22092
rect 9548 22040 9554 22092
rect 9585 22083 9643 22089
rect 9585 22049 9597 22083
rect 9631 22080 9643 22083
rect 9674 22080 9680 22092
rect 9631 22052 9680 22080
rect 9631 22049 9643 22052
rect 9585 22043 9643 22049
rect 9674 22040 9680 22052
rect 9732 22040 9738 22092
rect 9122 21972 9128 22024
rect 9180 22012 9186 22024
rect 9508 22012 9536 22040
rect 9180 21984 9536 22012
rect 9180 21972 9186 21984
rect 10502 21972 10508 22024
rect 10560 22012 10566 22024
rect 10630 22015 10688 22021
rect 10630 22012 10642 22015
rect 10560 21984 10642 22012
rect 10560 21972 10566 21984
rect 10630 21981 10642 21984
rect 10676 21981 10688 22015
rect 11054 22012 11060 22024
rect 11015 21984 11060 22012
rect 10630 21975 10688 21981
rect 11054 21972 11060 21984
rect 11112 21972 11118 22024
rect 11164 22021 11192 22120
rect 13357 22117 13369 22151
rect 13403 22148 13415 22151
rect 13832 22148 13860 22188
rect 14826 22176 14832 22188
rect 14884 22216 14890 22228
rect 15289 22219 15347 22225
rect 15289 22216 15301 22219
rect 14884 22188 15301 22216
rect 14884 22176 14890 22188
rect 15289 22185 15301 22188
rect 15335 22216 15347 22219
rect 15378 22216 15384 22228
rect 15335 22188 15384 22216
rect 15335 22185 15347 22188
rect 15289 22179 15347 22185
rect 15378 22176 15384 22188
rect 15436 22176 15442 22228
rect 15473 22219 15531 22225
rect 15473 22185 15485 22219
rect 15519 22216 15531 22219
rect 15930 22216 15936 22228
rect 15519 22188 15936 22216
rect 15519 22185 15531 22188
rect 15473 22179 15531 22185
rect 15930 22176 15936 22188
rect 15988 22216 15994 22228
rect 18601 22219 18659 22225
rect 18601 22216 18613 22219
rect 15988 22188 16427 22216
rect 15988 22176 15994 22188
rect 13403 22120 13860 22148
rect 13403 22117 13415 22120
rect 13357 22111 13415 22117
rect 13906 22108 13912 22160
rect 13964 22148 13970 22160
rect 14182 22148 14188 22160
rect 13964 22120 14188 22148
rect 13964 22108 13970 22120
rect 14182 22108 14188 22120
rect 14240 22108 14246 22160
rect 11701 22083 11759 22089
rect 11701 22049 11713 22083
rect 11747 22080 11759 22083
rect 12894 22080 12900 22092
rect 11747 22052 12900 22080
rect 11747 22049 11759 22052
rect 11701 22043 11759 22049
rect 12894 22040 12900 22052
rect 12952 22040 12958 22092
rect 13538 22080 13544 22092
rect 13499 22052 13544 22080
rect 13538 22040 13544 22052
rect 13596 22040 13602 22092
rect 14016 22052 14964 22080
rect 11149 22015 11207 22021
rect 11149 21981 11161 22015
rect 11195 22012 11207 22015
rect 11422 22012 11428 22024
rect 11195 21984 11428 22012
rect 11195 21981 11207 21984
rect 11149 21975 11207 21981
rect 11422 21972 11428 21984
rect 11480 21972 11486 22024
rect 11514 21972 11520 22024
rect 11572 22012 11578 22024
rect 11609 22015 11667 22021
rect 11609 22012 11621 22015
rect 11572 21984 11621 22012
rect 11572 21972 11578 21984
rect 11609 21981 11621 21984
rect 11655 21981 11667 22015
rect 11609 21975 11667 21981
rect 11793 22015 11851 22021
rect 11793 21981 11805 22015
rect 11839 22012 11851 22015
rect 11882 22012 11888 22024
rect 11839 21984 11888 22012
rect 11839 21981 11851 21984
rect 11793 21975 11851 21981
rect 11882 21972 11888 21984
rect 11940 21972 11946 22024
rect 12342 21972 12348 22024
rect 12400 22012 12406 22024
rect 12437 22015 12495 22021
rect 12437 22012 12449 22015
rect 12400 21984 12449 22012
rect 12400 21972 12406 21984
rect 12437 21981 12449 21984
rect 12483 21981 12495 22015
rect 12437 21975 12495 21981
rect 12526 21972 12532 22024
rect 12584 22012 12590 22024
rect 12710 22012 12716 22024
rect 12584 21984 12629 22012
rect 12671 21984 12716 22012
rect 12584 21972 12590 21984
rect 12710 21972 12716 21984
rect 12768 21972 12774 22024
rect 12802 21972 12808 22024
rect 12860 22012 12866 22024
rect 13265 22015 13323 22021
rect 12860 21984 12905 22012
rect 12860 21972 12866 21984
rect 13265 21981 13277 22015
rect 13311 22012 13323 22015
rect 13354 22012 13360 22024
rect 13311 21984 13360 22012
rect 13311 21981 13323 21984
rect 13265 21975 13323 21981
rect 13354 21972 13360 21984
rect 13412 22012 13418 22024
rect 14016 22012 14044 22052
rect 14936 22024 14964 22052
rect 13412 21984 14044 22012
rect 14093 22015 14151 22021
rect 13412 21972 13418 21984
rect 14093 21981 14105 22015
rect 14139 21981 14151 22015
rect 14918 22012 14924 22024
rect 14879 21984 14924 22012
rect 14093 21975 14151 21981
rect 9309 21947 9367 21953
rect 9309 21913 9321 21947
rect 9355 21944 9367 21947
rect 9582 21944 9588 21956
rect 9355 21916 9588 21944
rect 9355 21913 9367 21916
rect 9309 21907 9367 21913
rect 9582 21904 9588 21916
rect 9640 21904 9646 21956
rect 10520 21916 12020 21944
rect 9490 21876 9496 21888
rect 9048 21848 9496 21876
rect 8941 21839 8999 21845
rect 9490 21836 9496 21848
rect 9548 21836 9554 21888
rect 10520 21885 10548 21916
rect 10505 21879 10563 21885
rect 10505 21845 10517 21879
rect 10551 21845 10563 21879
rect 10505 21839 10563 21845
rect 10689 21879 10747 21885
rect 10689 21845 10701 21879
rect 10735 21876 10747 21879
rect 10778 21876 10784 21888
rect 10735 21848 10784 21876
rect 10735 21845 10747 21848
rect 10689 21839 10747 21845
rect 10778 21836 10784 21848
rect 10836 21836 10842 21888
rect 11992 21876 12020 21916
rect 12066 21904 12072 21956
rect 12124 21944 12130 21956
rect 13541 21947 13599 21953
rect 13541 21944 13553 21947
rect 12124 21916 13553 21944
rect 12124 21904 12130 21916
rect 13541 21913 13553 21916
rect 13587 21913 13599 21947
rect 13541 21907 13599 21913
rect 12618 21876 12624 21888
rect 11992 21848 12624 21876
rect 12618 21836 12624 21848
rect 12676 21836 12682 21888
rect 13446 21836 13452 21888
rect 13504 21876 13510 21888
rect 14108 21876 14136 21975
rect 14918 21972 14924 21984
rect 14976 21972 14982 22024
rect 16399 22021 16427 22188
rect 18432 22188 18613 22216
rect 18230 22108 18236 22160
rect 18288 22148 18294 22160
rect 18432 22148 18460 22188
rect 18601 22185 18613 22188
rect 18647 22185 18659 22219
rect 18601 22179 18659 22185
rect 21450 22176 21456 22228
rect 21508 22216 21514 22228
rect 28258 22216 28264 22228
rect 21508 22188 28264 22216
rect 21508 22176 21514 22188
rect 28258 22176 28264 22188
rect 28316 22216 28322 22228
rect 28626 22216 28632 22228
rect 28316 22188 28632 22216
rect 28316 22176 28322 22188
rect 28626 22176 28632 22188
rect 28684 22216 28690 22228
rect 28684 22188 28764 22216
rect 28684 22176 28690 22188
rect 18288 22120 18460 22148
rect 20625 22151 20683 22157
rect 18288 22108 18294 22120
rect 20625 22117 20637 22151
rect 20671 22148 20683 22151
rect 20714 22148 20720 22160
rect 20671 22120 20720 22148
rect 20671 22117 20683 22120
rect 20625 22111 20683 22117
rect 20714 22108 20720 22120
rect 20772 22108 20778 22160
rect 22462 22148 22468 22160
rect 21376 22120 22468 22148
rect 18598 22040 18604 22092
rect 18656 22080 18662 22092
rect 21376 22080 21404 22120
rect 22462 22108 22468 22120
rect 22520 22108 22526 22160
rect 21542 22080 21548 22092
rect 18656 22052 21404 22080
rect 21503 22052 21548 22080
rect 18656 22040 18662 22052
rect 21542 22040 21548 22052
rect 21600 22040 21606 22092
rect 24397 22083 24455 22089
rect 24397 22080 24409 22083
rect 21652 22052 24409 22080
rect 16393 22015 16451 22021
rect 16393 21981 16405 22015
rect 16439 21981 16451 22015
rect 16393 21975 16451 21981
rect 16669 22015 16727 22021
rect 16669 21981 16681 22015
rect 16715 21981 16727 22015
rect 17218 22012 17224 22024
rect 17179 21984 17224 22012
rect 16669 21975 16727 21981
rect 16684 21944 16712 21975
rect 17218 21972 17224 21984
rect 17276 21972 17282 22024
rect 17494 22021 17500 22024
rect 17488 21975 17500 22021
rect 17552 22012 17558 22024
rect 17552 21984 17588 22012
rect 17494 21972 17500 21975
rect 17552 21972 17558 21984
rect 20162 21972 20168 22024
rect 20220 22012 20226 22024
rect 20346 22012 20352 22024
rect 20220 21984 20352 22012
rect 20220 21972 20226 21984
rect 20346 21972 20352 21984
rect 20404 21972 20410 22024
rect 20806 22012 20812 22024
rect 20767 21984 20812 22012
rect 20806 21972 20812 21984
rect 20864 21972 20870 22024
rect 21652 22012 21680 22052
rect 24397 22049 24409 22052
rect 24443 22080 24455 22083
rect 26237 22083 26295 22089
rect 26237 22080 26249 22083
rect 24443 22052 26249 22080
rect 24443 22049 24455 22052
rect 24397 22043 24455 22049
rect 26237 22049 26249 22052
rect 26283 22049 26295 22083
rect 26237 22043 26295 22049
rect 26513 22083 26571 22089
rect 26513 22049 26525 22083
rect 26559 22080 26571 22083
rect 28074 22080 28080 22092
rect 26559 22052 28080 22080
rect 26559 22049 26571 22052
rect 26513 22043 26571 22049
rect 20916 21984 21680 22012
rect 17310 21944 17316 21956
rect 16684 21916 17316 21944
rect 17310 21904 17316 21916
rect 17368 21944 17374 21956
rect 20916 21944 20944 21984
rect 21818 21972 21824 22024
rect 21876 22012 21882 22024
rect 22005 22015 22063 22021
rect 22005 22012 22017 22015
rect 21876 21984 22017 22012
rect 21876 21972 21882 21984
rect 22005 21981 22017 21984
rect 22051 21981 22063 22015
rect 22005 21975 22063 21981
rect 22094 21972 22100 22024
rect 22152 22012 22158 22024
rect 22152 21984 22197 22012
rect 22152 21972 22158 21984
rect 22462 21972 22468 22024
rect 22520 22021 22526 22024
rect 22520 22012 22528 22021
rect 22520 21984 22565 22012
rect 22520 21975 22528 21984
rect 22520 21972 22526 21975
rect 22922 21972 22928 22024
rect 22980 22012 22986 22024
rect 23109 22015 23167 22021
rect 23109 22012 23121 22015
rect 22980 21984 23121 22012
rect 22980 21972 22986 21984
rect 23109 21981 23121 21984
rect 23155 21981 23167 22015
rect 23385 22015 23443 22021
rect 23385 22012 23397 22015
rect 23109 21975 23167 21981
rect 23216 21984 23397 22012
rect 21358 21944 21364 21956
rect 17368 21916 20944 21944
rect 21319 21916 21364 21944
rect 17368 21904 17374 21916
rect 21358 21904 21364 21916
rect 21416 21904 21422 21956
rect 22278 21944 22284 21956
rect 22239 21916 22284 21944
rect 22278 21904 22284 21916
rect 22336 21904 22342 21956
rect 22373 21947 22431 21953
rect 22373 21913 22385 21947
rect 22419 21944 22431 21947
rect 22419 21916 22784 21944
rect 22419 21913 22431 21916
rect 22373 21907 22431 21913
rect 13504 21848 14136 21876
rect 13504 21836 13510 21848
rect 14182 21836 14188 21888
rect 14240 21876 14246 21888
rect 15289 21879 15347 21885
rect 14240 21848 14285 21876
rect 14240 21836 14246 21848
rect 15289 21845 15301 21879
rect 15335 21876 15347 21879
rect 15378 21876 15384 21888
rect 15335 21848 15384 21876
rect 15335 21845 15347 21848
rect 15289 21839 15347 21845
rect 15378 21836 15384 21848
rect 15436 21836 15442 21888
rect 16669 21879 16727 21885
rect 16669 21845 16681 21879
rect 16715 21876 16727 21879
rect 22094 21876 22100 21888
rect 16715 21848 22100 21876
rect 16715 21845 16727 21848
rect 16669 21839 16727 21845
rect 22094 21836 22100 21848
rect 22152 21836 22158 21888
rect 22646 21876 22652 21888
rect 22607 21848 22652 21876
rect 22646 21836 22652 21848
rect 22704 21836 22710 21888
rect 22756 21876 22784 21916
rect 22830 21904 22836 21956
rect 22888 21944 22894 21956
rect 23216 21944 23244 21984
rect 23385 21981 23397 21984
rect 23431 21981 23443 22015
rect 23385 21975 23443 21981
rect 23477 22015 23535 22021
rect 23477 21981 23489 22015
rect 23523 22012 23535 22015
rect 23750 22012 23756 22024
rect 23523 21984 23756 22012
rect 23523 21981 23535 21984
rect 23477 21975 23535 21981
rect 23750 21972 23756 21984
rect 23808 22012 23814 22024
rect 24670 22012 24676 22024
rect 23808 21984 24676 22012
rect 23808 21972 23814 21984
rect 24670 21972 24676 21984
rect 24728 21972 24734 22024
rect 26694 21972 26700 22024
rect 26752 22012 26758 22024
rect 27908 22021 27936 22052
rect 28074 22040 28080 22052
rect 28132 22040 28138 22092
rect 28537 22083 28595 22089
rect 28537 22049 28549 22083
rect 28583 22080 28595 22083
rect 28626 22080 28632 22092
rect 28583 22052 28632 22080
rect 28583 22049 28595 22052
rect 28537 22043 28595 22049
rect 28626 22040 28632 22052
rect 28684 22040 28690 22092
rect 28736 22080 28764 22188
rect 29549 22083 29607 22089
rect 29549 22080 29561 22083
rect 28736 22052 29561 22080
rect 29549 22049 29561 22052
rect 29595 22049 29607 22083
rect 29914 22080 29920 22092
rect 29875 22052 29920 22080
rect 29549 22043 29607 22049
rect 29914 22040 29920 22052
rect 29972 22040 29978 22092
rect 27525 22015 27583 22021
rect 27525 22012 27537 22015
rect 26752 21984 27537 22012
rect 26752 21972 26758 21984
rect 27525 21981 27537 21984
rect 27571 21981 27583 22015
rect 27525 21975 27583 21981
rect 27893 22015 27951 22021
rect 27893 21981 27905 22015
rect 27939 21981 27951 22015
rect 28718 22012 28724 22024
rect 28679 21984 28724 22012
rect 27893 21975 27951 21981
rect 28718 21972 28724 21984
rect 28776 21972 28782 22024
rect 29733 22015 29791 22021
rect 29733 21981 29745 22015
rect 29779 21981 29791 22015
rect 29733 21975 29791 21981
rect 22888 21916 23244 21944
rect 23293 21947 23351 21953
rect 22888 21904 22894 21916
rect 23293 21913 23305 21947
rect 23339 21944 23351 21947
rect 24394 21944 24400 21956
rect 23339 21916 24400 21944
rect 23339 21913 23351 21916
rect 23293 21907 23351 21913
rect 24394 21904 24400 21916
rect 24452 21904 24458 21956
rect 26234 21904 26240 21956
rect 26292 21944 26298 21956
rect 27709 21947 27767 21953
rect 27709 21944 27721 21947
rect 26292 21916 27721 21944
rect 26292 21904 26298 21916
rect 27709 21913 27721 21916
rect 27755 21913 27767 21947
rect 27709 21907 27767 21913
rect 27801 21947 27859 21953
rect 27801 21913 27813 21947
rect 27847 21944 27859 21947
rect 29748 21944 29776 21975
rect 27847 21916 28028 21944
rect 27847 21913 27859 21916
rect 27801 21907 27859 21913
rect 23014 21876 23020 21888
rect 22756 21848 23020 21876
rect 23014 21836 23020 21848
rect 23072 21836 23078 21888
rect 23658 21876 23664 21888
rect 23619 21848 23664 21876
rect 23658 21836 23664 21848
rect 23716 21836 23722 21888
rect 27724 21876 27752 21907
rect 28000 21888 28028 21916
rect 28092 21916 29776 21944
rect 27890 21876 27896 21888
rect 27724 21848 27896 21876
rect 27890 21836 27896 21848
rect 27948 21836 27954 21888
rect 27982 21836 27988 21888
rect 28040 21836 28046 21888
rect 28092 21885 28120 21916
rect 28077 21879 28135 21885
rect 28077 21845 28089 21879
rect 28123 21845 28135 21879
rect 28077 21839 28135 21845
rect 28350 21836 28356 21888
rect 28408 21876 28414 21888
rect 28905 21879 28963 21885
rect 28905 21876 28917 21879
rect 28408 21848 28917 21876
rect 28408 21836 28414 21848
rect 28905 21845 28917 21848
rect 28951 21845 28963 21879
rect 28905 21839 28963 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 9214 21632 9220 21684
rect 9272 21632 9278 21684
rect 9490 21632 9496 21684
rect 9548 21672 9554 21684
rect 10229 21675 10287 21681
rect 10229 21672 10241 21675
rect 9548 21644 10241 21672
rect 9548 21632 9554 21644
rect 10229 21641 10241 21644
rect 10275 21641 10287 21675
rect 11698 21672 11704 21684
rect 11659 21644 11704 21672
rect 10229 21635 10287 21641
rect 11698 21632 11704 21644
rect 11756 21632 11762 21684
rect 13906 21672 13912 21684
rect 12912 21644 13912 21672
rect 9232 21604 9260 21632
rect 8128 21576 9352 21604
rect 7742 21536 7748 21548
rect 7703 21508 7748 21536
rect 7742 21496 7748 21508
rect 7800 21496 7806 21548
rect 7926 21536 7932 21548
rect 7887 21508 7932 21536
rect 7926 21496 7932 21508
rect 7984 21496 7990 21548
rect 8128 21545 8156 21576
rect 8113 21539 8171 21545
rect 8113 21505 8125 21539
rect 8159 21505 8171 21539
rect 8113 21499 8171 21505
rect 8297 21539 8355 21545
rect 8297 21505 8309 21539
rect 8343 21536 8355 21539
rect 8478 21536 8484 21548
rect 8343 21508 8484 21536
rect 8343 21505 8355 21508
rect 8297 21499 8355 21505
rect 8478 21496 8484 21508
rect 8536 21496 8542 21548
rect 9324 21545 9352 21576
rect 12342 21564 12348 21616
rect 12400 21604 12406 21616
rect 12912 21604 12940 21644
rect 13906 21632 13912 21644
rect 13964 21632 13970 21684
rect 14826 21672 14832 21684
rect 14016 21644 14832 21672
rect 14016 21604 14044 21644
rect 14826 21632 14832 21644
rect 14884 21632 14890 21684
rect 14921 21675 14979 21681
rect 14921 21641 14933 21675
rect 14967 21672 14979 21675
rect 15194 21672 15200 21684
rect 14967 21644 15200 21672
rect 14967 21641 14979 21644
rect 14921 21635 14979 21641
rect 15194 21632 15200 21644
rect 15252 21632 15258 21684
rect 15378 21632 15384 21684
rect 15436 21672 15442 21684
rect 16482 21672 16488 21684
rect 15436 21644 16488 21672
rect 15436 21632 15442 21644
rect 16482 21632 16488 21644
rect 16540 21672 16546 21684
rect 17037 21675 17095 21681
rect 17037 21672 17049 21675
rect 16540 21644 17049 21672
rect 16540 21632 16546 21644
rect 17037 21641 17049 21644
rect 17083 21641 17095 21675
rect 17310 21672 17316 21684
rect 17271 21644 17316 21672
rect 17037 21635 17095 21641
rect 17310 21632 17316 21644
rect 17368 21632 17374 21684
rect 17586 21632 17592 21684
rect 17644 21672 17650 21684
rect 17865 21675 17923 21681
rect 17865 21672 17877 21675
rect 17644 21644 17877 21672
rect 17644 21632 17650 21644
rect 17865 21641 17877 21644
rect 17911 21641 17923 21675
rect 17865 21635 17923 21641
rect 20806 21632 20812 21684
rect 20864 21672 20870 21684
rect 23477 21675 23535 21681
rect 23477 21672 23489 21675
rect 20864 21644 23489 21672
rect 20864 21632 20870 21644
rect 23477 21641 23489 21644
rect 23523 21641 23535 21675
rect 23477 21635 23535 21641
rect 24305 21675 24363 21681
rect 24305 21641 24317 21675
rect 24351 21672 24363 21675
rect 25590 21672 25596 21684
rect 24351 21644 25596 21672
rect 24351 21641 24363 21644
rect 24305 21635 24363 21641
rect 25590 21632 25596 21644
rect 25648 21632 25654 21684
rect 26878 21632 26884 21684
rect 26936 21672 26942 21684
rect 26973 21675 27031 21681
rect 26973 21672 26985 21675
rect 26936 21644 26985 21672
rect 26936 21632 26942 21644
rect 26973 21641 26985 21644
rect 27019 21641 27031 21675
rect 26973 21635 27031 21641
rect 28169 21675 28227 21681
rect 28169 21641 28181 21675
rect 28215 21641 28227 21675
rect 28169 21635 28227 21641
rect 12400 21576 12940 21604
rect 13372 21576 14044 21604
rect 14185 21607 14243 21613
rect 12400 21564 12406 21576
rect 9217 21539 9275 21545
rect 9217 21505 9229 21539
rect 9263 21505 9275 21539
rect 9217 21499 9275 21505
rect 9309 21539 9367 21545
rect 9309 21505 9321 21539
rect 9355 21505 9367 21539
rect 9309 21499 9367 21505
rect 8018 21468 8024 21480
rect 7979 21440 8024 21468
rect 8018 21428 8024 21440
rect 8076 21428 8082 21480
rect 9232 21400 9260 21499
rect 9398 21496 9404 21548
rect 9456 21536 9462 21548
rect 9456 21508 9501 21536
rect 9456 21496 9462 21508
rect 9582 21496 9588 21548
rect 9640 21536 9646 21548
rect 10597 21539 10655 21545
rect 9640 21508 9685 21536
rect 9640 21496 9646 21508
rect 10597 21505 10609 21539
rect 10643 21536 10655 21539
rect 11054 21536 11060 21548
rect 10643 21508 11060 21536
rect 10643 21505 10655 21508
rect 10597 21499 10655 21505
rect 11054 21496 11060 21508
rect 11112 21536 11118 21548
rect 11698 21539 11756 21545
rect 11698 21536 11710 21539
rect 11112 21508 11710 21536
rect 11112 21496 11118 21508
rect 11698 21505 11710 21508
rect 11744 21536 11756 21539
rect 11882 21536 11888 21548
rect 11744 21508 11888 21536
rect 11744 21505 11756 21508
rect 11698 21499 11756 21505
rect 11882 21496 11888 21508
rect 11940 21496 11946 21548
rect 12066 21496 12072 21548
rect 12124 21496 12130 21548
rect 13262 21536 13268 21548
rect 13223 21508 13268 21536
rect 13262 21496 13268 21508
rect 13320 21496 13326 21548
rect 13372 21545 13400 21576
rect 14185 21573 14197 21607
rect 14231 21604 14243 21607
rect 14231 21576 15240 21604
rect 14231 21573 14243 21576
rect 14185 21567 14243 21573
rect 13357 21539 13415 21545
rect 13357 21505 13369 21539
rect 13403 21505 13415 21539
rect 13357 21499 13415 21505
rect 13449 21539 13507 21545
rect 13449 21505 13461 21539
rect 13495 21536 13507 21539
rect 13538 21536 13544 21548
rect 13495 21508 13544 21536
rect 13495 21505 13507 21508
rect 13449 21499 13507 21505
rect 13538 21496 13544 21508
rect 13596 21496 13602 21548
rect 13633 21539 13691 21545
rect 13633 21505 13645 21539
rect 13679 21536 13691 21539
rect 13814 21536 13820 21548
rect 13679 21508 13820 21536
rect 13679 21505 13691 21508
rect 13633 21499 13691 21505
rect 10686 21468 10692 21480
rect 10647 21440 10692 21468
rect 10686 21428 10692 21440
rect 10744 21428 10750 21480
rect 10873 21471 10931 21477
rect 10873 21437 10885 21471
rect 10919 21468 10931 21471
rect 11330 21468 11336 21480
rect 10919 21440 11336 21468
rect 10919 21437 10931 21440
rect 10873 21431 10931 21437
rect 11330 21428 11336 21440
rect 11388 21468 11394 21480
rect 12084 21468 12112 21496
rect 11388 21440 12112 21468
rect 11388 21428 11394 21440
rect 12158 21428 12164 21480
rect 12216 21468 12222 21480
rect 12216 21440 12261 21468
rect 12216 21428 12222 21440
rect 10410 21400 10416 21412
rect 9232 21372 10416 21400
rect 10410 21360 10416 21372
rect 10468 21360 10474 21412
rect 11517 21403 11575 21409
rect 11517 21369 11529 21403
rect 11563 21400 11575 21403
rect 11974 21400 11980 21412
rect 11563 21372 11980 21400
rect 11563 21369 11575 21372
rect 11517 21363 11575 21369
rect 11974 21360 11980 21372
rect 12032 21360 12038 21412
rect 12069 21403 12127 21409
rect 12069 21369 12081 21403
rect 12115 21400 12127 21403
rect 12342 21400 12348 21412
rect 12115 21372 12348 21400
rect 12115 21369 12127 21372
rect 12069 21363 12127 21369
rect 12342 21360 12348 21372
rect 12400 21400 12406 21412
rect 13648 21400 13676 21499
rect 13814 21496 13820 21508
rect 13872 21496 13878 21548
rect 14093 21539 14151 21545
rect 14093 21505 14105 21539
rect 14139 21505 14151 21539
rect 14093 21499 14151 21505
rect 14737 21539 14795 21545
rect 14737 21505 14749 21539
rect 14783 21536 14795 21539
rect 14826 21536 14832 21548
rect 14783 21508 14832 21536
rect 14783 21505 14795 21508
rect 14737 21499 14795 21505
rect 12400 21372 13676 21400
rect 14108 21400 14136 21499
rect 14826 21496 14832 21508
rect 14884 21496 14890 21548
rect 15212 21536 15240 21576
rect 15286 21564 15292 21616
rect 15344 21604 15350 21616
rect 15933 21607 15991 21613
rect 15933 21604 15945 21607
rect 15344 21576 15945 21604
rect 15344 21564 15350 21576
rect 15933 21573 15945 21576
rect 15979 21573 15991 21607
rect 15933 21567 15991 21573
rect 16022 21564 16028 21616
rect 16080 21604 16086 21616
rect 17154 21607 17212 21613
rect 17154 21604 17166 21607
rect 16080 21576 17166 21604
rect 16080 21564 16086 21576
rect 17154 21573 17166 21576
rect 17200 21604 17212 21607
rect 18690 21604 18696 21616
rect 17200 21576 18696 21604
rect 17200 21573 17212 21576
rect 17154 21567 17212 21573
rect 18690 21564 18696 21576
rect 18748 21564 18754 21616
rect 21085 21607 21143 21613
rect 21085 21573 21097 21607
rect 21131 21604 21143 21607
rect 21542 21604 21548 21616
rect 21131 21576 21548 21604
rect 21131 21573 21143 21576
rect 21085 21567 21143 21573
rect 21542 21564 21548 21576
rect 21600 21564 21606 21616
rect 21634 21564 21640 21616
rect 21692 21604 21698 21616
rect 22189 21607 22247 21613
rect 22189 21604 22201 21607
rect 21692 21576 22201 21604
rect 21692 21564 21698 21576
rect 22189 21573 22201 21576
rect 22235 21573 22247 21607
rect 22922 21604 22928 21616
rect 22189 21567 22247 21573
rect 22480 21576 22928 21604
rect 22480 21548 22508 21576
rect 22922 21564 22928 21576
rect 22980 21604 22986 21616
rect 23750 21604 23756 21616
rect 22980 21576 23756 21604
rect 22980 21564 22986 21576
rect 23750 21564 23756 21576
rect 23808 21604 23814 21616
rect 23808 21576 24624 21604
rect 23808 21564 23814 21576
rect 15838 21536 15844 21548
rect 15212 21508 15844 21536
rect 15838 21496 15844 21508
rect 15896 21496 15902 21548
rect 16669 21539 16727 21545
rect 16669 21505 16681 21539
rect 16715 21536 16727 21539
rect 16850 21536 16856 21548
rect 16715 21508 16856 21536
rect 16715 21505 16727 21508
rect 16669 21499 16727 21505
rect 16850 21496 16856 21508
rect 16908 21496 16914 21548
rect 17310 21496 17316 21548
rect 17368 21536 17374 21548
rect 19334 21545 19340 21548
rect 17773 21539 17831 21545
rect 17773 21536 17785 21539
rect 17368 21508 17785 21536
rect 17368 21496 17374 21508
rect 17773 21505 17785 21508
rect 17819 21505 17831 21539
rect 17773 21499 17831 21505
rect 19328 21499 19340 21545
rect 19392 21536 19398 21548
rect 21818 21536 21824 21548
rect 19392 21508 19428 21536
rect 21779 21508 21824 21536
rect 19334 21496 19340 21499
rect 19392 21496 19398 21508
rect 21818 21496 21824 21508
rect 21876 21496 21882 21548
rect 21969 21539 22027 21545
rect 21969 21505 21981 21539
rect 22015 21536 22027 21539
rect 22015 21505 22048 21536
rect 21969 21499 22048 21505
rect 15105 21471 15163 21477
rect 15105 21437 15117 21471
rect 15151 21468 15163 21471
rect 15378 21468 15384 21480
rect 15151 21440 15384 21468
rect 15151 21437 15163 21440
rect 15105 21431 15163 21437
rect 15378 21428 15384 21440
rect 15436 21428 15442 21480
rect 16945 21471 17003 21477
rect 16945 21468 16957 21471
rect 15580 21440 16957 21468
rect 15580 21412 15608 21440
rect 16945 21437 16957 21440
rect 16991 21437 17003 21471
rect 16945 21431 17003 21437
rect 19061 21471 19119 21477
rect 19061 21437 19073 21471
rect 19107 21437 19119 21471
rect 22020 21468 22048 21499
rect 22094 21496 22100 21548
rect 22152 21536 22158 21548
rect 22327 21539 22385 21545
rect 22152 21508 22197 21536
rect 22152 21496 22158 21508
rect 22327 21505 22339 21539
rect 22373 21536 22385 21539
rect 22462 21536 22468 21548
rect 22373 21508 22468 21536
rect 22373 21505 22385 21508
rect 22327 21499 22385 21505
rect 22462 21496 22468 21508
rect 22520 21496 22526 21548
rect 23293 21539 23351 21545
rect 23293 21505 23305 21539
rect 23339 21536 23351 21539
rect 23658 21536 23664 21548
rect 23339 21508 23664 21536
rect 23339 21505 23351 21508
rect 23293 21499 23351 21505
rect 23658 21496 23664 21508
rect 23716 21496 23722 21548
rect 23934 21536 23940 21548
rect 23895 21508 23940 21536
rect 23934 21496 23940 21508
rect 23992 21496 23998 21548
rect 24118 21536 24124 21548
rect 24079 21508 24124 21536
rect 24118 21496 24124 21508
rect 24176 21496 24182 21548
rect 24596 21536 24624 21576
rect 24670 21564 24676 21616
rect 24728 21604 24734 21616
rect 24857 21607 24915 21613
rect 24857 21604 24869 21607
rect 24728 21576 24869 21604
rect 24728 21564 24734 21576
rect 24857 21573 24869 21576
rect 24903 21573 24915 21607
rect 26234 21604 26240 21616
rect 26195 21576 26240 21604
rect 24857 21567 24915 21573
rect 26234 21564 26240 21576
rect 26292 21564 26298 21616
rect 28184 21604 28212 21635
rect 29058 21607 29116 21613
rect 29058 21604 29070 21607
rect 28184 21576 29070 21604
rect 29058 21573 29070 21576
rect 29104 21573 29116 21607
rect 29058 21567 29116 21573
rect 25041 21539 25099 21545
rect 25041 21536 25053 21539
rect 24596 21508 25053 21536
rect 25041 21505 25053 21508
rect 25087 21505 25099 21539
rect 25041 21499 25099 21505
rect 27154 21496 27160 21548
rect 27212 21536 27218 21548
rect 27341 21539 27399 21545
rect 27341 21536 27353 21539
rect 27212 21508 27353 21536
rect 27212 21496 27218 21508
rect 27341 21505 27353 21508
rect 27387 21505 27399 21539
rect 27341 21499 27399 21505
rect 27433 21539 27491 21545
rect 27433 21505 27445 21539
rect 27479 21536 27491 21539
rect 27706 21536 27712 21548
rect 27479 21508 27712 21536
rect 27479 21505 27491 21508
rect 27433 21499 27491 21505
rect 27706 21496 27712 21508
rect 27764 21536 27770 21548
rect 28350 21536 28356 21548
rect 27764 21508 28212 21536
rect 28311 21508 28356 21536
rect 27764 21496 27770 21508
rect 22554 21468 22560 21480
rect 22020 21440 22560 21468
rect 19061 21431 19119 21437
rect 15562 21400 15568 21412
rect 14108 21372 15568 21400
rect 12400 21360 12406 21372
rect 15562 21360 15568 21372
rect 15620 21360 15626 21412
rect 16117 21403 16175 21409
rect 16117 21369 16129 21403
rect 16163 21400 16175 21403
rect 16574 21400 16580 21412
rect 16163 21372 16580 21400
rect 16163 21369 16175 21372
rect 16117 21363 16175 21369
rect 16574 21360 16580 21372
rect 16632 21360 16638 21412
rect 8294 21292 8300 21344
rect 8352 21332 8358 21344
rect 8481 21335 8539 21341
rect 8481 21332 8493 21335
rect 8352 21304 8493 21332
rect 8352 21292 8358 21304
rect 8481 21301 8493 21304
rect 8527 21301 8539 21335
rect 8938 21332 8944 21344
rect 8899 21304 8944 21332
rect 8481 21295 8539 21301
rect 8938 21292 8944 21304
rect 8996 21292 9002 21344
rect 9030 21292 9036 21344
rect 9088 21332 9094 21344
rect 9582 21332 9588 21344
rect 9088 21304 9588 21332
rect 9088 21292 9094 21304
rect 9582 21292 9588 21304
rect 9640 21292 9646 21344
rect 10134 21292 10140 21344
rect 10192 21332 10198 21344
rect 10778 21332 10784 21344
rect 10192 21304 10784 21332
rect 10192 21292 10198 21304
rect 10778 21292 10784 21304
rect 10836 21332 10842 21344
rect 12158 21332 12164 21344
rect 10836 21304 12164 21332
rect 10836 21292 10842 21304
rect 12158 21292 12164 21304
rect 12216 21292 12222 21344
rect 12894 21292 12900 21344
rect 12952 21332 12958 21344
rect 12989 21335 13047 21341
rect 12989 21332 13001 21335
rect 12952 21304 13001 21332
rect 12952 21292 12958 21304
rect 12989 21301 13001 21304
rect 13035 21301 13047 21335
rect 12989 21295 13047 21301
rect 14918 21292 14924 21344
rect 14976 21332 14982 21344
rect 15105 21335 15163 21341
rect 15105 21332 15117 21335
rect 14976 21304 15117 21332
rect 14976 21292 14982 21304
rect 15105 21301 15117 21304
rect 15151 21301 15163 21335
rect 19076 21332 19104 21431
rect 22554 21428 22560 21440
rect 22612 21468 22618 21480
rect 22830 21468 22836 21480
rect 22612 21440 22836 21468
rect 22612 21428 22618 21440
rect 22830 21428 22836 21440
rect 22888 21428 22894 21480
rect 23109 21471 23167 21477
rect 23109 21437 23121 21471
rect 23155 21468 23167 21471
rect 23952 21468 23980 21496
rect 23155 21440 23980 21468
rect 27525 21471 27583 21477
rect 23155 21437 23167 21440
rect 23109 21431 23167 21437
rect 27525 21437 27537 21471
rect 27571 21437 27583 21471
rect 27525 21431 27583 21437
rect 21269 21403 21327 21409
rect 21269 21400 21281 21403
rect 19996 21372 21281 21400
rect 19996 21344 20024 21372
rect 21269 21369 21281 21372
rect 21315 21400 21327 21403
rect 23658 21400 23664 21412
rect 21315 21372 23664 21400
rect 21315 21369 21327 21372
rect 21269 21363 21327 21369
rect 23658 21360 23664 21372
rect 23716 21360 23722 21412
rect 27338 21360 27344 21412
rect 27396 21400 27402 21412
rect 27540 21400 27568 21431
rect 27396 21372 27568 21400
rect 27396 21360 27402 21372
rect 19978 21332 19984 21344
rect 19076 21304 19984 21332
rect 15105 21295 15163 21301
rect 19978 21292 19984 21304
rect 20036 21292 20042 21344
rect 20441 21335 20499 21341
rect 20441 21301 20453 21335
rect 20487 21332 20499 21335
rect 20530 21332 20536 21344
rect 20487 21304 20536 21332
rect 20487 21301 20499 21304
rect 20441 21295 20499 21301
rect 20530 21292 20536 21304
rect 20588 21332 20594 21344
rect 22002 21332 22008 21344
rect 20588 21304 22008 21332
rect 20588 21292 20594 21304
rect 22002 21292 22008 21304
rect 22060 21292 22066 21344
rect 22462 21332 22468 21344
rect 22423 21304 22468 21332
rect 22462 21292 22468 21304
rect 22520 21292 22526 21344
rect 24394 21292 24400 21344
rect 24452 21332 24458 21344
rect 26329 21335 26387 21341
rect 26329 21332 26341 21335
rect 24452 21304 26341 21332
rect 24452 21292 24458 21304
rect 26329 21301 26341 21304
rect 26375 21332 26387 21335
rect 26878 21332 26884 21344
rect 26375 21304 26884 21332
rect 26375 21301 26387 21304
rect 26329 21295 26387 21301
rect 26878 21292 26884 21304
rect 26936 21292 26942 21344
rect 28184 21332 28212 21508
rect 28350 21496 28356 21508
rect 28408 21496 28414 21548
rect 28810 21468 28816 21480
rect 28771 21440 28816 21468
rect 28810 21428 28816 21440
rect 28868 21428 28874 21480
rect 30193 21335 30251 21341
rect 30193 21332 30205 21335
rect 28184 21304 30205 21332
rect 30193 21301 30205 21304
rect 30239 21301 30251 21335
rect 30193 21295 30251 21301
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 8018 21088 8024 21140
rect 8076 21128 8082 21140
rect 8389 21131 8447 21137
rect 8389 21128 8401 21131
rect 8076 21100 8401 21128
rect 8076 21088 8082 21100
rect 8389 21097 8401 21100
rect 8435 21097 8447 21131
rect 8389 21091 8447 21097
rect 8478 21088 8484 21140
rect 8536 21128 8542 21140
rect 11054 21128 11060 21140
rect 8536 21100 11060 21128
rect 8536 21088 8542 21100
rect 7745 20995 7803 21001
rect 7745 20961 7757 20995
rect 7791 20992 7803 20995
rect 8662 20992 8668 21004
rect 7791 20964 8668 20992
rect 7791 20961 7803 20964
rect 7745 20955 7803 20961
rect 8662 20952 8668 20964
rect 8720 20952 8726 21004
rect 9122 20952 9128 21004
rect 9180 20992 9186 21004
rect 9508 21001 9536 21100
rect 11054 21088 11060 21100
rect 11112 21088 11118 21140
rect 19245 21131 19303 21137
rect 19245 21097 19257 21131
rect 19291 21128 19303 21131
rect 19334 21128 19340 21140
rect 19291 21100 19340 21128
rect 19291 21097 19303 21100
rect 19245 21091 19303 21097
rect 19334 21088 19340 21100
rect 19392 21088 19398 21140
rect 21545 21131 21603 21137
rect 21545 21097 21557 21131
rect 21591 21128 21603 21131
rect 22186 21128 22192 21140
rect 21591 21100 22192 21128
rect 21591 21097 21603 21100
rect 21545 21091 21603 21097
rect 22186 21088 22192 21100
rect 22244 21088 22250 21140
rect 25866 21088 25872 21140
rect 25924 21128 25930 21140
rect 27062 21128 27068 21140
rect 25924 21100 27068 21128
rect 25924 21088 25930 21100
rect 27062 21088 27068 21100
rect 27120 21088 27126 21140
rect 28261 21131 28319 21137
rect 28261 21097 28273 21131
rect 28307 21128 28319 21131
rect 28718 21128 28724 21140
rect 28307 21100 28724 21128
rect 28307 21097 28319 21100
rect 28261 21091 28319 21097
rect 28718 21088 28724 21100
rect 28776 21088 28782 21140
rect 9217 20995 9275 21001
rect 9217 20992 9229 20995
rect 9180 20964 9229 20992
rect 9180 20952 9186 20964
rect 9217 20961 9229 20964
rect 9263 20961 9275 20995
rect 9217 20955 9275 20961
rect 9493 20995 9551 21001
rect 9493 20961 9505 20995
rect 9539 20961 9551 20995
rect 9493 20955 9551 20961
rect 10410 20952 10416 21004
rect 10468 20992 10474 21004
rect 10781 20995 10839 21001
rect 10781 20992 10793 20995
rect 10468 20964 10793 20992
rect 10468 20952 10474 20964
rect 10781 20961 10793 20964
rect 10827 20992 10839 20995
rect 12342 20992 12348 21004
rect 10827 20964 12348 20992
rect 10827 20961 10839 20964
rect 10781 20955 10839 20961
rect 12342 20952 12348 20964
rect 12400 20952 12406 21004
rect 13722 20992 13728 21004
rect 12820 20964 13728 20992
rect 8113 20927 8171 20933
rect 8113 20893 8125 20927
rect 8159 20893 8171 20927
rect 8113 20887 8171 20893
rect 8205 20927 8263 20933
rect 8205 20893 8217 20927
rect 8251 20924 8263 20927
rect 8386 20924 8392 20936
rect 8251 20896 8392 20924
rect 8251 20893 8263 20896
rect 8205 20887 8263 20893
rect 8128 20856 8156 20887
rect 8386 20884 8392 20896
rect 8444 20884 8450 20936
rect 10502 20924 10508 20936
rect 10463 20896 10508 20924
rect 10502 20884 10508 20896
rect 10560 20884 10566 20936
rect 11146 20884 11152 20936
rect 11204 20924 11210 20936
rect 12820 20933 12848 20964
rect 13722 20952 13728 20964
rect 13780 20952 13786 21004
rect 19334 20952 19340 21004
rect 19392 20992 19398 21004
rect 19613 20995 19671 21001
rect 19613 20992 19625 20995
rect 19392 20964 19625 20992
rect 19392 20952 19398 20964
rect 19613 20961 19625 20964
rect 19659 20961 19671 20995
rect 22204 20992 22232 21088
rect 23658 21020 23664 21072
rect 23716 21060 23722 21072
rect 23716 21032 25728 21060
rect 23716 21020 23722 21032
rect 25700 21001 25728 21032
rect 25685 20995 25743 21001
rect 19613 20955 19671 20961
rect 22113 20964 22232 20992
rect 23492 20964 24716 20992
rect 12437 20927 12495 20933
rect 12437 20924 12449 20927
rect 11204 20896 12449 20924
rect 11204 20884 11210 20896
rect 12437 20893 12449 20896
rect 12483 20893 12495 20927
rect 12437 20887 12495 20893
rect 12805 20927 12863 20933
rect 12805 20893 12817 20927
rect 12851 20893 12863 20927
rect 12805 20887 12863 20893
rect 12894 20884 12900 20936
rect 12952 20924 12958 20936
rect 13354 20924 13360 20936
rect 12952 20896 12997 20924
rect 13315 20896 13360 20924
rect 12952 20884 12958 20896
rect 13354 20884 13360 20896
rect 13412 20884 13418 20936
rect 14553 20927 14611 20933
rect 14553 20893 14565 20927
rect 14599 20924 14611 20927
rect 16574 20924 16580 20936
rect 14599 20896 16580 20924
rect 14599 20893 14611 20896
rect 14553 20887 14611 20893
rect 16574 20884 16580 20896
rect 16632 20924 16638 20936
rect 16853 20927 16911 20933
rect 16853 20924 16865 20927
rect 16632 20896 16865 20924
rect 16632 20884 16638 20896
rect 16853 20893 16865 20896
rect 16899 20924 16911 20927
rect 19426 20924 19432 20936
rect 16899 20896 17264 20924
rect 19387 20896 19432 20924
rect 16899 20893 16911 20896
rect 16853 20887 16911 20893
rect 17236 20868 17264 20896
rect 19426 20884 19432 20896
rect 19484 20884 19490 20936
rect 19705 20927 19763 20933
rect 19705 20893 19717 20927
rect 19751 20893 19763 20927
rect 19705 20887 19763 20893
rect 8128 20828 8248 20856
rect 8220 20788 8248 20828
rect 11974 20816 11980 20868
rect 12032 20856 12038 20868
rect 12529 20859 12587 20865
rect 12529 20856 12541 20859
rect 12032 20828 12541 20856
rect 12032 20816 12038 20828
rect 12529 20825 12541 20828
rect 12575 20825 12587 20859
rect 12529 20819 12587 20825
rect 8570 20788 8576 20800
rect 8220 20760 8576 20788
rect 8570 20748 8576 20760
rect 8628 20788 8634 20800
rect 12253 20791 12311 20797
rect 12253 20788 12265 20791
rect 8628 20760 12265 20788
rect 8628 20748 8634 20760
rect 12253 20757 12265 20760
rect 12299 20757 12311 20791
rect 12544 20788 12572 20819
rect 12618 20816 12624 20868
rect 12676 20856 12682 20868
rect 14182 20856 14188 20868
rect 12676 20828 14188 20856
rect 12676 20816 12682 20828
rect 14182 20816 14188 20828
rect 14240 20816 14246 20868
rect 14826 20865 14832 20868
rect 14820 20819 14832 20865
rect 14884 20856 14890 20868
rect 17126 20865 17132 20868
rect 17120 20856 17132 20865
rect 14884 20828 14920 20856
rect 17087 20828 17132 20856
rect 14826 20816 14832 20819
rect 14884 20816 14890 20828
rect 17120 20819 17132 20828
rect 17126 20816 17132 20819
rect 17184 20816 17190 20868
rect 17218 20816 17224 20868
rect 17276 20816 17282 20868
rect 13449 20791 13507 20797
rect 13449 20788 13461 20791
rect 12544 20760 13461 20788
rect 12253 20751 12311 20757
rect 13449 20757 13461 20760
rect 13495 20757 13507 20791
rect 13449 20751 13507 20757
rect 15933 20791 15991 20797
rect 15933 20757 15945 20791
rect 15979 20788 15991 20791
rect 16298 20788 16304 20800
rect 15979 20760 16304 20788
rect 15979 20757 15991 20760
rect 15933 20751 15991 20757
rect 16298 20748 16304 20760
rect 16356 20748 16362 20800
rect 17402 20748 17408 20800
rect 17460 20788 17466 20800
rect 18233 20791 18291 20797
rect 18233 20788 18245 20791
rect 17460 20760 18245 20788
rect 17460 20748 17466 20760
rect 18233 20757 18245 20760
rect 18279 20757 18291 20791
rect 19720 20788 19748 20887
rect 19978 20884 19984 20936
rect 20036 20924 20042 20936
rect 20165 20927 20223 20933
rect 20165 20924 20177 20927
rect 20036 20896 20177 20924
rect 20036 20884 20042 20896
rect 20165 20893 20177 20896
rect 20211 20893 20223 20927
rect 20165 20887 20223 20893
rect 20806 20884 20812 20936
rect 20864 20924 20870 20936
rect 20864 20896 21772 20924
rect 20864 20884 20870 20896
rect 20432 20859 20490 20865
rect 20432 20825 20444 20859
rect 20478 20856 20490 20859
rect 21744 20856 21772 20896
rect 21818 20884 21824 20936
rect 21876 20924 21882 20936
rect 22002 20924 22008 20936
rect 21876 20896 22008 20924
rect 21876 20884 21882 20896
rect 22002 20884 22008 20896
rect 22060 20884 22066 20936
rect 22113 20933 22141 20964
rect 22098 20927 22156 20933
rect 22098 20893 22110 20927
rect 22144 20893 22156 20927
rect 22373 20927 22431 20933
rect 22373 20924 22385 20927
rect 22098 20887 22156 20893
rect 22204 20896 22385 20924
rect 22204 20856 22232 20896
rect 22373 20893 22385 20896
rect 22419 20893 22431 20927
rect 22373 20887 22431 20893
rect 22511 20927 22569 20933
rect 22511 20893 22523 20927
rect 22557 20924 22569 20927
rect 22922 20924 22928 20936
rect 22557 20896 22928 20924
rect 22557 20893 22569 20896
rect 22511 20887 22569 20893
rect 22922 20884 22928 20896
rect 22980 20884 22986 20936
rect 23198 20924 23204 20936
rect 23159 20896 23204 20924
rect 23198 20884 23204 20896
rect 23256 20884 23262 20936
rect 23382 20933 23388 20936
rect 23349 20927 23388 20933
rect 23349 20893 23361 20927
rect 23349 20887 23388 20893
rect 23382 20884 23388 20887
rect 23440 20884 23446 20936
rect 23492 20933 23520 20964
rect 23750 20933 23756 20936
rect 23477 20927 23535 20933
rect 23477 20893 23489 20927
rect 23523 20893 23535 20927
rect 23477 20887 23535 20893
rect 23707 20927 23756 20933
rect 23707 20893 23719 20927
rect 23753 20893 23756 20927
rect 23707 20887 23756 20893
rect 20478 20828 21680 20856
rect 21744 20828 22232 20856
rect 20478 20825 20490 20828
rect 20432 20819 20490 20825
rect 20530 20788 20536 20800
rect 19720 20760 20536 20788
rect 18233 20751 18291 20757
rect 20530 20748 20536 20760
rect 20588 20788 20594 20800
rect 20714 20788 20720 20800
rect 20588 20760 20720 20788
rect 20588 20748 20594 20760
rect 20714 20748 20720 20760
rect 20772 20748 20778 20800
rect 21652 20788 21680 20828
rect 22278 20816 22284 20868
rect 22336 20856 22342 20868
rect 23492 20856 23520 20887
rect 23750 20884 23756 20887
rect 23808 20884 23814 20936
rect 24394 20924 24400 20936
rect 24355 20896 24400 20924
rect 24394 20884 24400 20896
rect 24452 20884 24458 20936
rect 24688 20933 24716 20964
rect 25685 20961 25697 20995
rect 25731 20961 25743 20995
rect 25685 20955 25743 20961
rect 27982 20952 27988 21004
rect 28040 20992 28046 21004
rect 28350 20992 28356 21004
rect 28040 20964 28356 20992
rect 28040 20952 28046 20964
rect 28350 20952 28356 20964
rect 28408 20952 28414 21004
rect 24673 20927 24731 20933
rect 24673 20893 24685 20927
rect 24719 20924 24731 20927
rect 25130 20924 25136 20936
rect 24719 20896 25136 20924
rect 24719 20893 24731 20896
rect 24673 20887 24731 20893
rect 25130 20884 25136 20896
rect 25188 20884 25194 20936
rect 27706 20924 27712 20936
rect 27667 20896 27712 20924
rect 27706 20884 27712 20896
rect 27764 20884 27770 20936
rect 27890 20924 27896 20936
rect 27851 20896 27896 20924
rect 27890 20884 27896 20896
rect 27948 20884 27954 20936
rect 28074 20884 28080 20936
rect 28132 20924 28138 20936
rect 28813 20927 28871 20933
rect 28813 20924 28825 20927
rect 28132 20896 28825 20924
rect 28132 20884 28138 20896
rect 28813 20893 28825 20896
rect 28859 20893 28871 20927
rect 28813 20887 28871 20893
rect 22336 20828 23520 20856
rect 22336 20816 22342 20828
rect 23566 20816 23572 20868
rect 23624 20856 23630 20868
rect 25952 20859 26010 20865
rect 23624 20828 23669 20856
rect 23624 20816 23630 20828
rect 25952 20825 25964 20859
rect 25998 20856 26010 20859
rect 26234 20856 26240 20868
rect 25998 20828 26240 20856
rect 25998 20825 26010 20828
rect 25952 20819 26010 20825
rect 26234 20816 26240 20828
rect 26292 20816 26298 20868
rect 26786 20816 26792 20868
rect 26844 20856 26850 20868
rect 27522 20856 27528 20868
rect 26844 20828 27528 20856
rect 26844 20816 26850 20828
rect 27522 20816 27528 20828
rect 27580 20816 27586 20868
rect 27982 20816 27988 20868
rect 28040 20856 28046 20868
rect 28040 20828 28085 20856
rect 28040 20816 28046 20828
rect 22649 20791 22707 20797
rect 22649 20788 22661 20791
rect 21652 20760 22661 20788
rect 22649 20757 22661 20760
rect 22695 20757 22707 20791
rect 22649 20751 22707 20757
rect 23845 20791 23903 20797
rect 23845 20757 23857 20791
rect 23891 20788 23903 20791
rect 23934 20788 23940 20800
rect 23891 20760 23940 20788
rect 23891 20757 23903 20760
rect 23845 20751 23903 20757
rect 23934 20748 23940 20760
rect 23992 20748 23998 20800
rect 27430 20748 27436 20800
rect 27488 20788 27494 20800
rect 28905 20791 28963 20797
rect 28905 20788 28917 20791
rect 27488 20760 28917 20788
rect 27488 20748 27494 20760
rect 28905 20757 28917 20760
rect 28951 20757 28963 20791
rect 28905 20751 28963 20757
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 8021 20587 8079 20593
rect 8021 20553 8033 20587
rect 8067 20584 8079 20587
rect 9122 20584 9128 20596
rect 8067 20556 9128 20584
rect 8067 20553 8079 20556
rect 8021 20547 8079 20553
rect 9122 20544 9128 20556
rect 9180 20544 9186 20596
rect 9861 20587 9919 20593
rect 9861 20553 9873 20587
rect 9907 20584 9919 20587
rect 10502 20584 10508 20596
rect 9907 20556 10508 20584
rect 9907 20553 9919 20556
rect 9861 20547 9919 20553
rect 10502 20544 10508 20556
rect 10560 20544 10566 20596
rect 10594 20544 10600 20596
rect 10652 20584 10658 20596
rect 10689 20587 10747 20593
rect 10689 20584 10701 20587
rect 10652 20556 10701 20584
rect 10652 20544 10658 20556
rect 10689 20553 10701 20556
rect 10735 20553 10747 20587
rect 12250 20584 12256 20596
rect 10689 20547 10747 20553
rect 11624 20556 12256 20584
rect 8748 20519 8806 20525
rect 6656 20488 8524 20516
rect 6656 20457 6684 20488
rect 8496 20460 8524 20488
rect 8748 20485 8760 20519
rect 8794 20516 8806 20519
rect 8938 20516 8944 20528
rect 8794 20488 8944 20516
rect 8794 20485 8806 20488
rect 8748 20479 8806 20485
rect 8938 20476 8944 20488
rect 8996 20476 9002 20528
rect 9398 20476 9404 20528
rect 9456 20516 9462 20528
rect 11624 20516 11652 20556
rect 12250 20544 12256 20556
rect 12308 20544 12314 20596
rect 12342 20544 12348 20596
rect 12400 20584 12406 20596
rect 13078 20584 13084 20596
rect 12400 20556 12445 20584
rect 13039 20556 13084 20584
rect 12400 20544 12406 20556
rect 13078 20544 13084 20556
rect 13136 20544 13142 20596
rect 15562 20584 15568 20596
rect 15523 20556 15568 20584
rect 15562 20544 15568 20556
rect 15620 20544 15626 20596
rect 17126 20584 17132 20596
rect 17087 20556 17132 20584
rect 17126 20544 17132 20556
rect 17184 20544 17190 20596
rect 20806 20584 20812 20596
rect 18800 20556 20812 20584
rect 11790 20516 11796 20528
rect 9456 20488 11652 20516
rect 11751 20488 11796 20516
rect 9456 20476 9462 20488
rect 11790 20476 11796 20488
rect 11848 20476 11854 20528
rect 12710 20516 12716 20528
rect 12268 20488 12716 20516
rect 6641 20451 6699 20457
rect 6641 20417 6653 20451
rect 6687 20417 6699 20451
rect 6641 20411 6699 20417
rect 6908 20451 6966 20457
rect 6908 20417 6920 20451
rect 6954 20448 6966 20451
rect 8294 20448 8300 20460
rect 6954 20420 8300 20448
rect 6954 20417 6966 20420
rect 6908 20411 6966 20417
rect 8294 20408 8300 20420
rect 8352 20408 8358 20460
rect 8478 20448 8484 20460
rect 8391 20420 8484 20448
rect 8478 20408 8484 20420
rect 8536 20408 8542 20460
rect 10226 20408 10232 20460
rect 10284 20448 10290 20460
rect 10597 20451 10655 20457
rect 10597 20448 10609 20451
rect 10284 20420 10609 20448
rect 10284 20408 10290 20420
rect 10597 20417 10609 20420
rect 10643 20417 10655 20451
rect 10778 20448 10784 20460
rect 10739 20420 10784 20448
rect 10597 20411 10655 20417
rect 10778 20408 10784 20420
rect 10836 20408 10842 20460
rect 10870 20408 10876 20460
rect 10928 20448 10934 20460
rect 10928 20420 10973 20448
rect 10928 20408 10934 20420
rect 11882 20408 11888 20460
rect 11940 20448 11946 20460
rect 12268 20457 12296 20488
rect 12710 20476 12716 20488
rect 12768 20476 12774 20528
rect 15470 20516 15476 20528
rect 13004 20488 15476 20516
rect 13004 20460 13032 20488
rect 15470 20476 15476 20488
rect 15528 20476 15534 20528
rect 12161 20451 12219 20457
rect 12161 20448 12173 20451
rect 11940 20420 12173 20448
rect 11940 20408 11946 20420
rect 12161 20417 12173 20420
rect 12207 20417 12219 20451
rect 12161 20411 12219 20417
rect 12253 20451 12311 20457
rect 12253 20417 12265 20451
rect 12299 20417 12311 20451
rect 12986 20448 12992 20460
rect 12947 20420 12992 20448
rect 12253 20411 12311 20417
rect 12986 20408 12992 20420
rect 13044 20408 13050 20460
rect 14441 20451 14499 20457
rect 14441 20448 14453 20451
rect 13464 20420 14453 20448
rect 9490 20340 9496 20392
rect 9548 20380 9554 20392
rect 13464 20380 13492 20420
rect 14441 20417 14453 20420
rect 14487 20417 14499 20451
rect 14441 20411 14499 20417
rect 16758 20408 16764 20460
rect 16816 20448 16822 20460
rect 17034 20448 17040 20460
rect 16816 20420 17040 20448
rect 16816 20408 16822 20420
rect 17034 20408 17040 20420
rect 17092 20448 17098 20460
rect 17402 20448 17408 20460
rect 17092 20420 17408 20448
rect 17092 20408 17098 20420
rect 17402 20408 17408 20420
rect 17460 20408 17466 20460
rect 17497 20451 17555 20457
rect 17497 20417 17509 20451
rect 17543 20417 17555 20451
rect 17497 20411 17555 20417
rect 9548 20352 13492 20380
rect 9548 20340 9554 20352
rect 14090 20340 14096 20392
rect 14148 20380 14154 20392
rect 14185 20383 14243 20389
rect 14185 20380 14197 20383
rect 14148 20352 14197 20380
rect 14148 20340 14154 20352
rect 14185 20349 14197 20352
rect 14231 20349 14243 20383
rect 14185 20343 14243 20349
rect 17512 20324 17540 20411
rect 17586 20408 17592 20460
rect 17644 20448 17650 20460
rect 17773 20451 17831 20457
rect 17644 20420 17689 20448
rect 17644 20408 17650 20420
rect 17773 20417 17785 20451
rect 17819 20417 17831 20451
rect 17773 20411 17831 20417
rect 18509 20451 18567 20457
rect 18509 20417 18521 20451
rect 18555 20448 18567 20451
rect 18690 20448 18696 20460
rect 18555 20420 18696 20448
rect 18555 20417 18567 20420
rect 18509 20411 18567 20417
rect 17788 20380 17816 20411
rect 18690 20408 18696 20420
rect 18748 20408 18754 20460
rect 18800 20457 18828 20556
rect 20806 20544 20812 20556
rect 20864 20544 20870 20596
rect 22186 20544 22192 20596
rect 22244 20584 22250 20596
rect 23198 20584 23204 20596
rect 22244 20556 23204 20584
rect 22244 20544 22250 20556
rect 23198 20544 23204 20556
rect 23256 20544 23262 20596
rect 23474 20544 23480 20596
rect 23532 20584 23538 20596
rect 25041 20587 25099 20593
rect 25041 20584 25053 20587
rect 23532 20556 25053 20584
rect 23532 20544 23538 20556
rect 25041 20553 25053 20556
rect 25087 20553 25099 20587
rect 25041 20547 25099 20553
rect 25130 20544 25136 20596
rect 25188 20584 25194 20596
rect 25188 20556 25820 20584
rect 25188 20544 25194 20556
rect 19978 20516 19984 20528
rect 19260 20488 19984 20516
rect 19260 20457 19288 20488
rect 19978 20476 19984 20488
rect 20036 20476 20042 20528
rect 22088 20519 22146 20525
rect 22088 20485 22100 20519
rect 22134 20516 22146 20519
rect 22462 20516 22468 20528
rect 22134 20488 22468 20516
rect 22134 20485 22146 20488
rect 22088 20479 22146 20485
rect 22462 20476 22468 20488
rect 22520 20476 22526 20528
rect 23216 20516 23244 20544
rect 25792 20525 25820 20556
rect 26878 20544 26884 20596
rect 26936 20584 26942 20596
rect 27338 20584 27344 20596
rect 26936 20556 27344 20584
rect 26936 20544 26942 20556
rect 25777 20519 25835 20525
rect 23216 20488 25544 20516
rect 18785 20451 18843 20457
rect 18785 20417 18797 20451
rect 18831 20417 18843 20451
rect 18785 20411 18843 20417
rect 19245 20451 19303 20457
rect 19245 20417 19257 20451
rect 19291 20417 19303 20451
rect 19501 20451 19559 20457
rect 19501 20448 19513 20451
rect 19245 20411 19303 20417
rect 19352 20420 19513 20448
rect 19150 20380 19156 20392
rect 17788 20352 19156 20380
rect 11054 20272 11060 20324
rect 11112 20312 11118 20324
rect 11112 20284 12112 20312
rect 11112 20272 11118 20284
rect 11974 20244 11980 20256
rect 11935 20216 11980 20244
rect 11974 20204 11980 20216
rect 12032 20204 12038 20256
rect 12084 20253 12112 20284
rect 17494 20272 17500 20324
rect 17552 20272 17558 20324
rect 12069 20247 12127 20253
rect 12069 20213 12081 20247
rect 12115 20244 12127 20247
rect 12342 20244 12348 20256
rect 12115 20216 12348 20244
rect 12115 20213 12127 20216
rect 12069 20207 12127 20213
rect 12342 20204 12348 20216
rect 12400 20244 12406 20256
rect 13446 20244 13452 20256
rect 12400 20216 13452 20244
rect 12400 20204 12406 20216
rect 13446 20204 13452 20216
rect 13504 20204 13510 20256
rect 15470 20204 15476 20256
rect 15528 20244 15534 20256
rect 17788 20244 17816 20352
rect 19150 20340 19156 20352
rect 19208 20340 19214 20392
rect 19352 20380 19380 20420
rect 19501 20417 19513 20420
rect 19547 20417 19559 20451
rect 19501 20411 19559 20417
rect 21174 20408 21180 20460
rect 21232 20448 21238 20460
rect 21542 20448 21548 20460
rect 21232 20420 21548 20448
rect 21232 20408 21238 20420
rect 21542 20408 21548 20420
rect 21600 20448 21606 20460
rect 21821 20451 21879 20457
rect 21821 20448 21833 20451
rect 21600 20420 21833 20448
rect 21600 20408 21606 20420
rect 21821 20417 21833 20420
rect 21867 20417 21879 20451
rect 23658 20448 23664 20460
rect 23619 20420 23664 20448
rect 21821 20411 21879 20417
rect 23658 20408 23664 20420
rect 23716 20408 23722 20460
rect 23934 20457 23940 20460
rect 23928 20448 23940 20457
rect 23895 20420 23940 20448
rect 23928 20411 23940 20420
rect 23934 20408 23940 20411
rect 23992 20408 23998 20460
rect 25516 20457 25544 20488
rect 25777 20485 25789 20519
rect 25823 20485 25835 20519
rect 25777 20479 25835 20485
rect 25682 20457 25688 20460
rect 25501 20451 25559 20457
rect 25501 20417 25513 20451
rect 25547 20417 25559 20451
rect 25501 20411 25559 20417
rect 25649 20451 25688 20457
rect 25649 20417 25661 20451
rect 25649 20411 25688 20417
rect 25682 20408 25688 20411
rect 25740 20408 25746 20460
rect 25866 20451 25924 20457
rect 25866 20448 25878 20451
rect 25848 20417 25878 20448
rect 25912 20417 25924 20451
rect 25848 20411 25924 20417
rect 25966 20451 26024 20457
rect 25966 20417 25978 20451
rect 26012 20417 26024 20451
rect 25966 20411 26024 20417
rect 19260 20352 19380 20380
rect 18325 20315 18383 20321
rect 18325 20281 18337 20315
rect 18371 20312 18383 20315
rect 19260 20312 19288 20352
rect 25848 20324 25876 20411
rect 25976 20324 26004 20411
rect 26878 20408 26884 20460
rect 26936 20448 26942 20460
rect 27264 20457 27292 20556
rect 27338 20544 27344 20556
rect 27396 20544 27402 20596
rect 27522 20476 27528 20528
rect 27580 20516 27586 20528
rect 28169 20519 28227 20525
rect 28169 20516 28181 20519
rect 27580 20488 28181 20516
rect 27580 20476 27586 20488
rect 28169 20485 28181 20488
rect 28215 20485 28227 20519
rect 28169 20479 28227 20485
rect 26973 20451 27031 20457
rect 26973 20448 26985 20451
rect 26936 20420 26985 20448
rect 26936 20408 26942 20420
rect 26973 20417 26985 20420
rect 27019 20417 27031 20451
rect 26973 20411 27031 20417
rect 27066 20451 27124 20457
rect 27066 20417 27078 20451
rect 27112 20417 27124 20451
rect 27066 20411 27124 20417
rect 27249 20451 27307 20457
rect 27249 20417 27261 20451
rect 27295 20417 27307 20451
rect 27249 20411 27307 20417
rect 27341 20451 27399 20457
rect 27341 20417 27353 20451
rect 27387 20417 27399 20451
rect 27341 20411 27399 20417
rect 18371 20284 19288 20312
rect 18371 20281 18383 20284
rect 18325 20275 18383 20281
rect 22830 20272 22836 20324
rect 22888 20312 22894 20324
rect 23201 20315 23259 20321
rect 23201 20312 23213 20315
rect 22888 20284 23213 20312
rect 22888 20272 22894 20284
rect 23201 20281 23213 20284
rect 23247 20281 23259 20315
rect 25848 20284 25872 20324
rect 23201 20275 23259 20281
rect 25866 20272 25872 20284
rect 25924 20272 25930 20324
rect 25958 20272 25964 20324
rect 26016 20272 26022 20324
rect 27080 20312 27108 20411
rect 27356 20380 27384 20411
rect 27430 20408 27436 20460
rect 27488 20457 27494 20460
rect 27488 20448 27496 20457
rect 27488 20420 27533 20448
rect 27488 20411 27496 20420
rect 27488 20408 27494 20411
rect 28350 20380 28356 20392
rect 27356 20352 28356 20380
rect 28350 20340 28356 20352
rect 28408 20340 28414 20392
rect 27246 20312 27252 20324
rect 27080 20284 27252 20312
rect 27246 20272 27252 20284
rect 27304 20272 27310 20324
rect 27522 20272 27528 20324
rect 27580 20312 27586 20324
rect 28810 20312 28816 20324
rect 27580 20284 28816 20312
rect 27580 20272 27586 20284
rect 15528 20216 17816 20244
rect 15528 20204 15534 20216
rect 18138 20204 18144 20256
rect 18196 20244 18202 20256
rect 18693 20247 18751 20253
rect 18693 20244 18705 20247
rect 18196 20216 18705 20244
rect 18196 20204 18202 20216
rect 18693 20213 18705 20216
rect 18739 20244 18751 20247
rect 19242 20244 19248 20256
rect 18739 20216 19248 20244
rect 18739 20213 18751 20216
rect 18693 20207 18751 20213
rect 19242 20204 19248 20216
rect 19300 20244 19306 20256
rect 20530 20244 20536 20256
rect 19300 20216 20536 20244
rect 19300 20204 19306 20216
rect 20530 20204 20536 20216
rect 20588 20204 20594 20256
rect 20625 20247 20683 20253
rect 20625 20213 20637 20247
rect 20671 20244 20683 20247
rect 20806 20244 20812 20256
rect 20671 20216 20812 20244
rect 20671 20213 20683 20216
rect 20625 20207 20683 20213
rect 20806 20204 20812 20216
rect 20864 20204 20870 20256
rect 26142 20244 26148 20256
rect 26103 20216 26148 20244
rect 26142 20204 26148 20216
rect 26200 20204 26206 20256
rect 27614 20244 27620 20256
rect 27575 20216 27620 20244
rect 27614 20204 27620 20216
rect 27672 20204 27678 20256
rect 28276 20253 28304 20284
rect 28810 20272 28816 20284
rect 28868 20272 28874 20324
rect 28261 20247 28319 20253
rect 28261 20213 28273 20247
rect 28307 20213 28319 20247
rect 28261 20207 28319 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 9309 20043 9367 20049
rect 9309 20009 9321 20043
rect 9355 20040 9367 20043
rect 9490 20040 9496 20052
rect 9355 20012 9496 20040
rect 9355 20009 9367 20012
rect 9309 20003 9367 20009
rect 9490 20000 9496 20012
rect 9548 20000 9554 20052
rect 10137 20043 10195 20049
rect 10137 20009 10149 20043
rect 10183 20040 10195 20043
rect 10686 20040 10692 20052
rect 10183 20012 10692 20040
rect 10183 20009 10195 20012
rect 10137 20003 10195 20009
rect 10686 20000 10692 20012
rect 10744 20000 10750 20052
rect 10778 20000 10784 20052
rect 10836 20040 10842 20052
rect 10836 20012 11652 20040
rect 10836 20000 10842 20012
rect 9950 19932 9956 19984
rect 10008 19972 10014 19984
rect 11057 19975 11115 19981
rect 11057 19972 11069 19975
rect 10008 19944 11069 19972
rect 10008 19932 10014 19944
rect 11057 19941 11069 19944
rect 11103 19941 11115 19975
rect 11624 19972 11652 20012
rect 11698 20000 11704 20052
rect 11756 20040 11762 20052
rect 12345 20043 12403 20049
rect 12345 20040 12357 20043
rect 11756 20012 12357 20040
rect 11756 20000 11762 20012
rect 12345 20009 12357 20012
rect 12391 20009 12403 20043
rect 12345 20003 12403 20009
rect 12989 20043 13047 20049
rect 12989 20009 13001 20043
rect 13035 20009 13047 20043
rect 13170 20040 13176 20052
rect 13131 20012 13176 20040
rect 12989 20003 13047 20009
rect 13004 19972 13032 20003
rect 13170 20000 13176 20012
rect 13228 20000 13234 20052
rect 14737 20043 14795 20049
rect 14737 20009 14749 20043
rect 14783 20040 14795 20043
rect 14826 20040 14832 20052
rect 14783 20012 14832 20040
rect 14783 20009 14795 20012
rect 14737 20003 14795 20009
rect 14826 20000 14832 20012
rect 14884 20000 14890 20052
rect 17402 20040 17408 20052
rect 14936 20012 17408 20040
rect 13354 19972 13360 19984
rect 11624 19944 13360 19972
rect 11057 19935 11115 19941
rect 9309 19839 9367 19845
rect 9309 19805 9321 19839
rect 9355 19805 9367 19839
rect 9490 19836 9496 19848
rect 9451 19808 9496 19836
rect 9309 19799 9367 19805
rect 9324 19768 9352 19799
rect 9490 19796 9496 19808
rect 9548 19796 9554 19848
rect 10134 19836 10140 19848
rect 10095 19808 10140 19836
rect 10134 19796 10140 19808
rect 10192 19796 10198 19848
rect 10594 19796 10600 19848
rect 10652 19836 10658 19848
rect 10781 19839 10839 19845
rect 10781 19836 10793 19839
rect 10652 19808 10793 19836
rect 10652 19796 10658 19808
rect 10781 19805 10793 19808
rect 10827 19805 10839 19839
rect 10781 19799 10839 19805
rect 10965 19839 11023 19845
rect 10965 19805 10977 19839
rect 11011 19836 11023 19839
rect 11054 19836 11060 19848
rect 11011 19808 11060 19836
rect 11011 19805 11023 19808
rect 10965 19799 11023 19805
rect 11054 19796 11060 19808
rect 11112 19796 11118 19848
rect 11241 19839 11299 19845
rect 11241 19805 11253 19839
rect 11287 19805 11299 19839
rect 11241 19799 11299 19805
rect 10686 19768 10692 19780
rect 9324 19740 10692 19768
rect 10686 19728 10692 19740
rect 10744 19728 10750 19780
rect 11256 19768 11284 19799
rect 11790 19796 11796 19848
rect 11848 19836 11854 19848
rect 12176 19845 12204 19944
rect 13354 19932 13360 19944
rect 13412 19972 13418 19984
rect 13722 19972 13728 19984
rect 13412 19944 13728 19972
rect 13412 19932 13418 19944
rect 13722 19932 13728 19944
rect 13780 19932 13786 19984
rect 12820 19876 14136 19904
rect 12820 19845 12848 19876
rect 11977 19839 12035 19845
rect 11977 19836 11989 19839
rect 11848 19808 11989 19836
rect 11848 19796 11854 19808
rect 11977 19805 11989 19808
rect 12023 19805 12035 19839
rect 11977 19799 12035 19805
rect 12069 19839 12127 19845
rect 12069 19805 12081 19839
rect 12115 19805 12127 19839
rect 12069 19799 12127 19805
rect 12161 19839 12219 19845
rect 12161 19805 12173 19839
rect 12207 19805 12219 19839
rect 12805 19839 12863 19845
rect 12805 19836 12817 19839
rect 12161 19799 12219 19805
rect 12268 19808 12817 19836
rect 12084 19768 12112 19799
rect 12268 19780 12296 19808
rect 12805 19805 12817 19808
rect 12851 19805 12863 19839
rect 12805 19799 12863 19805
rect 12989 19839 13047 19845
rect 12989 19805 13001 19839
rect 13035 19836 13047 19839
rect 13446 19836 13452 19848
rect 13035 19808 13452 19836
rect 13035 19805 13047 19808
rect 12989 19799 13047 19805
rect 13446 19796 13452 19808
rect 13504 19796 13510 19848
rect 14108 19845 14136 19876
rect 14093 19839 14151 19845
rect 14093 19805 14105 19839
rect 14139 19805 14151 19839
rect 14093 19799 14151 19805
rect 12250 19768 12256 19780
rect 11256 19740 12256 19768
rect 12250 19728 12256 19740
rect 12308 19728 12314 19780
rect 14936 19768 14964 20012
rect 17402 20000 17408 20012
rect 17460 20000 17466 20052
rect 17497 20043 17555 20049
rect 17497 20009 17509 20043
rect 17543 20040 17555 20043
rect 17586 20040 17592 20052
rect 17543 20012 17592 20040
rect 17543 20009 17555 20012
rect 17497 20003 17555 20009
rect 17586 20000 17592 20012
rect 17644 20000 17650 20052
rect 18690 20040 18696 20052
rect 18651 20012 18696 20040
rect 18690 20000 18696 20012
rect 18748 20000 18754 20052
rect 19426 20000 19432 20052
rect 19484 20040 19490 20052
rect 19981 20043 20039 20049
rect 19981 20040 19993 20043
rect 19484 20012 19993 20040
rect 19484 20000 19490 20012
rect 19981 20009 19993 20012
rect 20027 20009 20039 20043
rect 19981 20003 20039 20009
rect 20530 20000 20536 20052
rect 20588 20040 20594 20052
rect 20809 20043 20867 20049
rect 20809 20040 20821 20043
rect 20588 20012 20821 20040
rect 20588 20000 20594 20012
rect 20809 20009 20821 20012
rect 20855 20009 20867 20043
rect 20809 20003 20867 20009
rect 22738 20000 22744 20052
rect 22796 20040 22802 20052
rect 22925 20043 22983 20049
rect 22925 20040 22937 20043
rect 22796 20012 22937 20040
rect 22796 20000 22802 20012
rect 22925 20009 22937 20012
rect 22971 20009 22983 20043
rect 22925 20003 22983 20009
rect 25682 20000 25688 20052
rect 25740 20040 25746 20052
rect 26050 20040 26056 20052
rect 25740 20012 26056 20040
rect 25740 20000 25746 20012
rect 26050 20000 26056 20012
rect 26108 20040 26114 20052
rect 26145 20043 26203 20049
rect 26145 20040 26157 20043
rect 26108 20012 26157 20040
rect 26108 20000 26114 20012
rect 26145 20009 26157 20012
rect 26191 20009 26203 20043
rect 26786 20040 26792 20052
rect 26747 20012 26792 20040
rect 26145 20003 26203 20009
rect 26786 20000 26792 20012
rect 26844 20000 26850 20052
rect 27246 20000 27252 20052
rect 27304 20040 27310 20052
rect 28813 20043 28871 20049
rect 28813 20040 28825 20043
rect 27304 20012 28825 20040
rect 27304 20000 27310 20012
rect 28813 20009 28825 20012
rect 28859 20009 28871 20043
rect 28813 20003 28871 20009
rect 15010 19932 15016 19984
rect 15068 19972 15074 19984
rect 16298 19972 16304 19984
rect 15068 19944 16304 19972
rect 15068 19932 15074 19944
rect 16298 19932 16304 19944
rect 16356 19932 16362 19984
rect 18966 19972 18972 19984
rect 18248 19944 18972 19972
rect 15028 19845 15056 19932
rect 16209 19907 16267 19913
rect 16209 19904 16221 19907
rect 15212 19876 16221 19904
rect 15212 19845 15240 19876
rect 16209 19873 16221 19876
rect 16255 19873 16267 19907
rect 18248 19904 18276 19944
rect 18966 19932 18972 19944
rect 19024 19932 19030 19984
rect 19610 19972 19616 19984
rect 19306 19944 19616 19972
rect 16209 19867 16267 19873
rect 17236 19876 18276 19904
rect 15013 19839 15071 19845
rect 15013 19805 15025 19839
rect 15059 19805 15071 19839
rect 15013 19799 15071 19805
rect 15105 19839 15163 19845
rect 15105 19805 15117 19839
rect 15151 19805 15163 19839
rect 15105 19799 15163 19805
rect 15197 19839 15255 19845
rect 15197 19805 15209 19839
rect 15243 19805 15255 19839
rect 15197 19799 15255 19805
rect 15381 19839 15439 19845
rect 15381 19805 15393 19839
rect 15427 19836 15439 19839
rect 15470 19836 15476 19848
rect 15427 19808 15476 19836
rect 15427 19805 15439 19808
rect 15381 19799 15439 19805
rect 15120 19768 15148 19799
rect 12406 19740 14320 19768
rect 14936 19740 15148 19768
rect 9582 19660 9588 19712
rect 9640 19700 9646 19712
rect 12406 19700 12434 19740
rect 9640 19672 12434 19700
rect 9640 19660 9646 19672
rect 12710 19660 12716 19712
rect 12768 19700 12774 19712
rect 14185 19703 14243 19709
rect 14185 19700 14197 19703
rect 12768 19672 14197 19700
rect 12768 19660 12774 19672
rect 14185 19669 14197 19672
rect 14231 19669 14243 19703
rect 14292 19700 14320 19740
rect 15396 19700 15424 19799
rect 15470 19796 15476 19808
rect 15528 19796 15534 19848
rect 15841 19839 15899 19845
rect 15841 19805 15853 19839
rect 15887 19836 15899 19839
rect 16390 19836 16396 19848
rect 15887 19808 16396 19836
rect 15887 19805 15899 19808
rect 15841 19799 15899 19805
rect 16390 19796 16396 19808
rect 16448 19836 16454 19848
rect 17129 19839 17187 19845
rect 17129 19836 17141 19839
rect 16448 19808 17141 19836
rect 16448 19796 16454 19808
rect 17129 19805 17141 19808
rect 17175 19805 17187 19839
rect 17129 19799 17187 19805
rect 16025 19771 16083 19777
rect 16025 19737 16037 19771
rect 16071 19768 16083 19771
rect 17236 19768 17264 19876
rect 17957 19839 18015 19845
rect 17957 19805 17969 19839
rect 18003 19805 18015 19839
rect 18138 19836 18144 19848
rect 18099 19808 18144 19836
rect 17957 19799 18015 19805
rect 16071 19740 17264 19768
rect 17313 19771 17371 19777
rect 16071 19737 16083 19740
rect 16025 19731 16083 19737
rect 17313 19737 17325 19771
rect 17359 19768 17371 19771
rect 17586 19768 17592 19780
rect 17359 19740 17592 19768
rect 17359 19737 17371 19740
rect 17313 19731 17371 19737
rect 17586 19728 17592 19740
rect 17644 19728 17650 19780
rect 17862 19728 17868 19780
rect 17920 19768 17926 19780
rect 17972 19768 18000 19799
rect 18138 19796 18144 19808
rect 18196 19796 18202 19848
rect 18248 19845 18276 19876
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19904 18383 19907
rect 19306 19904 19334 19944
rect 19610 19932 19616 19944
rect 19668 19932 19674 19984
rect 20254 19972 20260 19984
rect 19812 19944 20260 19972
rect 18371 19876 19334 19904
rect 19521 19907 19579 19913
rect 18371 19873 18383 19876
rect 18325 19867 18383 19873
rect 19521 19873 19533 19907
rect 19567 19904 19579 19907
rect 19702 19904 19708 19916
rect 19567 19876 19708 19904
rect 19567 19873 19579 19876
rect 19521 19867 19579 19873
rect 19702 19864 19708 19876
rect 19760 19864 19766 19916
rect 18233 19839 18291 19845
rect 18233 19805 18245 19839
rect 18279 19805 18291 19839
rect 18506 19836 18512 19848
rect 18467 19808 18512 19836
rect 18233 19799 18291 19805
rect 18506 19796 18512 19808
rect 18564 19796 18570 19848
rect 19245 19839 19303 19845
rect 19245 19805 19257 19839
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 19260 19768 19288 19799
rect 19334 19796 19340 19848
rect 19392 19836 19398 19848
rect 19429 19839 19487 19845
rect 19429 19836 19441 19839
rect 19392 19808 19441 19836
rect 19392 19796 19398 19808
rect 19429 19805 19441 19808
rect 19475 19805 19487 19839
rect 19610 19836 19616 19848
rect 19523 19808 19616 19836
rect 19429 19799 19487 19805
rect 19610 19796 19616 19808
rect 19668 19836 19674 19848
rect 19812 19845 19840 19944
rect 20254 19932 20260 19944
rect 20312 19932 20318 19984
rect 21542 19904 21548 19916
rect 21503 19876 21548 19904
rect 21542 19864 21548 19876
rect 21600 19864 21606 19916
rect 24486 19864 24492 19916
rect 24544 19904 24550 19916
rect 24765 19907 24823 19913
rect 24765 19904 24777 19907
rect 24544 19876 24777 19904
rect 24544 19864 24550 19876
rect 24765 19873 24777 19876
rect 24811 19873 24823 19907
rect 24765 19867 24823 19873
rect 19797 19839 19855 19845
rect 19668 19808 19748 19836
rect 19668 19796 19674 19808
rect 17920 19740 19288 19768
rect 19720 19768 19748 19808
rect 19797 19805 19809 19839
rect 19843 19805 19855 19839
rect 20622 19836 20628 19848
rect 20583 19808 20628 19836
rect 19797 19799 19855 19805
rect 20622 19796 20628 19808
rect 20680 19796 20686 19848
rect 20898 19836 20904 19848
rect 20811 19808 20904 19836
rect 20898 19796 20904 19808
rect 20956 19836 20962 19848
rect 21174 19836 21180 19848
rect 20956 19808 21180 19836
rect 20956 19796 20962 19808
rect 21174 19796 21180 19808
rect 21232 19796 21238 19848
rect 21812 19839 21870 19845
rect 21812 19805 21824 19839
rect 21858 19836 21870 19839
rect 22646 19836 22652 19848
rect 21858 19808 22652 19836
rect 21858 19805 21870 19808
rect 21812 19799 21870 19805
rect 22646 19796 22652 19808
rect 22704 19796 22710 19848
rect 25032 19839 25090 19845
rect 25032 19805 25044 19839
rect 25078 19836 25090 19839
rect 26142 19836 26148 19848
rect 25078 19808 26148 19836
rect 25078 19805 25090 19808
rect 25032 19799 25090 19805
rect 26142 19796 26148 19808
rect 26200 19796 26206 19848
rect 26970 19796 26976 19848
rect 27028 19836 27034 19848
rect 27433 19839 27491 19845
rect 27433 19836 27445 19839
rect 27028 19808 27445 19836
rect 27028 19796 27034 19808
rect 27433 19805 27445 19808
rect 27479 19836 27491 19839
rect 27522 19836 27528 19848
rect 27479 19808 27528 19836
rect 27479 19805 27491 19808
rect 27433 19799 27491 19805
rect 27522 19796 27528 19808
rect 27580 19796 27586 19848
rect 27700 19839 27758 19845
rect 27700 19805 27712 19839
rect 27746 19805 27758 19839
rect 27700 19799 27758 19805
rect 26694 19768 26700 19780
rect 19720 19740 20300 19768
rect 26655 19740 26700 19768
rect 17920 19728 17926 19740
rect 20272 19712 20300 19740
rect 26694 19728 26700 19740
rect 26752 19728 26758 19780
rect 27614 19728 27620 19780
rect 27672 19768 27678 19780
rect 27724 19768 27752 19799
rect 27672 19740 27752 19768
rect 27672 19728 27678 19740
rect 14292 19672 15424 19700
rect 14185 19663 14243 19669
rect 15746 19660 15752 19712
rect 15804 19700 15810 19712
rect 19426 19700 19432 19712
rect 15804 19672 19432 19700
rect 15804 19660 15810 19672
rect 19426 19660 19432 19672
rect 19484 19660 19490 19712
rect 20254 19660 20260 19712
rect 20312 19660 20318 19712
rect 20438 19700 20444 19712
rect 20399 19672 20444 19700
rect 20438 19660 20444 19672
rect 20496 19660 20502 19712
rect 27246 19660 27252 19712
rect 27304 19700 27310 19712
rect 27706 19700 27712 19712
rect 27304 19672 27712 19700
rect 27304 19660 27310 19672
rect 27706 19660 27712 19672
rect 27764 19660 27770 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 9401 19499 9459 19505
rect 9401 19465 9413 19499
rect 9447 19496 9459 19499
rect 9766 19496 9772 19508
rect 9447 19468 9772 19496
rect 9447 19465 9459 19468
rect 9401 19459 9459 19465
rect 9766 19456 9772 19468
rect 9824 19456 9830 19508
rect 12069 19499 12127 19505
rect 12069 19465 12081 19499
rect 12115 19496 12127 19499
rect 12526 19496 12532 19508
rect 12115 19468 12532 19496
rect 12115 19465 12127 19468
rect 12069 19459 12127 19465
rect 12526 19456 12532 19468
rect 12584 19456 12590 19508
rect 14277 19499 14335 19505
rect 14277 19465 14289 19499
rect 14323 19496 14335 19499
rect 14366 19496 14372 19508
rect 14323 19468 14372 19496
rect 14323 19465 14335 19468
rect 14277 19459 14335 19465
rect 14366 19456 14372 19468
rect 14424 19456 14430 19508
rect 23014 19496 23020 19508
rect 16960 19468 23020 19496
rect 10502 19428 10508 19440
rect 10152 19400 10508 19428
rect 10152 19360 10180 19400
rect 9508 19332 10180 19360
rect 9217 19295 9275 19301
rect 9217 19261 9229 19295
rect 9263 19292 9275 19295
rect 9508 19292 9536 19332
rect 10226 19320 10232 19372
rect 10284 19360 10290 19372
rect 10428 19369 10456 19400
rect 10502 19388 10508 19400
rect 10560 19428 10566 19440
rect 10870 19428 10876 19440
rect 10560 19400 10876 19428
rect 10560 19388 10566 19400
rect 10870 19388 10876 19400
rect 10928 19428 10934 19440
rect 11790 19428 11796 19440
rect 10928 19400 11796 19428
rect 10928 19388 10934 19400
rect 11790 19388 11796 19400
rect 11848 19388 11854 19440
rect 12621 19431 12679 19437
rect 12621 19397 12633 19431
rect 12667 19428 12679 19431
rect 13078 19428 13084 19440
rect 12667 19400 13084 19428
rect 12667 19397 12679 19400
rect 12621 19391 12679 19397
rect 13078 19388 13084 19400
rect 13136 19388 13142 19440
rect 14918 19428 14924 19440
rect 14879 19400 14924 19428
rect 14918 19388 14924 19400
rect 14976 19388 14982 19440
rect 15470 19388 15476 19440
rect 15528 19428 15534 19440
rect 15654 19428 15660 19440
rect 15528 19400 15660 19428
rect 15528 19388 15534 19400
rect 15654 19388 15660 19400
rect 15712 19428 15718 19440
rect 16960 19437 16988 19468
rect 16945 19431 17003 19437
rect 15712 19400 16160 19428
rect 15712 19388 15718 19400
rect 10321 19363 10379 19369
rect 10321 19360 10333 19363
rect 10284 19332 10333 19360
rect 10284 19320 10290 19332
rect 10321 19329 10333 19332
rect 10367 19329 10379 19363
rect 10321 19323 10379 19329
rect 10413 19363 10471 19369
rect 10413 19329 10425 19363
rect 10459 19329 10471 19363
rect 10594 19360 10600 19372
rect 10555 19332 10600 19360
rect 10413 19323 10471 19329
rect 10594 19320 10600 19332
rect 10652 19320 10658 19372
rect 10686 19320 10692 19372
rect 10744 19360 10750 19372
rect 11514 19360 11520 19372
rect 10744 19332 11100 19360
rect 11475 19332 11520 19360
rect 10744 19320 10750 19332
rect 9263 19264 9536 19292
rect 9585 19295 9643 19301
rect 9263 19261 9275 19264
rect 9217 19255 9275 19261
rect 9585 19261 9597 19295
rect 9631 19292 9643 19295
rect 10612 19292 10640 19320
rect 10962 19292 10968 19304
rect 9631 19264 10640 19292
rect 10923 19264 10968 19292
rect 9631 19261 9643 19264
rect 9585 19255 9643 19261
rect 10962 19252 10968 19264
rect 11020 19252 11026 19304
rect 11072 19292 11100 19332
rect 11514 19320 11520 19332
rect 11572 19320 11578 19372
rect 11808 19360 11836 19388
rect 11885 19363 11943 19369
rect 11885 19360 11897 19363
rect 11808 19332 11897 19360
rect 11885 19329 11897 19332
rect 11931 19329 11943 19363
rect 11885 19323 11943 19329
rect 13449 19363 13507 19369
rect 13449 19329 13461 19363
rect 13495 19360 13507 19363
rect 14093 19363 14151 19369
rect 14093 19360 14105 19363
rect 13495 19332 14105 19360
rect 13495 19329 13507 19332
rect 13449 19323 13507 19329
rect 14093 19329 14105 19332
rect 14139 19360 14151 19363
rect 14936 19360 14964 19388
rect 15746 19360 15752 19372
rect 14139 19332 14964 19360
rect 15707 19332 15752 19360
rect 14139 19329 14151 19332
rect 14093 19323 14151 19329
rect 15746 19320 15752 19332
rect 15804 19320 15810 19372
rect 15838 19320 15844 19372
rect 15896 19360 15902 19372
rect 16132 19369 16160 19400
rect 16945 19397 16957 19431
rect 16991 19397 17003 19431
rect 16945 19391 17003 19397
rect 17310 19388 17316 19440
rect 17368 19428 17374 19440
rect 17586 19428 17592 19440
rect 17368 19400 17592 19428
rect 17368 19388 17374 19400
rect 17586 19388 17592 19400
rect 17644 19388 17650 19440
rect 18138 19388 18144 19440
rect 18196 19428 18202 19440
rect 18196 19400 19380 19428
rect 18196 19388 18202 19400
rect 19352 19372 19380 19400
rect 20732 19400 22140 19428
rect 16117 19363 16175 19369
rect 15896 19332 15941 19360
rect 15896 19320 15902 19332
rect 16117 19329 16129 19363
rect 16163 19329 16175 19363
rect 16117 19323 16175 19329
rect 16390 19320 16396 19372
rect 16448 19360 16454 19372
rect 16761 19363 16819 19369
rect 16761 19360 16773 19363
rect 16448 19332 16773 19360
rect 16448 19320 16454 19332
rect 16761 19329 16773 19332
rect 16807 19329 16819 19363
rect 17862 19360 17868 19372
rect 17823 19332 17868 19360
rect 16761 19323 16819 19329
rect 17862 19320 17868 19332
rect 17920 19320 17926 19372
rect 19334 19320 19340 19372
rect 19392 19360 19398 19372
rect 20732 19369 20760 19400
rect 22112 19372 22140 19400
rect 19429 19363 19487 19369
rect 19429 19360 19441 19363
rect 19392 19332 19441 19360
rect 19392 19320 19398 19332
rect 19429 19329 19441 19332
rect 19475 19329 19487 19363
rect 19429 19323 19487 19329
rect 20533 19363 20591 19369
rect 20533 19329 20545 19363
rect 20579 19360 20591 19363
rect 20717 19363 20775 19369
rect 20579 19332 20668 19360
rect 20579 19329 20591 19332
rect 20533 19323 20591 19329
rect 15565 19295 15623 19301
rect 15565 19292 15577 19295
rect 11072 19264 15577 19292
rect 15565 19261 15577 19264
rect 15611 19261 15623 19295
rect 15565 19255 15623 19261
rect 16022 19252 16028 19304
rect 16080 19292 16086 19304
rect 17589 19295 17647 19301
rect 17589 19292 17601 19295
rect 16080 19264 17601 19292
rect 16080 19252 16086 19264
rect 17589 19261 17601 19264
rect 17635 19292 17647 19295
rect 18690 19292 18696 19304
rect 17635 19264 18696 19292
rect 17635 19261 17647 19264
rect 17589 19255 17647 19261
rect 18690 19252 18696 19264
rect 18748 19252 18754 19304
rect 19150 19292 19156 19304
rect 18800 19264 19156 19292
rect 8478 19184 8484 19236
rect 8536 19224 8542 19236
rect 12805 19227 12863 19233
rect 12805 19224 12817 19227
rect 8536 19196 12817 19224
rect 8536 19184 8542 19196
rect 12805 19193 12817 19196
rect 12851 19224 12863 19227
rect 14090 19224 14096 19236
rect 12851 19196 14096 19224
rect 12851 19193 12863 19196
rect 12805 19187 12863 19193
rect 14090 19184 14096 19196
rect 14148 19184 14154 19236
rect 18800 19224 18828 19264
rect 19150 19252 19156 19264
rect 19208 19252 19214 19304
rect 16040 19196 18828 19224
rect 20640 19224 20668 19332
rect 20717 19329 20729 19363
rect 20763 19329 20775 19363
rect 20717 19323 20775 19329
rect 20809 19363 20867 19369
rect 20809 19329 20821 19363
rect 20855 19360 20867 19363
rect 20990 19360 20996 19372
rect 20855 19332 20996 19360
rect 20855 19329 20867 19332
rect 20809 19323 20867 19329
rect 20990 19320 20996 19332
rect 21048 19320 21054 19372
rect 21085 19363 21143 19369
rect 21085 19329 21097 19363
rect 21131 19360 21143 19363
rect 21726 19360 21732 19372
rect 21131 19332 21732 19360
rect 21131 19329 21143 19332
rect 21085 19323 21143 19329
rect 21726 19320 21732 19332
rect 21784 19320 21790 19372
rect 21910 19360 21916 19372
rect 21871 19332 21916 19360
rect 21910 19320 21916 19332
rect 21968 19320 21974 19372
rect 22094 19360 22100 19372
rect 22007 19332 22100 19360
rect 22094 19320 22100 19332
rect 22152 19320 22158 19372
rect 22204 19369 22232 19468
rect 23014 19456 23020 19468
rect 23072 19456 23078 19508
rect 26234 19456 26240 19508
rect 26292 19496 26298 19508
rect 26329 19499 26387 19505
rect 26329 19496 26341 19499
rect 26292 19468 26341 19496
rect 26292 19456 26298 19468
rect 26329 19465 26341 19468
rect 26375 19465 26387 19499
rect 26329 19459 26387 19465
rect 27154 19456 27160 19508
rect 27212 19496 27218 19508
rect 28997 19499 29055 19505
rect 28997 19496 29009 19499
rect 27212 19468 29009 19496
rect 27212 19456 27218 19468
rect 28997 19465 29009 19468
rect 29043 19465 29055 19499
rect 28997 19459 29055 19465
rect 25961 19431 26019 19437
rect 25961 19397 25973 19431
rect 26007 19397 26019 19431
rect 25961 19391 26019 19397
rect 22189 19363 22247 19369
rect 22189 19329 22201 19363
rect 22235 19329 22247 19363
rect 22189 19323 22247 19329
rect 22370 19320 22376 19372
rect 22428 19360 22434 19372
rect 22465 19363 22523 19369
rect 22465 19360 22477 19363
rect 22428 19332 22477 19360
rect 22428 19320 22434 19332
rect 22465 19329 22477 19332
rect 22511 19329 22523 19363
rect 22465 19323 22523 19329
rect 23198 19320 23204 19372
rect 23256 19360 23262 19372
rect 23937 19363 23995 19369
rect 23937 19360 23949 19363
rect 23256 19332 23949 19360
rect 23256 19320 23262 19332
rect 23937 19329 23949 19332
rect 23983 19329 23995 19363
rect 23937 19323 23995 19329
rect 25685 19363 25743 19369
rect 25685 19329 25697 19363
rect 25731 19329 25743 19363
rect 25685 19323 25743 19329
rect 20901 19295 20959 19301
rect 20901 19261 20913 19295
rect 20947 19292 20959 19295
rect 22281 19295 22339 19301
rect 22281 19292 22293 19295
rect 20947 19264 22293 19292
rect 20947 19261 20959 19264
rect 20901 19255 20959 19261
rect 22204 19236 22232 19264
rect 22281 19261 22293 19264
rect 22327 19261 22339 19295
rect 22281 19255 22339 19261
rect 23661 19295 23719 19301
rect 23661 19261 23673 19295
rect 23707 19292 23719 19295
rect 25700 19292 25728 19323
rect 25774 19320 25780 19372
rect 25832 19360 25838 19372
rect 25832 19332 25877 19360
rect 25967 19358 25995 19391
rect 25832 19320 25838 19332
rect 25967 19330 26004 19358
rect 23707 19264 25728 19292
rect 25976 19292 26004 19330
rect 26050 19320 26056 19372
rect 26108 19369 26114 19372
rect 26234 19369 26240 19372
rect 26108 19363 26131 19369
rect 26119 19329 26131 19363
rect 26108 19323 26131 19329
rect 26191 19363 26240 19369
rect 26191 19329 26203 19363
rect 26237 19329 26240 19363
rect 26191 19323 26240 19329
rect 26108 19320 26114 19323
rect 26234 19320 26240 19323
rect 26292 19320 26298 19372
rect 26970 19320 26976 19372
rect 27028 19360 27034 19372
rect 27617 19363 27675 19369
rect 27617 19360 27629 19363
rect 27028 19332 27629 19360
rect 27028 19320 27034 19332
rect 27617 19329 27629 19332
rect 27663 19329 27675 19363
rect 27617 19323 27675 19329
rect 27706 19320 27712 19372
rect 27764 19360 27770 19372
rect 27873 19363 27931 19369
rect 27873 19360 27885 19363
rect 27764 19332 27885 19360
rect 27764 19320 27770 19332
rect 27873 19329 27885 19332
rect 27919 19329 27931 19363
rect 27873 19323 27931 19329
rect 27338 19292 27344 19304
rect 25976 19264 27344 19292
rect 23707 19261 23719 19264
rect 23661 19255 23719 19261
rect 21910 19224 21916 19236
rect 20640 19196 21916 19224
rect 9766 19156 9772 19168
rect 9727 19128 9772 19156
rect 9766 19116 9772 19128
rect 9824 19116 9830 19168
rect 10594 19116 10600 19168
rect 10652 19156 10658 19168
rect 11609 19159 11667 19165
rect 11609 19156 11621 19159
rect 10652 19128 11621 19156
rect 10652 19116 10658 19128
rect 11609 19125 11621 19128
rect 11655 19125 11667 19159
rect 13538 19156 13544 19168
rect 13499 19128 13544 19156
rect 11609 19119 11667 19125
rect 13538 19116 13544 19128
rect 13596 19116 13602 19168
rect 14458 19116 14464 19168
rect 14516 19156 14522 19168
rect 15013 19159 15071 19165
rect 15013 19156 15025 19159
rect 14516 19128 15025 19156
rect 14516 19116 14522 19128
rect 15013 19125 15025 19128
rect 15059 19125 15071 19159
rect 15013 19119 15071 19125
rect 15102 19116 15108 19168
rect 15160 19156 15166 19168
rect 16040 19165 16068 19196
rect 21910 19184 21916 19196
rect 21968 19184 21974 19236
rect 22186 19184 22192 19236
rect 22244 19184 22250 19236
rect 22462 19184 22468 19236
rect 22520 19224 22526 19236
rect 23676 19224 23704 19255
rect 22520 19196 23704 19224
rect 22520 19184 22526 19196
rect 16025 19159 16083 19165
rect 16025 19156 16037 19159
rect 15160 19128 16037 19156
rect 15160 19116 15166 19128
rect 16025 19125 16037 19128
rect 16071 19125 16083 19159
rect 16025 19119 16083 19125
rect 17129 19159 17187 19165
rect 17129 19125 17141 19159
rect 17175 19156 17187 19159
rect 18138 19156 18144 19168
rect 17175 19128 18144 19156
rect 17175 19125 17187 19128
rect 17129 19119 17187 19125
rect 18138 19116 18144 19128
rect 18196 19116 18202 19168
rect 19058 19116 19064 19168
rect 19116 19156 19122 19168
rect 20162 19156 20168 19168
rect 19116 19128 20168 19156
rect 19116 19116 19122 19128
rect 20162 19116 20168 19128
rect 20220 19116 20226 19168
rect 21269 19159 21327 19165
rect 21269 19125 21281 19159
rect 21315 19156 21327 19159
rect 21726 19156 21732 19168
rect 21315 19128 21732 19156
rect 21315 19125 21327 19128
rect 21269 19119 21327 19125
rect 21726 19116 21732 19128
rect 21784 19116 21790 19168
rect 22370 19116 22376 19168
rect 22428 19156 22434 19168
rect 22649 19159 22707 19165
rect 22649 19156 22661 19159
rect 22428 19128 22661 19156
rect 22428 19116 22434 19128
rect 22649 19125 22661 19128
rect 22695 19125 22707 19159
rect 22649 19119 22707 19125
rect 23382 19116 23388 19168
rect 23440 19156 23446 19168
rect 24946 19156 24952 19168
rect 23440 19128 24952 19156
rect 23440 19116 23446 19128
rect 24946 19116 24952 19128
rect 25004 19116 25010 19168
rect 25700 19156 25728 19264
rect 27338 19252 27344 19264
rect 27396 19252 27402 19304
rect 26234 19156 26240 19168
rect 25700 19128 26240 19156
rect 26234 19116 26240 19128
rect 26292 19116 26298 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 9766 18912 9772 18964
rect 9824 18952 9830 18964
rect 10226 18952 10232 18964
rect 9824 18924 10232 18952
rect 9824 18912 9830 18924
rect 10226 18912 10232 18924
rect 10284 18952 10290 18964
rect 10778 18952 10784 18964
rect 10284 18924 10784 18952
rect 10284 18912 10290 18924
rect 10778 18912 10784 18924
rect 10836 18952 10842 18964
rect 11514 18952 11520 18964
rect 10836 18924 11520 18952
rect 10836 18912 10842 18924
rect 11514 18912 11520 18924
rect 11572 18952 11578 18964
rect 11793 18955 11851 18961
rect 11793 18952 11805 18955
rect 11572 18924 11805 18952
rect 11572 18912 11578 18924
rect 11793 18921 11805 18924
rect 11839 18921 11851 18955
rect 11793 18915 11851 18921
rect 12158 18912 12164 18964
rect 12216 18952 12222 18964
rect 12253 18955 12311 18961
rect 12253 18952 12265 18955
rect 12216 18924 12265 18952
rect 12216 18912 12222 18924
rect 12253 18921 12265 18924
rect 12299 18921 12311 18955
rect 12253 18915 12311 18921
rect 14366 18912 14372 18964
rect 14424 18952 14430 18964
rect 17678 18952 17684 18964
rect 14424 18924 17448 18952
rect 17639 18924 17684 18952
rect 14424 18912 14430 18924
rect 14918 18884 14924 18896
rect 14569 18856 14924 18884
rect 11977 18819 12035 18825
rect 11977 18816 11989 18819
rect 10428 18788 11989 18816
rect 10428 18760 10456 18788
rect 11977 18785 11989 18788
rect 12023 18785 12035 18819
rect 13814 18816 13820 18828
rect 11977 18779 12035 18785
rect 13188 18788 13820 18816
rect 10410 18748 10416 18760
rect 10371 18720 10416 18748
rect 10410 18708 10416 18720
rect 10468 18708 10474 18760
rect 10502 18708 10508 18760
rect 10560 18748 10566 18760
rect 10689 18751 10747 18757
rect 10689 18748 10701 18751
rect 10560 18720 10701 18748
rect 10560 18708 10566 18720
rect 10689 18717 10701 18720
rect 10735 18717 10747 18751
rect 11701 18751 11759 18757
rect 11701 18748 11713 18751
rect 10689 18711 10747 18717
rect 10796 18720 11713 18748
rect 10594 18640 10600 18692
rect 10652 18680 10658 18692
rect 10796 18680 10824 18720
rect 11701 18717 11713 18720
rect 11747 18717 11759 18751
rect 13078 18748 13084 18760
rect 13039 18720 13084 18748
rect 11701 18711 11759 18717
rect 13078 18708 13084 18720
rect 13136 18708 13142 18760
rect 13188 18757 13216 18788
rect 13814 18776 13820 18788
rect 13872 18776 13878 18828
rect 13173 18751 13231 18757
rect 13173 18717 13185 18751
rect 13219 18717 13231 18751
rect 13173 18711 13231 18717
rect 13265 18751 13323 18757
rect 13265 18717 13277 18751
rect 13311 18717 13323 18751
rect 13265 18711 13323 18717
rect 13449 18751 13507 18757
rect 13449 18717 13461 18751
rect 13495 18748 13507 18751
rect 14366 18748 14372 18760
rect 13495 18720 14372 18748
rect 13495 18717 13507 18720
rect 13449 18711 13507 18717
rect 10652 18652 10824 18680
rect 10652 18640 10658 18652
rect 10870 18640 10876 18692
rect 10928 18680 10934 18692
rect 13280 18680 13308 18711
rect 14366 18708 14372 18720
rect 14424 18708 14430 18760
rect 14569 18757 14597 18856
rect 14918 18844 14924 18856
rect 14976 18844 14982 18896
rect 15470 18816 15476 18828
rect 14660 18788 15476 18816
rect 14660 18757 14688 18788
rect 15470 18776 15476 18788
rect 15528 18776 15534 18828
rect 16117 18819 16175 18825
rect 16117 18785 16129 18819
rect 16163 18816 16175 18819
rect 16574 18816 16580 18828
rect 16163 18788 16580 18816
rect 16163 18785 16175 18788
rect 16117 18779 16175 18785
rect 16574 18776 16580 18788
rect 16632 18776 16638 18828
rect 17126 18816 17132 18828
rect 17052 18788 17132 18816
rect 14553 18751 14611 18757
rect 14553 18717 14565 18751
rect 14599 18717 14611 18751
rect 14553 18711 14611 18717
rect 14645 18751 14703 18757
rect 14645 18717 14657 18751
rect 14691 18717 14703 18751
rect 14645 18711 14703 18717
rect 14758 18748 14816 18754
rect 14758 18714 14770 18748
rect 14804 18714 14816 18748
rect 14758 18708 14816 18714
rect 14918 18708 14924 18760
rect 14976 18748 14982 18760
rect 14976 18720 15021 18748
rect 14976 18708 14982 18720
rect 15286 18708 15292 18760
rect 15344 18748 15350 18760
rect 15749 18751 15807 18757
rect 15749 18748 15761 18751
rect 15344 18720 15761 18748
rect 15344 18708 15350 18720
rect 15749 18717 15761 18720
rect 15795 18748 15807 18751
rect 15838 18748 15844 18760
rect 15795 18720 15844 18748
rect 15795 18717 15807 18720
rect 15749 18711 15807 18717
rect 15838 18708 15844 18720
rect 15896 18708 15902 18760
rect 16022 18748 16028 18760
rect 15983 18720 16028 18748
rect 16022 18708 16028 18720
rect 16080 18708 16086 18760
rect 16850 18748 16856 18760
rect 16811 18720 16856 18748
rect 16850 18708 16856 18720
rect 16908 18708 16914 18760
rect 17052 18757 17080 18788
rect 17126 18776 17132 18788
rect 17184 18776 17190 18828
rect 16942 18748 17000 18754
rect 16942 18714 16954 18748
rect 16988 18714 17000 18748
rect 16942 18708 17000 18714
rect 17037 18751 17095 18757
rect 17037 18717 17049 18751
rect 17083 18717 17095 18751
rect 17037 18711 17095 18717
rect 17233 18751 17291 18757
rect 17233 18717 17245 18751
rect 17279 18748 17291 18751
rect 17420 18748 17448 18924
rect 17678 18912 17684 18924
rect 17736 18912 17742 18964
rect 17862 18912 17868 18964
rect 17920 18952 17926 18964
rect 21085 18955 21143 18961
rect 17920 18924 20668 18952
rect 17920 18912 17926 18924
rect 20530 18884 20536 18896
rect 17926 18856 20536 18884
rect 17926 18757 17954 18856
rect 20530 18844 20536 18856
rect 20588 18844 20594 18896
rect 20640 18884 20668 18924
rect 21085 18921 21097 18955
rect 21131 18952 21143 18955
rect 21358 18952 21364 18964
rect 21131 18924 21364 18952
rect 21131 18921 21143 18924
rect 21085 18915 21143 18921
rect 21358 18912 21364 18924
rect 21416 18952 21422 18964
rect 26694 18952 26700 18964
rect 21416 18924 26700 18952
rect 21416 18912 21422 18924
rect 26694 18912 26700 18924
rect 26752 18912 26758 18964
rect 27617 18955 27675 18961
rect 27617 18921 27629 18955
rect 27663 18952 27675 18955
rect 27706 18952 27712 18964
rect 27663 18924 27712 18952
rect 27663 18921 27675 18924
rect 27617 18915 27675 18921
rect 27706 18912 27712 18924
rect 27764 18912 27770 18964
rect 22278 18884 22284 18896
rect 20640 18856 22284 18884
rect 22278 18844 22284 18856
rect 22336 18844 22342 18896
rect 27798 18844 27804 18896
rect 27856 18884 27862 18896
rect 27856 18856 28580 18884
rect 27856 18844 27862 18856
rect 18506 18816 18512 18828
rect 18064 18788 18512 18816
rect 18064 18757 18092 18788
rect 18506 18776 18512 18788
rect 18564 18776 18570 18828
rect 19978 18776 19984 18828
rect 20036 18816 20042 18828
rect 22462 18816 22468 18828
rect 20036 18788 22468 18816
rect 20036 18776 20042 18788
rect 22462 18776 22468 18788
rect 22520 18776 22526 18828
rect 26418 18776 26424 18828
rect 26476 18816 26482 18828
rect 26476 18788 28304 18816
rect 26476 18776 26482 18788
rect 17279 18720 17448 18748
rect 17911 18751 17969 18757
rect 17279 18717 17291 18720
rect 17233 18711 17291 18717
rect 17911 18717 17923 18751
rect 17957 18717 17969 18751
rect 17911 18711 17969 18717
rect 18049 18751 18107 18757
rect 18049 18717 18061 18751
rect 18095 18717 18107 18751
rect 18049 18711 18107 18717
rect 18138 18708 18144 18760
rect 18196 18748 18202 18760
rect 18196 18720 18241 18748
rect 18196 18708 18202 18720
rect 18322 18708 18328 18760
rect 18380 18748 18386 18760
rect 18380 18720 18425 18748
rect 18380 18708 18386 18720
rect 19150 18708 19156 18760
rect 19208 18748 19214 18760
rect 22554 18748 22560 18760
rect 19208 18720 22560 18748
rect 19208 18708 19214 18720
rect 22554 18708 22560 18720
rect 22612 18708 22618 18760
rect 23934 18708 23940 18760
rect 23992 18748 23998 18760
rect 24486 18748 24492 18760
rect 23992 18720 24492 18748
rect 23992 18708 23998 18720
rect 24486 18708 24492 18720
rect 24544 18708 24550 18760
rect 26234 18708 26240 18760
rect 26292 18748 26298 18760
rect 26878 18748 26884 18760
rect 26292 18720 26884 18748
rect 26292 18708 26298 18720
rect 26878 18708 26884 18720
rect 26936 18748 26942 18760
rect 27154 18757 27160 18760
rect 26973 18751 27031 18757
rect 26973 18748 26985 18751
rect 26936 18720 26985 18748
rect 26936 18708 26942 18720
rect 26973 18717 26985 18720
rect 27019 18717 27031 18751
rect 26973 18711 27031 18717
rect 27121 18751 27160 18757
rect 27121 18717 27133 18751
rect 27121 18711 27160 18717
rect 27154 18708 27160 18711
rect 27212 18708 27218 18760
rect 27430 18708 27436 18760
rect 27488 18757 27494 18760
rect 28276 18757 28304 18788
rect 28552 18760 28580 18856
rect 27488 18748 27496 18757
rect 28261 18751 28319 18757
rect 27488 18720 27533 18748
rect 27488 18711 27496 18720
rect 28261 18717 28273 18751
rect 28307 18717 28319 18751
rect 28261 18711 28319 18717
rect 28445 18751 28503 18757
rect 28445 18717 28457 18751
rect 28491 18717 28503 18751
rect 28445 18711 28503 18717
rect 27488 18708 27494 18711
rect 10928 18652 13308 18680
rect 14773 18680 14801 18708
rect 15194 18680 15200 18692
rect 14773 18652 15200 18680
rect 10928 18640 10934 18652
rect 15194 18640 15200 18652
rect 15252 18640 15258 18692
rect 16960 18624 16988 18708
rect 17126 18640 17132 18692
rect 17184 18680 17190 18692
rect 18506 18680 18512 18692
rect 17184 18652 18512 18680
rect 17184 18640 17190 18652
rect 18506 18640 18512 18652
rect 18564 18640 18570 18692
rect 19426 18640 19432 18692
rect 19484 18680 19490 18692
rect 19613 18683 19671 18689
rect 19613 18680 19625 18683
rect 19484 18652 19625 18680
rect 19484 18640 19490 18652
rect 19613 18649 19625 18652
rect 19659 18649 19671 18683
rect 19613 18643 19671 18649
rect 21818 18640 21824 18692
rect 21876 18680 21882 18692
rect 22710 18683 22768 18689
rect 22710 18680 22722 18683
rect 21876 18652 22722 18680
rect 21876 18640 21882 18652
rect 22710 18649 22722 18652
rect 22756 18649 22768 18683
rect 22710 18643 22768 18649
rect 24756 18683 24814 18689
rect 24756 18649 24768 18683
rect 24802 18680 24814 18683
rect 25774 18680 25780 18692
rect 24802 18652 25780 18680
rect 24802 18649 24814 18652
rect 24756 18643 24814 18649
rect 25774 18640 25780 18652
rect 25832 18640 25838 18692
rect 27249 18683 27307 18689
rect 27249 18649 27261 18683
rect 27295 18649 27307 18683
rect 27249 18643 27307 18649
rect 27341 18683 27399 18689
rect 27341 18649 27353 18683
rect 27387 18680 27399 18683
rect 27890 18680 27896 18692
rect 27387 18652 27896 18680
rect 27387 18649 27399 18652
rect 27341 18643 27399 18649
rect 12802 18612 12808 18624
rect 12763 18584 12808 18612
rect 12802 18572 12808 18584
rect 12860 18572 12866 18624
rect 14277 18615 14335 18621
rect 14277 18581 14289 18615
rect 14323 18612 14335 18615
rect 14366 18612 14372 18624
rect 14323 18584 14372 18612
rect 14323 18581 14335 18584
rect 14277 18575 14335 18581
rect 14366 18572 14372 18584
rect 14424 18572 14430 18624
rect 16574 18612 16580 18624
rect 16535 18584 16580 18612
rect 16574 18572 16580 18584
rect 16632 18572 16638 18624
rect 16942 18572 16948 18624
rect 17000 18572 17006 18624
rect 17310 18572 17316 18624
rect 17368 18612 17374 18624
rect 23658 18612 23664 18624
rect 17368 18584 23664 18612
rect 17368 18572 17374 18584
rect 23658 18572 23664 18584
rect 23716 18572 23722 18624
rect 23842 18612 23848 18624
rect 23803 18584 23848 18612
rect 23842 18572 23848 18584
rect 23900 18572 23906 18624
rect 25869 18615 25927 18621
rect 25869 18581 25881 18615
rect 25915 18612 25927 18615
rect 26234 18612 26240 18624
rect 25915 18584 26240 18612
rect 25915 18581 25927 18584
rect 25869 18575 25927 18581
rect 26234 18572 26240 18584
rect 26292 18612 26298 18624
rect 27154 18612 27160 18624
rect 26292 18584 27160 18612
rect 26292 18572 26298 18584
rect 27154 18572 27160 18584
rect 27212 18572 27218 18624
rect 27264 18612 27292 18643
rect 27890 18640 27896 18652
rect 27948 18640 27954 18692
rect 28460 18680 28488 18711
rect 28534 18708 28540 18760
rect 28592 18748 28598 18760
rect 28592 18720 28637 18748
rect 28592 18708 28598 18720
rect 28626 18680 28632 18692
rect 28460 18652 28632 18680
rect 28626 18640 28632 18652
rect 28684 18640 28690 18692
rect 27430 18612 27436 18624
rect 27264 18584 27436 18612
rect 27430 18572 27436 18584
rect 27488 18572 27494 18624
rect 28074 18612 28080 18624
rect 28035 18584 28080 18612
rect 28074 18572 28080 18584
rect 28132 18572 28138 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 10045 18411 10103 18417
rect 10045 18377 10057 18411
rect 10091 18408 10103 18411
rect 10502 18408 10508 18420
rect 10091 18380 10508 18408
rect 10091 18377 10103 18380
rect 10045 18371 10103 18377
rect 10502 18368 10508 18380
rect 10560 18408 10566 18420
rect 10560 18380 10640 18408
rect 10560 18368 10566 18380
rect 10612 18349 10640 18380
rect 10686 18368 10692 18420
rect 10744 18408 10750 18420
rect 10744 18380 10789 18408
rect 10744 18368 10750 18380
rect 13078 18368 13084 18420
rect 13136 18408 13142 18420
rect 13136 18380 19840 18408
rect 13136 18368 13142 18380
rect 10597 18343 10655 18349
rect 10597 18309 10609 18343
rect 10643 18309 10655 18343
rect 10597 18303 10655 18309
rect 16574 18300 16580 18352
rect 16632 18340 16638 18352
rect 17466 18343 17524 18349
rect 17466 18340 17478 18343
rect 16632 18312 17478 18340
rect 16632 18300 16638 18312
rect 17466 18309 17478 18312
rect 17512 18309 17524 18343
rect 19058 18340 19064 18352
rect 17466 18303 17524 18309
rect 17696 18312 19064 18340
rect 8478 18232 8484 18284
rect 8536 18272 8542 18284
rect 8665 18275 8723 18281
rect 8665 18272 8677 18275
rect 8536 18244 8677 18272
rect 8536 18232 8542 18244
rect 8665 18241 8677 18244
rect 8711 18241 8723 18275
rect 8665 18235 8723 18241
rect 8932 18275 8990 18281
rect 8932 18241 8944 18275
rect 8978 18272 8990 18275
rect 8978 18244 10548 18272
rect 8978 18241 8990 18244
rect 8932 18235 8990 18241
rect 10520 18204 10548 18244
rect 10962 18232 10968 18284
rect 11020 18272 11026 18284
rect 11517 18275 11575 18281
rect 11517 18272 11529 18275
rect 11020 18244 11529 18272
rect 11020 18232 11026 18244
rect 11517 18241 11529 18244
rect 11563 18241 11575 18275
rect 13078 18272 13084 18284
rect 13039 18244 13084 18272
rect 11517 18235 11575 18241
rect 13078 18232 13084 18244
rect 13136 18232 13142 18284
rect 13173 18275 13231 18281
rect 13173 18241 13185 18275
rect 13219 18241 13231 18275
rect 13173 18235 13231 18241
rect 12805 18207 12863 18213
rect 12805 18204 12817 18207
rect 10520 18176 12817 18204
rect 12805 18173 12817 18176
rect 12851 18173 12863 18207
rect 13188 18204 13216 18235
rect 13262 18232 13268 18284
rect 13320 18272 13326 18284
rect 13449 18275 13507 18281
rect 13320 18244 13365 18272
rect 13320 18232 13326 18244
rect 13449 18241 13461 18275
rect 13495 18272 13507 18275
rect 13538 18272 13544 18284
rect 13495 18244 13544 18272
rect 13495 18241 13507 18244
rect 13449 18235 13507 18241
rect 13538 18232 13544 18244
rect 13596 18232 13602 18284
rect 14182 18272 14188 18284
rect 14143 18244 14188 18272
rect 14182 18232 14188 18244
rect 14240 18232 14246 18284
rect 14277 18275 14335 18281
rect 14277 18241 14289 18275
rect 14323 18241 14335 18275
rect 14277 18235 14335 18241
rect 14369 18275 14427 18281
rect 14369 18241 14381 18275
rect 14415 18272 14427 18275
rect 14458 18272 14464 18284
rect 14415 18244 14464 18272
rect 14415 18241 14427 18244
rect 14369 18235 14427 18241
rect 13814 18204 13820 18216
rect 13188 18176 13820 18204
rect 12805 18167 12863 18173
rect 13814 18164 13820 18176
rect 13872 18204 13878 18216
rect 14292 18204 14320 18235
rect 14458 18232 14464 18244
rect 14516 18232 14522 18284
rect 14550 18232 14556 18284
rect 14608 18272 14614 18284
rect 15197 18275 15255 18281
rect 14608 18244 14653 18272
rect 14608 18232 14614 18244
rect 15197 18241 15209 18275
rect 15243 18272 15255 18275
rect 15470 18272 15476 18284
rect 15243 18244 15476 18272
rect 15243 18241 15255 18244
rect 15197 18235 15255 18241
rect 15470 18232 15476 18244
rect 15528 18232 15534 18284
rect 15746 18272 15752 18284
rect 15707 18244 15752 18272
rect 15746 18232 15752 18244
rect 15804 18232 15810 18284
rect 17696 18272 17724 18312
rect 19058 18300 19064 18312
rect 19116 18300 19122 18352
rect 19812 18340 19840 18380
rect 22002 18368 22008 18420
rect 22060 18408 22066 18420
rect 26786 18408 26792 18420
rect 22060 18380 23704 18408
rect 22060 18368 22066 18380
rect 20064 18343 20122 18349
rect 19812 18312 20024 18340
rect 17052 18244 17724 18272
rect 19797 18275 19855 18281
rect 16022 18204 16028 18216
rect 13872 18176 14320 18204
rect 15983 18176 16028 18204
rect 13872 18164 13878 18176
rect 16022 18164 16028 18176
rect 16080 18164 16086 18216
rect 15289 18139 15347 18145
rect 15289 18105 15301 18139
rect 15335 18136 15347 18139
rect 17052 18136 17080 18244
rect 19797 18241 19809 18275
rect 19843 18272 19855 18275
rect 19886 18272 19892 18284
rect 19843 18244 19892 18272
rect 19843 18241 19855 18244
rect 19797 18235 19855 18241
rect 19886 18232 19892 18244
rect 19944 18232 19950 18284
rect 19996 18272 20024 18312
rect 20064 18309 20076 18343
rect 20110 18340 20122 18343
rect 20438 18340 20444 18352
rect 20110 18312 20444 18340
rect 20110 18309 20122 18312
rect 20064 18303 20122 18309
rect 20438 18300 20444 18312
rect 20496 18300 20502 18352
rect 22094 18300 22100 18352
rect 22152 18340 22158 18352
rect 22922 18340 22928 18352
rect 22152 18312 22928 18340
rect 22152 18300 22158 18312
rect 22922 18300 22928 18312
rect 22980 18340 22986 18352
rect 22980 18312 23336 18340
rect 22980 18300 22986 18312
rect 22830 18272 22836 18284
rect 19996 18244 22836 18272
rect 22830 18232 22836 18244
rect 22888 18232 22894 18284
rect 23106 18272 23112 18284
rect 23067 18244 23112 18272
rect 23106 18232 23112 18244
rect 23164 18232 23170 18284
rect 23308 18281 23336 18312
rect 23676 18281 23704 18380
rect 25884 18380 26792 18408
rect 25314 18340 25320 18352
rect 24320 18312 25320 18340
rect 24320 18281 24348 18312
rect 25314 18300 25320 18312
rect 25372 18340 25378 18352
rect 25372 18312 25821 18340
rect 25372 18300 25378 18312
rect 23293 18275 23351 18281
rect 23293 18241 23305 18275
rect 23339 18241 23351 18275
rect 23293 18235 23351 18241
rect 23661 18275 23719 18281
rect 23661 18241 23673 18275
rect 23707 18241 23719 18275
rect 24305 18275 24363 18281
rect 24305 18272 24317 18275
rect 23661 18235 23719 18241
rect 23768 18244 24317 18272
rect 17218 18204 17224 18216
rect 17179 18176 17224 18204
rect 17218 18164 17224 18176
rect 17276 18164 17282 18216
rect 21821 18207 21879 18213
rect 21821 18204 21833 18207
rect 20824 18176 21833 18204
rect 15335 18108 17080 18136
rect 15335 18105 15347 18108
rect 15289 18099 15347 18105
rect 18690 18096 18696 18148
rect 18748 18136 18754 18148
rect 18748 18108 19840 18136
rect 18748 18096 18754 18108
rect 11701 18071 11759 18077
rect 11701 18037 11713 18071
rect 11747 18068 11759 18071
rect 12342 18068 12348 18080
rect 11747 18040 12348 18068
rect 11747 18037 11759 18040
rect 11701 18031 11759 18037
rect 12342 18028 12348 18040
rect 12400 18028 12406 18080
rect 13909 18071 13967 18077
rect 13909 18037 13921 18071
rect 13955 18068 13967 18071
rect 14182 18068 14188 18080
rect 13955 18040 14188 18068
rect 13955 18037 13967 18040
rect 13909 18031 13967 18037
rect 14182 18028 14188 18040
rect 14240 18028 14246 18080
rect 16850 18028 16856 18080
rect 16908 18068 16914 18080
rect 18230 18068 18236 18080
rect 16908 18040 18236 18068
rect 16908 18028 16914 18040
rect 18230 18028 18236 18040
rect 18288 18068 18294 18080
rect 18601 18071 18659 18077
rect 18601 18068 18613 18071
rect 18288 18040 18613 18068
rect 18288 18028 18294 18040
rect 18601 18037 18613 18040
rect 18647 18068 18659 18071
rect 18782 18068 18788 18080
rect 18647 18040 18788 18068
rect 18647 18037 18659 18040
rect 18601 18031 18659 18037
rect 18782 18028 18788 18040
rect 18840 18028 18846 18080
rect 19812 18068 19840 18108
rect 20438 18068 20444 18080
rect 19812 18040 20444 18068
rect 20438 18028 20444 18040
rect 20496 18068 20502 18080
rect 20824 18068 20852 18176
rect 21821 18173 21833 18176
rect 21867 18173 21879 18207
rect 21821 18167 21879 18173
rect 21910 18164 21916 18216
rect 21968 18204 21974 18216
rect 22097 18207 22155 18213
rect 22097 18204 22109 18207
rect 21968 18176 22109 18204
rect 21968 18164 21974 18176
rect 22097 18173 22109 18176
rect 22143 18173 22155 18207
rect 22848 18204 22876 18232
rect 23385 18207 23443 18213
rect 23385 18204 23397 18207
rect 22848 18176 23397 18204
rect 22097 18167 22155 18173
rect 23385 18173 23397 18176
rect 23431 18173 23443 18207
rect 23385 18167 23443 18173
rect 20990 18096 20996 18148
rect 21048 18136 21054 18148
rect 21266 18136 21272 18148
rect 21048 18108 21272 18136
rect 21048 18096 21054 18108
rect 21266 18096 21272 18108
rect 21324 18096 21330 18148
rect 22112 18136 22140 18167
rect 23474 18164 23480 18216
rect 23532 18204 23538 18216
rect 23532 18176 23577 18204
rect 23532 18164 23538 18176
rect 23768 18136 23796 18244
rect 24305 18241 24317 18244
rect 24351 18241 24363 18275
rect 24305 18235 24363 18241
rect 24489 18275 24547 18281
rect 24489 18241 24501 18275
rect 24535 18272 24547 18275
rect 24762 18272 24768 18284
rect 24535 18244 24768 18272
rect 24535 18241 24547 18244
rect 24489 18235 24547 18241
rect 24762 18232 24768 18244
rect 24820 18232 24826 18284
rect 24857 18275 24915 18281
rect 24857 18241 24869 18275
rect 24903 18272 24915 18275
rect 25038 18272 25044 18284
rect 24903 18244 25044 18272
rect 24903 18241 24915 18244
rect 24857 18235 24915 18241
rect 25038 18232 25044 18244
rect 25096 18232 25102 18284
rect 25689 18275 25747 18281
rect 25689 18241 25701 18275
rect 25735 18274 25747 18275
rect 25793 18274 25821 18312
rect 25884 18281 25912 18380
rect 26786 18368 26792 18380
rect 26844 18368 26850 18420
rect 26421 18343 26479 18349
rect 26421 18309 26433 18343
rect 26467 18340 26479 18343
rect 26467 18312 29040 18340
rect 26467 18309 26479 18312
rect 26421 18303 26479 18309
rect 25735 18246 25821 18274
rect 25857 18275 25915 18281
rect 25735 18241 25747 18246
rect 25689 18235 25747 18241
rect 25857 18241 25869 18275
rect 25903 18241 25915 18275
rect 25857 18235 25915 18241
rect 25961 18275 26019 18281
rect 25961 18241 25973 18275
rect 26007 18272 26019 18275
rect 26237 18275 26295 18281
rect 26007 18244 26188 18272
rect 26007 18241 26019 18244
rect 25961 18235 26019 18241
rect 26160 18216 26188 18244
rect 26237 18241 26249 18275
rect 26283 18272 26295 18275
rect 26326 18272 26332 18284
rect 26283 18244 26332 18272
rect 26283 18241 26295 18244
rect 26237 18235 26295 18241
rect 26326 18232 26332 18244
rect 26384 18232 26390 18284
rect 29012 18281 29040 18312
rect 27240 18275 27298 18281
rect 27240 18241 27252 18275
rect 27286 18272 27298 18275
rect 28813 18275 28871 18281
rect 28813 18272 28825 18275
rect 27286 18244 28825 18272
rect 27286 18241 27298 18244
rect 27240 18235 27298 18241
rect 28813 18241 28825 18244
rect 28859 18241 28871 18275
rect 28813 18235 28871 18241
rect 28997 18275 29055 18281
rect 28997 18241 29009 18275
rect 29043 18241 29055 18275
rect 28997 18235 29055 18241
rect 24210 18164 24216 18216
rect 24268 18204 24274 18216
rect 24581 18207 24639 18213
rect 24581 18204 24593 18207
rect 24268 18176 24593 18204
rect 24268 18164 24274 18176
rect 24581 18173 24593 18176
rect 24627 18173 24639 18207
rect 24581 18167 24639 18173
rect 24673 18207 24731 18213
rect 24673 18173 24685 18207
rect 24719 18204 24731 18207
rect 25590 18204 25596 18216
rect 24719 18176 25596 18204
rect 24719 18173 24731 18176
rect 24673 18167 24731 18173
rect 25590 18164 25596 18176
rect 25648 18204 25654 18216
rect 26053 18207 26111 18213
rect 26053 18204 26065 18207
rect 25648 18176 26065 18204
rect 25648 18164 25654 18176
rect 26053 18173 26065 18176
rect 26099 18173 26111 18207
rect 26053 18167 26111 18173
rect 26142 18164 26148 18216
rect 26200 18164 26206 18216
rect 26970 18204 26976 18216
rect 26883 18176 26976 18204
rect 26970 18164 26976 18176
rect 27028 18164 27034 18216
rect 28350 18204 28356 18216
rect 28263 18176 28356 18204
rect 28350 18164 28356 18176
rect 28408 18204 28414 18216
rect 29273 18207 29331 18213
rect 29273 18204 29285 18207
rect 28408 18176 29285 18204
rect 28408 18164 28414 18176
rect 29273 18173 29285 18176
rect 29319 18173 29331 18207
rect 29273 18167 29331 18173
rect 22112 18108 23796 18136
rect 24486 18096 24492 18148
rect 24544 18136 24550 18148
rect 26988 18136 27016 18164
rect 24544 18108 27016 18136
rect 24544 18096 24550 18108
rect 21174 18068 21180 18080
rect 20496 18040 20852 18068
rect 21135 18040 21180 18068
rect 20496 18028 20502 18040
rect 21174 18028 21180 18040
rect 21232 18028 21238 18080
rect 22094 18028 22100 18080
rect 22152 18068 22158 18080
rect 23845 18071 23903 18077
rect 23845 18068 23857 18071
rect 22152 18040 23857 18068
rect 22152 18028 22158 18040
rect 23845 18037 23857 18040
rect 23891 18037 23903 18071
rect 23845 18031 23903 18037
rect 25041 18071 25099 18077
rect 25041 18037 25053 18071
rect 25087 18068 25099 18071
rect 27246 18068 27252 18080
rect 25087 18040 27252 18068
rect 25087 18037 25099 18040
rect 25041 18031 25099 18037
rect 27246 18028 27252 18040
rect 27304 18028 27310 18080
rect 28258 18028 28264 18080
rect 28316 18068 28322 18080
rect 28368 18077 28396 18164
rect 28353 18071 28411 18077
rect 28353 18068 28365 18071
rect 28316 18040 28365 18068
rect 28316 18028 28322 18040
rect 28353 18037 28365 18040
rect 28399 18037 28411 18071
rect 28353 18031 28411 18037
rect 28626 18028 28632 18080
rect 28684 18068 28690 18080
rect 29181 18071 29239 18077
rect 29181 18068 29193 18071
rect 28684 18040 29193 18068
rect 28684 18028 28690 18040
rect 29181 18037 29193 18040
rect 29227 18037 29239 18071
rect 29181 18031 29239 18037
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 10321 17867 10379 17873
rect 10321 17833 10333 17867
rect 10367 17864 10379 17867
rect 10410 17864 10416 17876
rect 10367 17836 10416 17864
rect 10367 17833 10379 17836
rect 10321 17827 10379 17833
rect 10410 17824 10416 17836
rect 10468 17864 10474 17876
rect 10962 17864 10968 17876
rect 10468 17836 10968 17864
rect 10468 17824 10474 17836
rect 10962 17824 10968 17836
rect 11020 17824 11026 17876
rect 15470 17824 15476 17876
rect 15528 17864 15534 17876
rect 16390 17864 16396 17876
rect 15528 17836 16396 17864
rect 15528 17824 15534 17836
rect 16390 17824 16396 17836
rect 16448 17824 16454 17876
rect 17954 17864 17960 17876
rect 17926 17824 17960 17864
rect 18012 17824 18018 17876
rect 19981 17867 20039 17873
rect 18340 17836 18516 17864
rect 15562 17756 15568 17808
rect 15620 17796 15626 17808
rect 16482 17796 16488 17808
rect 15620 17768 16488 17796
rect 15620 17756 15626 17768
rect 16482 17756 16488 17768
rect 16540 17796 16546 17808
rect 17926 17796 17954 17824
rect 18340 17796 18368 17836
rect 16540 17768 16620 17796
rect 16540 17756 16546 17768
rect 8478 17688 8484 17740
rect 8536 17728 8542 17740
rect 8941 17731 8999 17737
rect 8941 17728 8953 17731
rect 8536 17700 8953 17728
rect 8536 17688 8542 17700
rect 8941 17697 8953 17700
rect 8987 17697 8999 17731
rect 12802 17728 12808 17740
rect 8941 17691 8999 17697
rect 10796 17700 12808 17728
rect 9208 17663 9266 17669
rect 9208 17629 9220 17663
rect 9254 17660 9266 17663
rect 10796 17660 10824 17700
rect 12802 17688 12808 17700
rect 12860 17688 12866 17740
rect 15838 17688 15844 17740
rect 15896 17728 15902 17740
rect 16390 17728 16396 17740
rect 15896 17700 16396 17728
rect 15896 17688 15902 17700
rect 16390 17688 16396 17700
rect 16448 17728 16454 17740
rect 16448 17700 16528 17728
rect 16448 17688 16454 17700
rect 9254 17632 10824 17660
rect 11149 17663 11207 17669
rect 9254 17629 9266 17632
rect 9208 17623 9266 17629
rect 11149 17629 11161 17663
rect 11195 17660 11207 17663
rect 11195 17632 11744 17660
rect 11195 17629 11207 17632
rect 11149 17623 11207 17629
rect 11716 17601 11744 17632
rect 11790 17620 11796 17672
rect 11848 17660 11854 17672
rect 12250 17660 12256 17672
rect 11848 17632 12256 17660
rect 11848 17620 11854 17632
rect 12250 17620 12256 17632
rect 12308 17620 12314 17672
rect 13170 17660 13176 17672
rect 13131 17632 13176 17660
rect 13170 17620 13176 17632
rect 13228 17620 13234 17672
rect 13265 17663 13323 17669
rect 13265 17629 13277 17663
rect 13311 17629 13323 17663
rect 13265 17623 13323 17629
rect 11701 17595 11759 17601
rect 11701 17561 11713 17595
rect 11747 17592 11759 17595
rect 11974 17592 11980 17604
rect 11747 17564 11980 17592
rect 11747 17561 11759 17564
rect 11701 17555 11759 17561
rect 11974 17552 11980 17564
rect 12032 17552 12038 17604
rect 13280 17592 13308 17623
rect 13354 17620 13360 17672
rect 13412 17660 13418 17672
rect 13412 17632 13457 17660
rect 13412 17620 13418 17632
rect 13538 17620 13544 17672
rect 13596 17660 13602 17672
rect 14090 17660 14096 17672
rect 13596 17632 13952 17660
rect 14051 17632 14096 17660
rect 13596 17620 13602 17632
rect 13814 17592 13820 17604
rect 13280 17564 13820 17592
rect 13814 17552 13820 17564
rect 13872 17552 13878 17604
rect 13924 17592 13952 17632
rect 14090 17620 14096 17632
rect 14148 17620 14154 17672
rect 14182 17620 14188 17672
rect 14240 17660 14246 17672
rect 14349 17663 14407 17669
rect 14349 17660 14361 17663
rect 14240 17632 14361 17660
rect 14240 17620 14246 17632
rect 14349 17629 14361 17632
rect 14395 17629 14407 17663
rect 14349 17623 14407 17629
rect 16022 17620 16028 17672
rect 16080 17660 16086 17672
rect 16500 17669 16528 17700
rect 16592 17669 16620 17768
rect 17328 17768 17954 17796
rect 18156 17768 18368 17796
rect 16209 17663 16267 17669
rect 16209 17660 16221 17663
rect 16080 17632 16221 17660
rect 16080 17620 16086 17632
rect 16209 17629 16221 17632
rect 16255 17629 16267 17663
rect 16209 17623 16267 17629
rect 16301 17663 16359 17669
rect 16301 17629 16313 17663
rect 16347 17629 16359 17663
rect 16301 17623 16359 17629
rect 16485 17663 16543 17669
rect 16485 17629 16497 17663
rect 16531 17629 16543 17663
rect 16485 17623 16543 17629
rect 16577 17663 16635 17669
rect 16577 17629 16589 17663
rect 16623 17629 16635 17663
rect 16577 17623 16635 17629
rect 17221 17663 17279 17669
rect 17221 17629 17233 17663
rect 17267 17660 17279 17663
rect 17328 17660 17356 17768
rect 17405 17731 17463 17737
rect 17405 17697 17417 17731
rect 17451 17728 17463 17731
rect 17862 17728 17868 17740
rect 17451 17700 17868 17728
rect 17451 17697 17463 17700
rect 17405 17691 17463 17697
rect 17862 17688 17868 17700
rect 17920 17688 17926 17740
rect 17267 17632 17356 17660
rect 17497 17663 17555 17669
rect 17267 17629 17279 17632
rect 17221 17623 17279 17629
rect 17497 17629 17509 17663
rect 17543 17660 17555 17663
rect 17770 17660 17776 17672
rect 17543 17632 17776 17660
rect 17543 17629 17555 17632
rect 17497 17623 17555 17629
rect 14918 17592 14924 17604
rect 13924 17564 14924 17592
rect 14918 17552 14924 17564
rect 14976 17552 14982 17604
rect 16316 17592 16344 17623
rect 17770 17620 17776 17632
rect 17828 17620 17834 17672
rect 17954 17620 17960 17672
rect 18012 17660 18018 17672
rect 18156 17669 18184 17768
rect 18322 17688 18328 17740
rect 18380 17728 18386 17740
rect 18488 17728 18516 17836
rect 19981 17833 19993 17867
rect 20027 17864 20039 17867
rect 20622 17864 20628 17876
rect 20027 17836 20628 17864
rect 20027 17833 20039 17836
rect 19981 17827 20039 17833
rect 20622 17824 20628 17836
rect 20680 17824 20686 17876
rect 21818 17864 21824 17876
rect 21779 17836 21824 17864
rect 21818 17824 21824 17836
rect 21876 17824 21882 17876
rect 22189 17867 22247 17873
rect 22189 17833 22201 17867
rect 22235 17864 22247 17867
rect 23290 17864 23296 17876
rect 22235 17836 23296 17864
rect 22235 17833 22247 17836
rect 22189 17827 22247 17833
rect 23290 17824 23296 17836
rect 23348 17824 23354 17876
rect 23474 17824 23480 17876
rect 23532 17864 23538 17876
rect 26418 17864 26424 17876
rect 23532 17836 24799 17864
rect 26379 17836 26424 17864
rect 23532 17824 23538 17836
rect 19426 17756 19432 17808
rect 19484 17756 19490 17808
rect 19518 17756 19524 17808
rect 19576 17796 19582 17808
rect 20162 17796 20168 17808
rect 19576 17768 20168 17796
rect 19576 17756 19582 17768
rect 20162 17756 20168 17768
rect 20220 17796 20226 17808
rect 20220 17768 20852 17796
rect 20220 17756 20226 17768
rect 19460 17728 19488 17756
rect 18380 17700 18425 17728
rect 18488 17700 19488 17728
rect 18380 17688 18386 17700
rect 18141 17663 18199 17669
rect 18012 17632 18057 17660
rect 18012 17620 18018 17632
rect 18141 17629 18153 17663
rect 18187 17629 18199 17663
rect 18141 17623 18199 17629
rect 18230 17620 18236 17672
rect 18288 17660 18294 17672
rect 18509 17663 18567 17669
rect 18288 17632 18333 17660
rect 18288 17620 18294 17632
rect 18509 17629 18521 17663
rect 18555 17660 18567 17663
rect 18874 17660 18880 17672
rect 18555 17632 18880 17660
rect 18555 17629 18567 17632
rect 18509 17623 18567 17629
rect 18874 17620 18880 17632
rect 18932 17620 18938 17672
rect 19242 17660 19248 17672
rect 19203 17632 19248 17660
rect 19242 17620 19248 17632
rect 19300 17620 19306 17672
rect 19460 17669 19488 17700
rect 19613 17731 19671 17737
rect 19613 17697 19625 17731
rect 19659 17728 19671 17731
rect 19978 17728 19984 17740
rect 19659 17700 19984 17728
rect 19659 17697 19671 17700
rect 19613 17691 19671 17697
rect 19978 17688 19984 17700
rect 20036 17728 20042 17740
rect 20254 17728 20260 17740
rect 20036 17700 20260 17728
rect 20036 17688 20042 17700
rect 20254 17688 20260 17700
rect 20312 17728 20318 17740
rect 20824 17737 20852 17768
rect 23198 17756 23204 17808
rect 23256 17796 23262 17808
rect 23842 17796 23848 17808
rect 23256 17768 23848 17796
rect 23256 17756 23262 17768
rect 23842 17756 23848 17768
rect 23900 17756 23906 17808
rect 20809 17731 20867 17737
rect 20312 17700 20668 17728
rect 20312 17688 20318 17700
rect 19433 17663 19491 17669
rect 19433 17660 19445 17663
rect 19355 17632 19445 17660
rect 19433 17629 19445 17632
rect 19479 17629 19491 17663
rect 19433 17623 19491 17629
rect 19521 17663 19579 17669
rect 19521 17629 19533 17663
rect 19567 17658 19579 17663
rect 19702 17660 19708 17672
rect 19628 17658 19708 17660
rect 19567 17632 19708 17658
rect 19567 17630 19656 17632
rect 19567 17629 19579 17630
rect 19521 17623 19579 17629
rect 15856 17564 16344 17592
rect 17037 17595 17095 17601
rect 15856 17536 15884 17564
rect 17037 17561 17049 17595
rect 17083 17592 17095 17595
rect 19460 17592 19488 17623
rect 19702 17620 19708 17632
rect 19760 17620 19766 17672
rect 19797 17663 19855 17669
rect 19797 17629 19809 17663
rect 19843 17662 19855 17663
rect 19843 17660 19923 17662
rect 20346 17660 20352 17672
rect 19843 17634 20352 17660
rect 19843 17629 19855 17634
rect 19895 17632 20352 17634
rect 19797 17623 19855 17629
rect 20346 17620 20352 17632
rect 20404 17620 20410 17672
rect 20438 17620 20444 17672
rect 20496 17660 20502 17672
rect 20533 17663 20591 17669
rect 20533 17660 20545 17663
rect 20496 17632 20545 17660
rect 20496 17620 20502 17632
rect 20533 17629 20545 17632
rect 20579 17629 20591 17663
rect 20640 17660 20668 17700
rect 20809 17697 20821 17731
rect 20855 17728 20867 17731
rect 24670 17728 24676 17740
rect 20855 17700 23152 17728
rect 24631 17700 24676 17728
rect 20855 17697 20867 17700
rect 20809 17691 20867 17697
rect 23124 17672 23152 17700
rect 24670 17688 24676 17700
rect 24728 17688 24734 17740
rect 24771 17737 24799 17836
rect 26418 17824 26424 17836
rect 26476 17824 26482 17876
rect 25590 17756 25596 17808
rect 25648 17796 25654 17808
rect 25648 17768 26096 17796
rect 25648 17756 25654 17768
rect 24765 17731 24823 17737
rect 24765 17697 24777 17731
rect 24811 17697 24823 17731
rect 24765 17691 24823 17697
rect 25498 17688 25504 17740
rect 25556 17728 25562 17740
rect 25961 17731 26019 17737
rect 25961 17728 25973 17731
rect 25556 17700 25973 17728
rect 25556 17688 25562 17700
rect 25961 17697 25973 17700
rect 26007 17697 26019 17731
rect 25961 17691 26019 17697
rect 21450 17660 21456 17672
rect 20640 17632 21456 17660
rect 20533 17623 20591 17629
rect 21450 17620 21456 17632
rect 21508 17620 21514 17672
rect 22005 17663 22063 17669
rect 22005 17629 22017 17663
rect 22051 17660 22063 17663
rect 22094 17660 22100 17672
rect 22051 17632 22100 17660
rect 22051 17629 22063 17632
rect 22005 17623 22063 17629
rect 22094 17620 22100 17632
rect 22152 17620 22158 17672
rect 22278 17660 22284 17672
rect 22239 17632 22284 17660
rect 22278 17620 22284 17632
rect 22336 17620 22342 17672
rect 22554 17620 22560 17672
rect 22612 17660 22618 17672
rect 22741 17663 22799 17669
rect 22741 17660 22753 17663
rect 22612 17632 22753 17660
rect 22612 17620 22618 17632
rect 22741 17629 22753 17632
rect 22787 17629 22799 17663
rect 22741 17623 22799 17629
rect 22922 17620 22928 17672
rect 22980 17660 22986 17672
rect 23017 17663 23075 17669
rect 23017 17660 23029 17663
rect 22980 17632 23029 17660
rect 22980 17620 22986 17632
rect 23017 17629 23029 17632
rect 23063 17629 23075 17663
rect 23017 17623 23075 17629
rect 23032 17592 23060 17623
rect 23106 17620 23112 17672
rect 23164 17660 23170 17672
rect 24397 17663 24455 17669
rect 24397 17660 24409 17663
rect 23164 17632 24409 17660
rect 23164 17620 23170 17632
rect 24397 17629 24409 17632
rect 24443 17629 24455 17663
rect 24397 17623 24455 17629
rect 24581 17663 24639 17669
rect 24581 17629 24593 17663
rect 24627 17660 24639 17663
rect 24854 17660 24860 17672
rect 24627 17632 24860 17660
rect 24627 17629 24639 17632
rect 24581 17623 24639 17629
rect 24596 17592 24624 17623
rect 24854 17620 24860 17632
rect 24912 17620 24918 17672
rect 24946 17620 24952 17672
rect 25004 17660 25010 17672
rect 25004 17632 25049 17660
rect 25004 17620 25010 17632
rect 25314 17620 25320 17672
rect 25372 17660 25378 17672
rect 25685 17663 25743 17669
rect 25685 17660 25697 17663
rect 25372 17632 25697 17660
rect 25372 17620 25378 17632
rect 25685 17629 25697 17632
rect 25731 17629 25743 17663
rect 25685 17623 25743 17629
rect 25866 17620 25872 17672
rect 25924 17669 25930 17672
rect 26068 17669 26096 17768
rect 26142 17756 26148 17808
rect 26200 17796 26206 17808
rect 27062 17796 27068 17808
rect 26200 17768 27068 17796
rect 26200 17756 26206 17768
rect 27062 17756 27068 17768
rect 27120 17756 27126 17808
rect 26970 17688 26976 17740
rect 27028 17728 27034 17740
rect 27433 17731 27491 17737
rect 27433 17728 27445 17731
rect 27028 17700 27445 17728
rect 27028 17688 27034 17700
rect 27433 17697 27445 17700
rect 27479 17697 27491 17731
rect 27433 17691 27491 17697
rect 25924 17660 25931 17669
rect 26053 17663 26111 17669
rect 25924 17632 25969 17660
rect 25924 17623 25931 17632
rect 26053 17629 26065 17663
rect 26099 17660 26111 17663
rect 26142 17660 26148 17672
rect 26099 17632 26148 17660
rect 26099 17629 26111 17632
rect 26053 17623 26111 17629
rect 25924 17620 25930 17623
rect 26142 17620 26148 17632
rect 26200 17620 26206 17672
rect 26237 17663 26295 17669
rect 26237 17629 26249 17663
rect 26283 17629 26295 17663
rect 26237 17623 26295 17629
rect 17083 17564 19380 17592
rect 19460 17564 20392 17592
rect 23032 17564 24624 17592
rect 26252 17592 26280 17623
rect 26510 17620 26516 17672
rect 26568 17660 26574 17672
rect 27522 17660 27528 17672
rect 26568 17632 27528 17660
rect 26568 17620 26574 17632
rect 27522 17620 27528 17632
rect 27580 17620 27586 17672
rect 27700 17663 27758 17669
rect 27700 17629 27712 17663
rect 27746 17660 27758 17663
rect 28074 17660 28080 17672
rect 27746 17632 28080 17660
rect 27746 17629 27758 17632
rect 27700 17623 27758 17629
rect 28074 17620 28080 17632
rect 28132 17620 28138 17672
rect 28166 17592 28172 17604
rect 26252 17564 28172 17592
rect 17083 17561 17095 17564
rect 17037 17555 17095 17561
rect 19352 17536 19380 17564
rect 20364 17536 20392 17564
rect 28166 17552 28172 17564
rect 28224 17552 28230 17604
rect 10778 17484 10784 17536
rect 10836 17524 10842 17536
rect 10965 17527 11023 17533
rect 10965 17524 10977 17527
rect 10836 17496 10977 17524
rect 10836 17484 10842 17496
rect 10965 17493 10977 17496
rect 11011 17493 11023 17527
rect 11790 17524 11796 17536
rect 11751 17496 11796 17524
rect 10965 17487 11023 17493
rect 11790 17484 11796 17496
rect 11848 17484 11854 17536
rect 11882 17484 11888 17536
rect 11940 17524 11946 17536
rect 12897 17527 12955 17533
rect 12897 17524 12909 17527
rect 11940 17496 12909 17524
rect 11940 17484 11946 17496
rect 12897 17493 12909 17496
rect 12943 17493 12955 17527
rect 12897 17487 12955 17493
rect 15473 17527 15531 17533
rect 15473 17493 15485 17527
rect 15519 17524 15531 17527
rect 15838 17524 15844 17536
rect 15519 17496 15844 17524
rect 15519 17493 15531 17496
rect 15473 17487 15531 17493
rect 15838 17484 15844 17496
rect 15896 17484 15902 17536
rect 16025 17527 16083 17533
rect 16025 17493 16037 17527
rect 16071 17524 16083 17527
rect 18598 17524 18604 17536
rect 16071 17496 18604 17524
rect 16071 17493 16083 17496
rect 16025 17487 16083 17493
rect 18598 17484 18604 17496
rect 18656 17484 18662 17536
rect 18693 17527 18751 17533
rect 18693 17493 18705 17527
rect 18739 17524 18751 17527
rect 19242 17524 19248 17536
rect 18739 17496 19248 17524
rect 18739 17493 18751 17496
rect 18693 17487 18751 17493
rect 19242 17484 19248 17496
rect 19300 17484 19306 17536
rect 19334 17484 19340 17536
rect 19392 17484 19398 17536
rect 20346 17484 20352 17536
rect 20404 17484 20410 17536
rect 22738 17484 22744 17536
rect 22796 17524 22802 17536
rect 25133 17527 25191 17533
rect 25133 17524 25145 17527
rect 22796 17496 25145 17524
rect 22796 17484 22802 17496
rect 25133 17493 25145 17496
rect 25179 17493 25191 17527
rect 25133 17487 25191 17493
rect 25314 17484 25320 17536
rect 25372 17524 25378 17536
rect 25958 17524 25964 17536
rect 25372 17496 25964 17524
rect 25372 17484 25378 17496
rect 25958 17484 25964 17496
rect 26016 17524 26022 17536
rect 27614 17524 27620 17536
rect 26016 17496 27620 17524
rect 26016 17484 26022 17496
rect 27614 17484 27620 17496
rect 27672 17484 27678 17536
rect 27706 17484 27712 17536
rect 27764 17524 27770 17536
rect 28534 17524 28540 17536
rect 27764 17496 28540 17524
rect 27764 17484 27770 17496
rect 28534 17484 28540 17496
rect 28592 17524 28598 17536
rect 28813 17527 28871 17533
rect 28813 17524 28825 17527
rect 28592 17496 28825 17524
rect 28592 17484 28598 17496
rect 28813 17493 28825 17496
rect 28859 17493 28871 17527
rect 28813 17487 28871 17493
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 10321 17323 10379 17329
rect 10321 17289 10333 17323
rect 10367 17320 10379 17323
rect 10594 17320 10600 17332
rect 10367 17292 10600 17320
rect 10367 17289 10379 17292
rect 10321 17283 10379 17289
rect 10594 17280 10600 17292
rect 10652 17280 10658 17332
rect 12713 17323 12771 17329
rect 12713 17289 12725 17323
rect 12759 17320 12771 17323
rect 13354 17320 13360 17332
rect 12759 17292 13360 17320
rect 12759 17289 12771 17292
rect 12713 17283 12771 17289
rect 13354 17280 13360 17292
rect 13412 17280 13418 17332
rect 15654 17280 15660 17332
rect 15712 17320 15718 17332
rect 15841 17323 15899 17329
rect 15841 17320 15853 17323
rect 15712 17292 15853 17320
rect 15712 17280 15718 17292
rect 15841 17289 15853 17292
rect 15887 17289 15899 17323
rect 15841 17283 15899 17289
rect 16025 17323 16083 17329
rect 16025 17289 16037 17323
rect 16071 17289 16083 17323
rect 20898 17320 20904 17332
rect 16025 17283 16083 17289
rect 17926 17292 20668 17320
rect 20859 17292 20904 17320
rect 8478 17252 8484 17264
rect 7852 17224 8484 17252
rect 7852 17193 7880 17224
rect 8478 17212 8484 17224
rect 8536 17212 8542 17264
rect 11977 17255 12035 17261
rect 11977 17221 11989 17255
rect 12023 17252 12035 17255
rect 13262 17252 13268 17264
rect 12023 17224 13268 17252
rect 12023 17221 12035 17224
rect 11977 17215 12035 17221
rect 13262 17212 13268 17224
rect 13320 17212 13326 17264
rect 15102 17212 15108 17264
rect 15160 17252 15166 17264
rect 16040 17252 16068 17283
rect 17926 17252 17954 17292
rect 15160 17224 16068 17252
rect 16132 17224 17954 17252
rect 15160 17212 15166 17224
rect 7837 17187 7895 17193
rect 7837 17153 7849 17187
rect 7883 17153 7895 17187
rect 7837 17147 7895 17153
rect 7926 17144 7932 17196
rect 7984 17184 7990 17196
rect 8093 17187 8151 17193
rect 8093 17184 8105 17187
rect 7984 17156 8105 17184
rect 7984 17144 7990 17156
rect 8093 17153 8105 17156
rect 8139 17153 8151 17187
rect 10502 17184 10508 17196
rect 10463 17156 10508 17184
rect 8093 17147 8151 17153
rect 10502 17144 10508 17156
rect 10560 17144 10566 17196
rect 11885 17187 11943 17193
rect 11885 17153 11897 17187
rect 11931 17153 11943 17187
rect 12066 17184 12072 17196
rect 12027 17156 12072 17184
rect 11885 17147 11943 17153
rect 11900 17116 11928 17147
rect 12066 17144 12072 17156
rect 12124 17144 12130 17196
rect 12529 17187 12587 17193
rect 12529 17184 12541 17187
rect 12406 17156 12541 17184
rect 12250 17116 12256 17128
rect 11900 17088 12256 17116
rect 12250 17076 12256 17088
rect 12308 17116 12314 17128
rect 12406 17116 12434 17156
rect 12529 17153 12541 17156
rect 12575 17153 12587 17187
rect 12710 17184 12716 17196
rect 12671 17156 12716 17184
rect 12529 17147 12587 17153
rect 12710 17144 12716 17156
rect 12768 17144 12774 17196
rect 14461 17187 14519 17193
rect 14461 17184 14473 17187
rect 13372 17156 14473 17184
rect 13372 17128 13400 17156
rect 14461 17153 14473 17156
rect 14507 17153 14519 17187
rect 14461 17147 14519 17153
rect 15194 17144 15200 17196
rect 15252 17184 15258 17196
rect 15749 17187 15807 17193
rect 15749 17184 15761 17187
rect 15252 17156 15761 17184
rect 15252 17144 15258 17156
rect 15749 17153 15761 17156
rect 15795 17153 15807 17187
rect 16132 17183 16160 17224
rect 20169 17197 20227 17203
rect 17494 17184 17500 17196
rect 15749 17147 15807 17153
rect 16117 17177 16175 17183
rect 16117 17143 16129 17177
rect 16163 17143 16175 17177
rect 17455 17156 17500 17184
rect 17494 17144 17500 17156
rect 17552 17144 17558 17196
rect 17589 17187 17647 17193
rect 17589 17153 17601 17187
rect 17635 17153 17647 17187
rect 17589 17147 17647 17153
rect 16117 17137 16175 17143
rect 12308 17088 12434 17116
rect 13173 17119 13231 17125
rect 12308 17076 12314 17088
rect 13173 17085 13185 17119
rect 13219 17116 13231 17119
rect 13354 17116 13360 17128
rect 13219 17088 13360 17116
rect 13219 17085 13231 17088
rect 13173 17079 13231 17085
rect 13354 17076 13360 17088
rect 13412 17076 13418 17128
rect 13449 17119 13507 17125
rect 13449 17085 13461 17119
rect 13495 17116 13507 17119
rect 13814 17116 13820 17128
rect 13495 17088 13820 17116
rect 13495 17085 13507 17088
rect 13449 17079 13507 17085
rect 13814 17076 13820 17088
rect 13872 17076 13878 17128
rect 14737 17119 14795 17125
rect 14737 17085 14749 17119
rect 14783 17116 14795 17119
rect 15470 17116 15476 17128
rect 14783 17088 15476 17116
rect 14783 17085 14795 17088
rect 14737 17079 14795 17085
rect 15470 17076 15476 17088
rect 15528 17076 15534 17128
rect 15933 17119 15991 17125
rect 15933 17085 15945 17119
rect 15979 17116 15991 17119
rect 15979 17085 15998 17116
rect 15933 17079 15998 17085
rect 15970 17048 15998 17079
rect 16666 17076 16672 17128
rect 16724 17116 16730 17128
rect 16942 17116 16948 17128
rect 16724 17088 16948 17116
rect 16724 17076 16730 17088
rect 16942 17076 16948 17088
rect 17000 17116 17006 17128
rect 17604 17116 17632 17147
rect 17678 17144 17684 17196
rect 17736 17184 17742 17196
rect 17865 17187 17923 17193
rect 17736 17156 17781 17184
rect 17736 17144 17742 17156
rect 17865 17153 17877 17187
rect 17911 17184 17923 17187
rect 18138 17184 18144 17196
rect 17911 17156 18144 17184
rect 17911 17153 17923 17156
rect 17865 17147 17923 17153
rect 18138 17144 18144 17156
rect 18196 17144 18202 17196
rect 18598 17144 18604 17196
rect 18656 17184 18662 17196
rect 18877 17187 18935 17193
rect 18877 17184 18889 17187
rect 18656 17156 18889 17184
rect 18656 17144 18662 17156
rect 18877 17153 18889 17156
rect 18923 17184 18935 17187
rect 19610 17184 19616 17196
rect 18923 17156 19616 17184
rect 18923 17153 18935 17156
rect 18877 17147 18935 17153
rect 19610 17144 19616 17156
rect 19668 17144 19674 17196
rect 20070 17144 20076 17196
rect 20128 17184 20134 17196
rect 20169 17184 20181 17197
rect 20128 17163 20181 17184
rect 20215 17163 20227 17197
rect 20128 17157 20227 17163
rect 20128 17156 20199 17157
rect 20128 17144 20134 17156
rect 20346 17144 20352 17196
rect 20404 17184 20410 17196
rect 20404 17156 20449 17184
rect 20404 17144 20410 17156
rect 17000 17088 17632 17116
rect 17000 17076 17006 17088
rect 18322 17076 18328 17128
rect 18380 17116 18386 17128
rect 19153 17119 19211 17125
rect 19153 17116 19165 17119
rect 18380 17088 19165 17116
rect 18380 17076 18386 17088
rect 19153 17085 19165 17088
rect 19199 17116 19211 17119
rect 19978 17116 19984 17128
rect 19199 17088 19984 17116
rect 19199 17085 19211 17088
rect 19153 17079 19211 17085
rect 19978 17076 19984 17088
rect 20036 17076 20042 17128
rect 20438 17116 20444 17128
rect 20399 17088 20444 17116
rect 20438 17076 20444 17088
rect 20496 17076 20502 17128
rect 20533 17119 20591 17125
rect 20533 17085 20545 17119
rect 20579 17085 20591 17119
rect 20640 17116 20668 17292
rect 20898 17280 20904 17292
rect 20956 17280 20962 17332
rect 20990 17280 20996 17332
rect 21048 17320 21054 17332
rect 22094 17329 22100 17332
rect 22051 17323 22100 17329
rect 22051 17320 22063 17323
rect 21048 17292 22063 17320
rect 21048 17280 21054 17292
rect 22051 17289 22063 17292
rect 22097 17289 22100 17323
rect 22051 17283 22100 17289
rect 22094 17280 22100 17283
rect 22152 17320 22158 17332
rect 23382 17320 23388 17332
rect 22152 17292 23388 17320
rect 22152 17280 22158 17292
rect 23382 17280 23388 17292
rect 23440 17280 23446 17332
rect 23474 17280 23480 17332
rect 23532 17320 23538 17332
rect 25774 17320 25780 17332
rect 23532 17292 25636 17320
rect 25735 17292 25780 17320
rect 23532 17280 23538 17292
rect 21082 17212 21088 17264
rect 21140 17252 21146 17264
rect 22186 17252 22192 17264
rect 21140 17224 22192 17252
rect 21140 17212 21146 17224
rect 22186 17212 22192 17224
rect 22244 17212 22250 17264
rect 22278 17212 22284 17264
rect 22336 17252 22342 17264
rect 23198 17252 23204 17264
rect 22336 17224 23204 17252
rect 22336 17212 22342 17224
rect 23198 17212 23204 17224
rect 23256 17212 23262 17264
rect 25608 17252 25636 17292
rect 25774 17280 25780 17292
rect 25832 17280 25838 17332
rect 26418 17320 26424 17332
rect 25884 17292 26424 17320
rect 25884 17252 25912 17292
rect 26418 17280 26424 17292
rect 26476 17320 26482 17332
rect 27154 17320 27160 17332
rect 26476 17292 27160 17320
rect 26476 17280 26482 17292
rect 27154 17280 27160 17292
rect 27212 17280 27218 17332
rect 27246 17280 27252 17332
rect 27304 17320 27310 17332
rect 27304 17292 28396 17320
rect 27304 17280 27310 17292
rect 28169 17255 28227 17261
rect 28169 17252 28181 17255
rect 25608 17224 25912 17252
rect 26436 17224 28181 17252
rect 20714 17144 20720 17196
rect 20772 17184 20778 17196
rect 20772 17156 20817 17184
rect 20772 17144 20778 17156
rect 21450 17144 21456 17196
rect 21508 17184 21514 17196
rect 23293 17187 23351 17193
rect 23293 17184 23305 17187
rect 21508 17156 23305 17184
rect 21508 17144 21514 17156
rect 23293 17153 23305 17156
rect 23339 17153 23351 17187
rect 23477 17187 23535 17193
rect 23477 17184 23489 17187
rect 23293 17147 23351 17153
rect 23400 17156 23489 17184
rect 21818 17116 21824 17128
rect 20640 17088 21680 17116
rect 21779 17088 21824 17116
rect 20533 17079 20591 17085
rect 16114 17048 16120 17060
rect 15970 17020 16120 17048
rect 16114 17008 16120 17020
rect 16172 17008 16178 17060
rect 17126 17008 17132 17060
rect 17184 17048 17190 17060
rect 20548 17048 20576 17079
rect 20990 17048 20996 17060
rect 17184 17020 20484 17048
rect 20548 17020 20996 17048
rect 17184 17008 17190 17020
rect 9214 16980 9220 16992
rect 9175 16952 9220 16980
rect 9214 16940 9220 16952
rect 9272 16940 9278 16992
rect 13078 16940 13084 16992
rect 13136 16980 13142 16992
rect 15654 16980 15660 16992
rect 13136 16952 15660 16980
rect 13136 16940 13142 16952
rect 15654 16940 15660 16952
rect 15712 16940 15718 16992
rect 17221 16983 17279 16989
rect 17221 16949 17233 16983
rect 17267 16980 17279 16983
rect 17402 16980 17408 16992
rect 17267 16952 17408 16980
rect 17267 16949 17279 16952
rect 17221 16943 17279 16949
rect 17402 16940 17408 16952
rect 17460 16940 17466 16992
rect 17770 16940 17776 16992
rect 17828 16980 17834 16992
rect 20346 16980 20352 16992
rect 17828 16952 20352 16980
rect 17828 16940 17834 16952
rect 20346 16940 20352 16952
rect 20404 16940 20410 16992
rect 20456 16980 20484 17020
rect 20990 17008 20996 17020
rect 21048 17008 21054 17060
rect 21652 17048 21680 17088
rect 21818 17076 21824 17088
rect 21876 17076 21882 17128
rect 23400 17048 23428 17156
rect 23477 17153 23489 17156
rect 23523 17153 23535 17187
rect 23934 17184 23940 17196
rect 23895 17156 23940 17184
rect 23477 17147 23535 17153
rect 23934 17144 23940 17156
rect 23992 17144 23998 17196
rect 24204 17187 24262 17193
rect 24204 17153 24216 17187
rect 24250 17184 24262 17187
rect 24250 17156 25912 17184
rect 24250 17153 24262 17156
rect 24204 17147 24262 17153
rect 23566 17048 23572 17060
rect 21652 17020 23572 17048
rect 23566 17008 23572 17020
rect 23624 17008 23630 17060
rect 25884 17048 25912 17156
rect 25958 17144 25964 17196
rect 26016 17184 26022 17196
rect 26016 17156 26061 17184
rect 26016 17144 26022 17156
rect 26237 17119 26295 17125
rect 26237 17085 26249 17119
rect 26283 17116 26295 17119
rect 26326 17116 26332 17128
rect 26283 17088 26332 17116
rect 26283 17085 26295 17088
rect 26237 17079 26295 17085
rect 26326 17076 26332 17088
rect 26384 17076 26390 17128
rect 26436 17048 26464 17224
rect 28169 17221 28181 17224
rect 28215 17221 28227 17255
rect 28169 17215 28227 17221
rect 26878 17144 26884 17196
rect 26936 17184 26942 17196
rect 26973 17187 27031 17193
rect 26973 17184 26985 17187
rect 26936 17156 26985 17184
rect 26936 17144 26942 17156
rect 26973 17153 26985 17156
rect 27019 17153 27031 17187
rect 26973 17147 27031 17153
rect 27157 17187 27215 17193
rect 27157 17153 27169 17187
rect 27203 17153 27215 17187
rect 27157 17147 27215 17153
rect 26786 17076 26792 17128
rect 26844 17116 26850 17128
rect 27172 17116 27200 17147
rect 27246 17144 27252 17196
rect 27304 17184 27310 17196
rect 27522 17184 27528 17196
rect 27304 17156 27349 17184
rect 27483 17156 27528 17184
rect 27304 17144 27310 17156
rect 27522 17144 27528 17156
rect 27580 17144 27586 17196
rect 28368 17193 28396 17292
rect 28353 17187 28411 17193
rect 28353 17153 28365 17187
rect 28399 17153 28411 17187
rect 28353 17147 28411 17153
rect 26844 17088 27200 17116
rect 26844 17076 26850 17088
rect 27338 17076 27344 17128
rect 27396 17116 27402 17128
rect 27396 17088 27441 17116
rect 27396 17076 27402 17088
rect 27614 17076 27620 17128
rect 27672 17116 27678 17128
rect 28629 17119 28687 17125
rect 28629 17116 28641 17119
rect 27672 17088 28641 17116
rect 27672 17076 27678 17088
rect 28629 17085 28641 17088
rect 28675 17085 28687 17119
rect 28629 17079 28687 17085
rect 28537 17051 28595 17057
rect 28537 17048 28549 17051
rect 25884 17020 26464 17048
rect 27356 17020 28549 17048
rect 21082 16980 21088 16992
rect 20456 16952 21088 16980
rect 21082 16940 21088 16952
rect 21140 16940 21146 16992
rect 22922 16940 22928 16992
rect 22980 16980 22986 16992
rect 23293 16983 23351 16989
rect 23293 16980 23305 16983
rect 22980 16952 23305 16980
rect 22980 16940 22986 16952
rect 23293 16949 23305 16952
rect 23339 16949 23351 16983
rect 23293 16943 23351 16949
rect 25130 16940 25136 16992
rect 25188 16980 25194 16992
rect 25314 16980 25320 16992
rect 25188 16952 25320 16980
rect 25188 16940 25194 16952
rect 25314 16940 25320 16952
rect 25372 16940 25378 16992
rect 25406 16940 25412 16992
rect 25464 16980 25470 16992
rect 26145 16983 26203 16989
rect 26145 16980 26157 16983
rect 25464 16952 26157 16980
rect 25464 16940 25470 16952
rect 26145 16949 26157 16952
rect 26191 16980 26203 16983
rect 27356 16980 27384 17020
rect 28537 17017 28549 17020
rect 28583 17017 28595 17051
rect 28537 17011 28595 17017
rect 26191 16952 27384 16980
rect 27709 16983 27767 16989
rect 26191 16949 26203 16952
rect 26145 16943 26203 16949
rect 27709 16949 27721 16983
rect 27755 16980 27767 16983
rect 28074 16980 28080 16992
rect 27755 16952 28080 16980
rect 27755 16949 27767 16952
rect 27709 16943 27767 16949
rect 28074 16940 28080 16952
rect 28132 16940 28138 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 11974 16776 11980 16788
rect 11935 16748 11980 16776
rect 11974 16736 11980 16748
rect 12032 16736 12038 16788
rect 15102 16776 15108 16788
rect 15063 16748 15108 16776
rect 15102 16736 15108 16748
rect 15160 16736 15166 16788
rect 15654 16736 15660 16788
rect 15712 16776 15718 16788
rect 19702 16776 19708 16788
rect 15712 16748 19708 16776
rect 15712 16736 15718 16748
rect 19702 16736 19708 16748
rect 19760 16736 19766 16788
rect 19812 16748 21680 16776
rect 7742 16668 7748 16720
rect 7800 16708 7806 16720
rect 9309 16711 9367 16717
rect 9309 16708 9321 16711
rect 7800 16680 9321 16708
rect 7800 16668 7806 16680
rect 9309 16677 9321 16680
rect 9355 16677 9367 16711
rect 15933 16711 15991 16717
rect 9309 16671 9367 16677
rect 13372 16680 15884 16708
rect 8478 16600 8484 16652
rect 8536 16640 8542 16652
rect 10597 16643 10655 16649
rect 10597 16640 10609 16643
rect 8536 16612 10609 16640
rect 8536 16600 8542 16612
rect 10597 16609 10609 16612
rect 10643 16609 10655 16643
rect 10597 16603 10655 16609
rect 8389 16575 8447 16581
rect 8389 16541 8401 16575
rect 8435 16572 8447 16575
rect 9125 16575 9183 16581
rect 8435 16544 9076 16572
rect 8435 16541 8447 16544
rect 8389 16535 8447 16541
rect 8941 16507 8999 16513
rect 8941 16473 8953 16507
rect 8987 16473 8999 16507
rect 9048 16504 9076 16544
rect 9125 16541 9137 16575
rect 9171 16572 9183 16575
rect 9214 16572 9220 16584
rect 9171 16544 9220 16572
rect 9171 16541 9183 16544
rect 9125 16535 9183 16541
rect 9214 16532 9220 16544
rect 9272 16532 9278 16584
rect 10864 16575 10922 16581
rect 10864 16541 10876 16575
rect 10910 16572 10922 16575
rect 11882 16572 11888 16584
rect 10910 16544 11888 16572
rect 10910 16541 10922 16544
rect 10864 16535 10922 16541
rect 11882 16532 11888 16544
rect 11940 16532 11946 16584
rect 12621 16575 12679 16581
rect 12621 16541 12633 16575
rect 12667 16572 12679 16575
rect 12802 16572 12808 16584
rect 12667 16544 12808 16572
rect 12667 16541 12679 16544
rect 12621 16535 12679 16541
rect 12802 16532 12808 16544
rect 12860 16532 12866 16584
rect 13372 16581 13400 16680
rect 15746 16640 15752 16652
rect 14292 16612 15752 16640
rect 13357 16575 13415 16581
rect 13357 16541 13369 16575
rect 13403 16541 13415 16575
rect 13357 16535 13415 16541
rect 13814 16532 13820 16584
rect 13872 16572 13878 16584
rect 14292 16581 14320 16612
rect 15746 16600 15752 16612
rect 15804 16600 15810 16652
rect 15856 16640 15884 16680
rect 15933 16677 15945 16711
rect 15979 16708 15991 16711
rect 16390 16708 16396 16720
rect 15979 16680 16396 16708
rect 15979 16677 15991 16680
rect 15933 16671 15991 16677
rect 16390 16668 16396 16680
rect 16448 16668 16454 16720
rect 16298 16640 16304 16652
rect 15856 16612 16304 16640
rect 16298 16600 16304 16612
rect 16356 16600 16362 16652
rect 16482 16640 16488 16652
rect 16408 16612 16488 16640
rect 14093 16575 14151 16581
rect 14093 16572 14105 16575
rect 13872 16544 14105 16572
rect 13872 16532 13878 16544
rect 14093 16541 14105 16544
rect 14139 16541 14151 16575
rect 14093 16535 14151 16541
rect 14277 16575 14335 16581
rect 14277 16541 14289 16575
rect 14323 16541 14335 16575
rect 14277 16535 14335 16541
rect 14550 16532 14556 16584
rect 14608 16572 14614 16584
rect 14921 16575 14979 16581
rect 14921 16572 14933 16575
rect 14608 16544 14933 16572
rect 14608 16532 14614 16544
rect 14921 16541 14933 16544
rect 14967 16541 14979 16575
rect 14921 16535 14979 16541
rect 15197 16575 15255 16581
rect 15197 16541 15209 16575
rect 15243 16572 15255 16575
rect 16025 16575 16083 16581
rect 15243 16544 15792 16572
rect 15243 16541 15255 16544
rect 15197 16535 15255 16541
rect 10042 16504 10048 16516
rect 9048 16476 10048 16504
rect 8941 16467 8999 16473
rect 8202 16436 8208 16448
rect 8163 16408 8208 16436
rect 8202 16396 8208 16408
rect 8260 16396 8266 16448
rect 8956 16436 8984 16467
rect 10042 16464 10048 16476
rect 10100 16464 10106 16516
rect 13449 16507 13507 16513
rect 13449 16473 13461 16507
rect 13495 16504 13507 16507
rect 14826 16504 14832 16516
rect 13495 16476 14832 16504
rect 13495 16473 13507 16476
rect 13449 16467 13507 16473
rect 14826 16464 14832 16476
rect 14884 16464 14890 16516
rect 14936 16504 14964 16535
rect 15286 16504 15292 16516
rect 14936 16476 15292 16504
rect 15286 16464 15292 16476
rect 15344 16464 15350 16516
rect 15654 16504 15660 16516
rect 15615 16476 15660 16504
rect 15654 16464 15660 16476
rect 15712 16464 15718 16516
rect 15764 16504 15792 16544
rect 16025 16541 16037 16575
rect 16071 16572 16083 16575
rect 16408 16572 16436 16612
rect 16482 16600 16488 16612
rect 16540 16600 16546 16652
rect 17218 16600 17224 16652
rect 17276 16640 17282 16652
rect 19812 16649 19840 16748
rect 17313 16643 17371 16649
rect 17313 16640 17325 16643
rect 17276 16612 17325 16640
rect 17276 16600 17282 16612
rect 17313 16609 17325 16612
rect 17359 16609 17371 16643
rect 17313 16603 17371 16609
rect 19797 16643 19855 16649
rect 19797 16609 19809 16643
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 16758 16572 16764 16584
rect 16071 16544 16436 16572
rect 16500 16544 16764 16572
rect 16071 16541 16083 16544
rect 16025 16535 16083 16541
rect 16500 16516 16528 16544
rect 16758 16532 16764 16544
rect 16816 16532 16822 16584
rect 17402 16532 17408 16584
rect 17460 16572 17466 16584
rect 17569 16575 17627 16581
rect 17569 16572 17581 16575
rect 17460 16544 17581 16572
rect 17460 16532 17466 16544
rect 17569 16541 17581 16544
rect 17615 16541 17627 16575
rect 17569 16535 17627 16541
rect 19334 16532 19340 16584
rect 19392 16572 19398 16584
rect 21652 16581 21680 16748
rect 21818 16736 21824 16788
rect 21876 16776 21882 16788
rect 21876 16748 23520 16776
rect 21876 16736 21882 16748
rect 20053 16575 20111 16581
rect 20053 16572 20065 16575
rect 19392 16544 20065 16572
rect 19392 16532 19398 16544
rect 20053 16541 20065 16544
rect 20099 16541 20111 16575
rect 20053 16535 20111 16541
rect 21637 16575 21695 16581
rect 21637 16541 21649 16575
rect 21683 16572 21695 16575
rect 22462 16572 22468 16584
rect 21683 16544 22468 16572
rect 21683 16541 21695 16544
rect 21637 16535 21695 16541
rect 22462 16532 22468 16544
rect 22520 16532 22526 16584
rect 23492 16581 23520 16748
rect 26786 16736 26792 16788
rect 26844 16736 26850 16788
rect 26881 16779 26939 16785
rect 26881 16745 26893 16779
rect 26927 16776 26939 16779
rect 28350 16776 28356 16788
rect 26927 16748 28356 16776
rect 26927 16745 26939 16748
rect 26881 16739 26939 16745
rect 28350 16736 28356 16748
rect 28408 16736 28414 16788
rect 26804 16708 26832 16736
rect 27062 16708 27068 16720
rect 26344 16680 27068 16708
rect 24854 16640 24860 16652
rect 24815 16612 24860 16640
rect 24854 16600 24860 16612
rect 24912 16600 24918 16652
rect 25774 16600 25780 16652
rect 25832 16640 25838 16652
rect 26344 16640 26372 16680
rect 27062 16668 27068 16680
rect 27120 16668 27126 16720
rect 25832 16612 26372 16640
rect 25832 16600 25838 16612
rect 23477 16575 23535 16581
rect 23477 16541 23489 16575
rect 23523 16541 23535 16575
rect 23477 16535 23535 16541
rect 25133 16575 25191 16581
rect 25133 16541 25145 16575
rect 25179 16541 25191 16575
rect 26142 16572 26148 16584
rect 26103 16544 26148 16572
rect 25133 16535 25191 16541
rect 16114 16504 16120 16516
rect 15764 16476 16120 16504
rect 16114 16464 16120 16476
rect 16172 16464 16178 16516
rect 16482 16464 16488 16516
rect 16540 16464 16546 16516
rect 16666 16504 16672 16516
rect 16627 16476 16672 16504
rect 16666 16464 16672 16476
rect 16724 16464 16730 16516
rect 16850 16464 16856 16516
rect 16908 16504 16914 16516
rect 17310 16504 17316 16516
rect 16908 16476 17316 16504
rect 16908 16464 16914 16476
rect 17310 16464 17316 16476
rect 17368 16464 17374 16516
rect 19794 16504 19800 16516
rect 17512 16476 19800 16504
rect 17512 16448 17540 16476
rect 19794 16464 19800 16476
rect 19852 16464 19858 16516
rect 21904 16507 21962 16513
rect 21904 16473 21916 16507
rect 21950 16504 21962 16507
rect 22186 16504 22192 16516
rect 21950 16476 22192 16504
rect 21950 16473 21962 16476
rect 21904 16467 21962 16473
rect 22186 16464 22192 16476
rect 22244 16464 22250 16516
rect 24578 16504 24584 16516
rect 22296 16476 24584 16504
rect 9674 16436 9680 16448
rect 8956 16408 9680 16436
rect 9674 16396 9680 16408
rect 9732 16396 9738 16448
rect 12434 16396 12440 16448
rect 12492 16436 12498 16448
rect 14277 16439 14335 16445
rect 12492 16408 12537 16436
rect 12492 16396 12498 16408
rect 14277 16405 14289 16439
rect 14323 16436 14335 16439
rect 14458 16436 14464 16448
rect 14323 16408 14464 16436
rect 14323 16405 14335 16408
rect 14277 16399 14335 16405
rect 14458 16396 14464 16408
rect 14516 16396 14522 16448
rect 14737 16439 14795 16445
rect 14737 16405 14749 16439
rect 14783 16436 14795 16439
rect 15102 16436 15108 16448
rect 14783 16408 15108 16436
rect 14783 16405 14795 16408
rect 14737 16399 14795 16405
rect 15102 16396 15108 16408
rect 15160 16396 15166 16448
rect 15749 16439 15807 16445
rect 15749 16405 15761 16439
rect 15795 16436 15807 16439
rect 15838 16436 15844 16448
rect 15795 16408 15844 16436
rect 15795 16405 15807 16408
rect 15749 16399 15807 16405
rect 15838 16396 15844 16408
rect 15896 16396 15902 16448
rect 17494 16396 17500 16448
rect 17552 16396 17558 16448
rect 17586 16396 17592 16448
rect 17644 16436 17650 16448
rect 17954 16436 17960 16448
rect 17644 16408 17960 16436
rect 17644 16396 17650 16408
rect 17954 16396 17960 16408
rect 18012 16436 18018 16448
rect 18693 16439 18751 16445
rect 18693 16436 18705 16439
rect 18012 16408 18705 16436
rect 18012 16396 18018 16408
rect 18693 16405 18705 16408
rect 18739 16405 18751 16439
rect 18693 16399 18751 16405
rect 20346 16396 20352 16448
rect 20404 16436 20410 16448
rect 21177 16439 21235 16445
rect 21177 16436 21189 16439
rect 20404 16408 21189 16436
rect 20404 16396 20410 16408
rect 21177 16405 21189 16408
rect 21223 16436 21235 16439
rect 21542 16436 21548 16448
rect 21223 16408 21548 16436
rect 21223 16405 21235 16408
rect 21177 16399 21235 16405
rect 21542 16396 21548 16408
rect 21600 16396 21606 16448
rect 22094 16396 22100 16448
rect 22152 16436 22158 16448
rect 22296 16436 22324 16476
rect 24578 16464 24584 16476
rect 24636 16464 24642 16516
rect 25148 16504 25176 16535
rect 26142 16532 26148 16544
rect 26200 16532 26206 16584
rect 26344 16581 26372 16612
rect 26421 16643 26479 16649
rect 26421 16609 26433 16643
rect 26467 16640 26479 16643
rect 26786 16640 26792 16652
rect 26467 16612 26792 16640
rect 26467 16609 26479 16612
rect 26421 16603 26479 16609
rect 26786 16600 26792 16612
rect 26844 16600 26850 16652
rect 26970 16600 26976 16652
rect 27028 16640 27034 16652
rect 27617 16643 27675 16649
rect 27617 16640 27629 16643
rect 27028 16612 27629 16640
rect 27028 16600 27034 16612
rect 27617 16609 27629 16612
rect 27663 16609 27675 16643
rect 27617 16603 27675 16609
rect 26329 16575 26387 16581
rect 26329 16541 26341 16575
rect 26375 16541 26387 16575
rect 26329 16535 26387 16541
rect 26513 16575 26571 16581
rect 26513 16541 26525 16575
rect 26559 16541 26571 16575
rect 26513 16535 26571 16541
rect 26697 16575 26755 16581
rect 26697 16541 26709 16575
rect 26743 16572 26755 16575
rect 28718 16572 28724 16584
rect 26743 16544 28724 16572
rect 26743 16541 26755 16544
rect 26697 16535 26755 16541
rect 26234 16504 26240 16516
rect 25148 16476 26240 16504
rect 26234 16464 26240 16476
rect 26292 16504 26298 16516
rect 26528 16504 26556 16535
rect 28718 16532 28724 16544
rect 28776 16532 28782 16584
rect 27338 16504 27344 16516
rect 26292 16476 27344 16504
rect 26292 16464 26298 16476
rect 27338 16464 27344 16476
rect 27396 16464 27402 16516
rect 27884 16507 27942 16513
rect 27884 16473 27896 16507
rect 27930 16504 27942 16507
rect 28166 16504 28172 16516
rect 27930 16476 28172 16504
rect 27930 16473 27942 16476
rect 27884 16467 27942 16473
rect 28166 16464 28172 16476
rect 28224 16464 28230 16516
rect 22152 16408 22324 16436
rect 22152 16396 22158 16408
rect 22646 16396 22652 16448
rect 22704 16436 22710 16448
rect 23014 16436 23020 16448
rect 22704 16408 23020 16436
rect 22704 16396 22710 16408
rect 23014 16396 23020 16408
rect 23072 16396 23078 16448
rect 23569 16439 23627 16445
rect 23569 16405 23581 16439
rect 23615 16436 23627 16439
rect 23750 16436 23756 16448
rect 23615 16408 23756 16436
rect 23615 16405 23627 16408
rect 23569 16399 23627 16405
rect 23750 16396 23756 16408
rect 23808 16396 23814 16448
rect 27798 16396 27804 16448
rect 27856 16436 27862 16448
rect 27982 16436 27988 16448
rect 27856 16408 27988 16436
rect 27856 16396 27862 16408
rect 27982 16396 27988 16408
rect 28040 16436 28046 16448
rect 28626 16436 28632 16448
rect 28040 16408 28632 16436
rect 28040 16396 28046 16408
rect 28626 16396 28632 16408
rect 28684 16436 28690 16448
rect 28997 16439 29055 16445
rect 28997 16436 29009 16439
rect 28684 16408 29009 16436
rect 28684 16396 28690 16408
rect 28997 16405 29009 16408
rect 29043 16405 29055 16439
rect 28997 16399 29055 16405
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 11054 16232 11060 16244
rect 10888 16204 11060 16232
rect 8104 16167 8162 16173
rect 8104 16133 8116 16167
rect 8150 16164 8162 16167
rect 8202 16164 8208 16176
rect 8150 16136 8208 16164
rect 8150 16133 8162 16136
rect 8104 16127 8162 16133
rect 8202 16124 8208 16136
rect 8260 16124 8266 16176
rect 7377 16099 7435 16105
rect 7377 16065 7389 16099
rect 7423 16096 7435 16099
rect 9214 16096 9220 16108
rect 7423 16068 9220 16096
rect 7423 16065 7435 16068
rect 7377 16059 7435 16065
rect 9214 16056 9220 16068
rect 9272 16056 9278 16108
rect 9674 16096 9680 16108
rect 9635 16068 9680 16096
rect 9674 16056 9680 16068
rect 9732 16056 9738 16108
rect 9766 16056 9772 16108
rect 9824 16096 9830 16108
rect 9861 16099 9919 16105
rect 9861 16096 9873 16099
rect 9824 16068 9873 16096
rect 9824 16056 9830 16068
rect 9861 16065 9873 16068
rect 9907 16065 9919 16099
rect 9861 16059 9919 16065
rect 10781 16099 10839 16105
rect 10781 16065 10793 16099
rect 10827 16096 10839 16099
rect 10888 16096 10916 16204
rect 11054 16192 11060 16204
rect 11112 16192 11118 16244
rect 13538 16192 13544 16244
rect 13596 16232 13602 16244
rect 13596 16204 15148 16232
rect 13596 16192 13602 16204
rect 11784 16167 11842 16173
rect 11784 16133 11796 16167
rect 11830 16164 11842 16167
rect 12434 16164 12440 16176
rect 11830 16136 12440 16164
rect 11830 16133 11842 16136
rect 11784 16127 11842 16133
rect 12434 16124 12440 16136
rect 12492 16124 12498 16176
rect 10827 16068 10916 16096
rect 10965 16099 11023 16105
rect 10827 16065 10839 16068
rect 10781 16059 10839 16065
rect 10965 16065 10977 16099
rect 11011 16096 11023 16099
rect 12618 16096 12624 16108
rect 11011 16094 11744 16096
rect 11900 16094 12624 16096
rect 11011 16068 12624 16094
rect 11011 16065 11023 16068
rect 11716 16066 11928 16068
rect 10965 16059 11023 16065
rect 12618 16056 12624 16068
rect 12676 16056 12682 16108
rect 13998 16056 14004 16108
rect 14056 16096 14062 16108
rect 15120 16105 15148 16204
rect 15746 16192 15752 16244
rect 15804 16232 15810 16244
rect 15841 16235 15899 16241
rect 15841 16232 15853 16235
rect 15804 16204 15853 16232
rect 15804 16192 15810 16204
rect 15841 16201 15853 16204
rect 15887 16201 15899 16235
rect 15841 16195 15899 16201
rect 17681 16235 17739 16241
rect 17681 16201 17693 16235
rect 17727 16232 17739 16235
rect 17770 16232 17776 16244
rect 17727 16204 17776 16232
rect 17727 16201 17739 16204
rect 17681 16195 17739 16201
rect 17770 16192 17776 16204
rect 17828 16192 17834 16244
rect 18506 16232 18512 16244
rect 18467 16204 18512 16232
rect 18506 16192 18512 16204
rect 18564 16192 18570 16244
rect 20254 16232 20260 16244
rect 19260 16204 20260 16232
rect 15654 16124 15660 16176
rect 15712 16164 15718 16176
rect 16022 16164 16028 16176
rect 15712 16136 16028 16164
rect 15712 16124 15718 16136
rect 16022 16124 16028 16136
rect 16080 16124 16086 16176
rect 17313 16167 17371 16173
rect 17313 16133 17325 16167
rect 17359 16164 17371 16167
rect 18141 16167 18199 16173
rect 18141 16164 18153 16167
rect 17359 16136 18153 16164
rect 17359 16133 17371 16136
rect 17313 16127 17371 16133
rect 18141 16133 18153 16136
rect 18187 16133 18199 16167
rect 19260 16164 19288 16204
rect 20254 16192 20260 16204
rect 20312 16232 20318 16244
rect 24670 16232 24676 16244
rect 20312 16204 24676 16232
rect 20312 16192 20318 16204
rect 24670 16192 24676 16204
rect 24728 16192 24734 16244
rect 26602 16192 26608 16244
rect 26660 16232 26666 16244
rect 28166 16232 28172 16244
rect 26660 16204 27568 16232
rect 28127 16204 28172 16232
rect 26660 16192 26666 16204
rect 18141 16127 18199 16133
rect 18340 16136 19288 16164
rect 14921 16099 14979 16105
rect 14921 16096 14933 16099
rect 14056 16068 14933 16096
rect 14056 16056 14062 16068
rect 14921 16065 14933 16068
rect 14967 16065 14979 16099
rect 14921 16059 14979 16065
rect 15013 16099 15071 16105
rect 15013 16065 15025 16099
rect 15059 16065 15071 16099
rect 15013 16059 15071 16065
rect 15105 16099 15163 16105
rect 15105 16065 15117 16099
rect 15151 16065 15163 16099
rect 15286 16096 15292 16108
rect 15247 16068 15292 16096
rect 15105 16059 15163 16065
rect 7834 16028 7840 16040
rect 7795 16000 7840 16028
rect 7834 15988 7840 16000
rect 7892 15988 7898 16040
rect 10318 15988 10324 16040
rect 10376 16028 10382 16040
rect 11517 16031 11575 16037
rect 11517 16028 11529 16031
rect 10376 16000 11529 16028
rect 10376 15988 10382 16000
rect 11517 15997 11529 16000
rect 11563 15997 11575 16031
rect 13354 16028 13360 16040
rect 13315 16000 13360 16028
rect 11517 15991 11575 15997
rect 13354 15988 13360 16000
rect 13412 15988 13418 16040
rect 13633 16031 13691 16037
rect 13633 15997 13645 16031
rect 13679 15997 13691 16031
rect 13633 15991 13691 15997
rect 8846 15920 8852 15972
rect 8904 15960 8910 15972
rect 10045 15963 10103 15969
rect 10045 15960 10057 15963
rect 8904 15932 10057 15960
rect 8904 15920 8910 15932
rect 10045 15929 10057 15932
rect 10091 15929 10103 15963
rect 10870 15960 10876 15972
rect 10831 15932 10876 15960
rect 10045 15923 10103 15929
rect 10870 15920 10876 15932
rect 10928 15920 10934 15972
rect 13648 15960 13676 15991
rect 12544 15932 13676 15960
rect 7193 15895 7251 15901
rect 7193 15861 7205 15895
rect 7239 15892 7251 15895
rect 8018 15892 8024 15904
rect 7239 15864 8024 15892
rect 7239 15861 7251 15864
rect 7193 15855 7251 15861
rect 8018 15852 8024 15864
rect 8076 15852 8082 15904
rect 9217 15895 9275 15901
rect 9217 15861 9229 15895
rect 9263 15892 9275 15895
rect 9858 15892 9864 15904
rect 9263 15864 9864 15892
rect 9263 15861 9275 15864
rect 9217 15855 9275 15861
rect 9858 15852 9864 15864
rect 9916 15852 9922 15904
rect 11054 15852 11060 15904
rect 11112 15892 11118 15904
rect 12250 15892 12256 15904
rect 11112 15864 12256 15892
rect 11112 15852 11118 15864
rect 12250 15852 12256 15864
rect 12308 15892 12314 15904
rect 12544 15892 12572 15932
rect 14734 15920 14740 15972
rect 14792 15960 14798 15972
rect 15028 15960 15056 16059
rect 15286 16056 15292 16068
rect 15344 16056 15350 16108
rect 15746 16096 15752 16108
rect 15707 16068 15752 16096
rect 15746 16056 15752 16068
rect 15804 16056 15810 16108
rect 16574 16056 16580 16108
rect 16632 16096 16638 16108
rect 16669 16099 16727 16105
rect 16669 16096 16681 16099
rect 16632 16068 16681 16096
rect 16632 16056 16638 16068
rect 16669 16065 16681 16068
rect 16715 16065 16727 16099
rect 16669 16059 16727 16065
rect 16758 16056 16764 16108
rect 16816 16096 16822 16108
rect 16853 16099 16911 16105
rect 16853 16096 16865 16099
rect 16816 16068 16865 16096
rect 16816 16056 16822 16068
rect 16853 16065 16865 16068
rect 16899 16065 16911 16099
rect 16853 16059 16911 16065
rect 15470 15988 15476 16040
rect 15528 16028 15534 16040
rect 17328 16028 17356 16127
rect 17494 16096 17500 16108
rect 17455 16068 17500 16096
rect 17494 16056 17500 16068
rect 17552 16056 17558 16108
rect 18340 16105 18368 16136
rect 19334 16124 19340 16176
rect 19392 16164 19398 16176
rect 22646 16173 22652 16176
rect 19392 16136 22600 16164
rect 19392 16124 19398 16136
rect 18325 16099 18383 16105
rect 18325 16065 18337 16099
rect 18371 16065 18383 16099
rect 19242 16096 19248 16108
rect 19203 16068 19248 16096
rect 18325 16059 18383 16065
rect 19242 16056 19248 16068
rect 19300 16056 19306 16108
rect 19429 16099 19487 16105
rect 19429 16065 19441 16099
rect 19475 16096 19487 16099
rect 19886 16096 19892 16108
rect 19475 16068 19892 16096
rect 19475 16065 19487 16068
rect 19429 16059 19487 16065
rect 15528 16000 17356 16028
rect 15528 15988 15534 16000
rect 17862 15988 17868 16040
rect 17920 16028 17926 16040
rect 19444 16028 19472 16059
rect 19886 16056 19892 16068
rect 19944 16056 19950 16108
rect 19981 16099 20039 16105
rect 19981 16065 19993 16099
rect 20027 16098 20039 16099
rect 20079 16098 20107 16136
rect 20027 16070 20107 16098
rect 20027 16065 20039 16070
rect 19981 16059 20039 16065
rect 20162 16056 20168 16108
rect 20220 16096 20226 16108
rect 20257 16099 20315 16105
rect 20257 16096 20269 16099
rect 20220 16068 20269 16096
rect 20220 16056 20226 16068
rect 20257 16065 20269 16068
rect 20303 16065 20315 16099
rect 22572 16096 22600 16136
rect 22640 16127 22652 16173
rect 22704 16164 22710 16176
rect 22704 16136 22740 16164
rect 23309 16136 24256 16164
rect 22646 16124 22652 16127
rect 22704 16124 22710 16136
rect 23309 16096 23337 16136
rect 22572 16068 23337 16096
rect 22655 16066 22692 16068
rect 20257 16059 20315 16065
rect 23382 16056 23388 16108
rect 23440 16056 23446 16108
rect 24228 16105 24256 16136
rect 24213 16099 24271 16105
rect 24213 16065 24225 16099
rect 24259 16096 24271 16099
rect 24946 16096 24952 16108
rect 24259 16068 24952 16096
rect 24259 16065 24271 16068
rect 24213 16059 24271 16065
rect 24946 16056 24952 16068
rect 25004 16056 25010 16108
rect 25774 16096 25780 16108
rect 25735 16068 25780 16096
rect 25774 16056 25780 16068
rect 25832 16056 25838 16108
rect 26234 16056 26240 16108
rect 26292 16096 26298 16108
rect 26878 16096 26884 16108
rect 26292 16068 26884 16096
rect 26292 16056 26298 16068
rect 26878 16056 26884 16068
rect 26936 16096 26942 16108
rect 26973 16099 27031 16105
rect 26973 16096 26985 16099
rect 26936 16068 26985 16096
rect 26936 16056 26942 16068
rect 26973 16065 26985 16068
rect 27019 16065 27031 16099
rect 26973 16059 27031 16065
rect 27062 16056 27068 16108
rect 27120 16096 27126 16108
rect 27157 16099 27215 16105
rect 27157 16096 27169 16099
rect 27120 16068 27169 16096
rect 27120 16056 27126 16068
rect 27157 16065 27169 16068
rect 27203 16065 27215 16099
rect 27338 16096 27344 16108
rect 27299 16068 27344 16096
rect 27157 16059 27215 16065
rect 27338 16056 27344 16068
rect 27396 16056 27402 16108
rect 27540 16105 27568 16204
rect 28166 16192 28172 16204
rect 28224 16192 28230 16244
rect 27525 16099 27583 16105
rect 27525 16065 27537 16099
rect 27571 16065 27583 16099
rect 28350 16096 28356 16108
rect 28311 16068 28356 16096
rect 27525 16059 27583 16065
rect 28350 16056 28356 16068
rect 28408 16056 28414 16108
rect 28626 16096 28632 16108
rect 28587 16068 28632 16096
rect 28626 16056 28632 16068
rect 28684 16056 28690 16108
rect 17920 16000 19472 16028
rect 19521 16031 19579 16037
rect 17920 15988 17926 16000
rect 19521 15997 19533 16031
rect 19567 16028 19579 16031
rect 21634 16028 21640 16040
rect 19567 16000 21640 16028
rect 19567 15997 19579 16000
rect 19521 15991 19579 15997
rect 21634 15988 21640 16000
rect 21692 15988 21698 16040
rect 22002 15988 22008 16040
rect 22060 16028 22066 16040
rect 22373 16031 22431 16037
rect 22373 16028 22385 16031
rect 22060 16000 22385 16028
rect 22060 15988 22066 16000
rect 22373 15997 22385 16000
rect 22419 15997 22431 16031
rect 23400 16028 23428 16056
rect 24489 16031 24547 16037
rect 24489 16028 24501 16031
rect 23400 16000 24501 16028
rect 22373 15991 22431 15997
rect 24489 15997 24501 16000
rect 24535 15997 24547 16031
rect 24489 15991 24547 15997
rect 16850 15960 16856 15972
rect 14792 15932 16856 15960
rect 14792 15920 14798 15932
rect 16850 15920 16856 15932
rect 16908 15920 16914 15972
rect 17678 15920 17684 15972
rect 17736 15960 17742 15972
rect 22278 15960 22284 15972
rect 17736 15932 22284 15960
rect 17736 15920 17742 15932
rect 22278 15920 22284 15932
rect 22336 15920 22342 15972
rect 23382 15920 23388 15972
rect 23440 15960 23446 15972
rect 23753 15963 23811 15969
rect 23753 15960 23765 15963
rect 23440 15932 23765 15960
rect 23440 15920 23446 15932
rect 23753 15929 23765 15932
rect 23799 15960 23811 15963
rect 24302 15960 24308 15972
rect 23799 15932 24308 15960
rect 23799 15929 23811 15932
rect 23753 15923 23811 15929
rect 24302 15920 24308 15932
rect 24360 15920 24366 15972
rect 24504 15960 24532 15991
rect 24578 15988 24584 16040
rect 24636 16028 24642 16040
rect 25501 16031 25559 16037
rect 25501 16028 25513 16031
rect 24636 16000 25513 16028
rect 24636 15988 24642 16000
rect 25501 15997 25513 16000
rect 25547 15997 25559 16031
rect 25501 15991 25559 15997
rect 26510 15988 26516 16040
rect 26568 16028 26574 16040
rect 27249 16031 27307 16037
rect 27249 16028 27261 16031
rect 26568 16000 27261 16028
rect 26568 15988 26574 16000
rect 27249 15997 27261 16000
rect 27295 15997 27307 16031
rect 27249 15991 27307 15997
rect 25406 15960 25412 15972
rect 24504 15932 25412 15960
rect 25406 15920 25412 15932
rect 25464 15920 25470 15972
rect 26326 15920 26332 15972
rect 26384 15960 26390 15972
rect 27338 15960 27344 15972
rect 26384 15932 27344 15960
rect 26384 15920 26390 15932
rect 27338 15920 27344 15932
rect 27396 15920 27402 15972
rect 12308 15864 12572 15892
rect 12308 15852 12314 15864
rect 12618 15852 12624 15904
rect 12676 15892 12682 15904
rect 12897 15895 12955 15901
rect 12897 15892 12909 15895
rect 12676 15864 12909 15892
rect 12676 15852 12682 15864
rect 12897 15861 12909 15864
rect 12943 15861 12955 15895
rect 12897 15855 12955 15861
rect 13078 15852 13084 15904
rect 13136 15892 13142 15904
rect 14645 15895 14703 15901
rect 14645 15892 14657 15895
rect 13136 15864 14657 15892
rect 13136 15852 13142 15864
rect 14645 15861 14657 15864
rect 14691 15861 14703 15895
rect 14645 15855 14703 15861
rect 16390 15852 16396 15904
rect 16448 15892 16454 15904
rect 16669 15895 16727 15901
rect 16669 15892 16681 15895
rect 16448 15864 16681 15892
rect 16448 15852 16454 15864
rect 16669 15861 16681 15864
rect 16715 15861 16727 15895
rect 16669 15855 16727 15861
rect 19061 15895 19119 15901
rect 19061 15861 19073 15895
rect 19107 15892 19119 15895
rect 20162 15892 20168 15904
rect 19107 15864 20168 15892
rect 19107 15861 19119 15864
rect 19061 15855 19119 15861
rect 20162 15852 20168 15864
rect 20220 15852 20226 15904
rect 27614 15852 27620 15904
rect 27672 15892 27678 15904
rect 27709 15895 27767 15901
rect 27709 15892 27721 15895
rect 27672 15864 27721 15892
rect 27672 15852 27678 15864
rect 27709 15861 27721 15864
rect 27755 15861 27767 15895
rect 28534 15892 28540 15904
rect 28495 15864 28540 15892
rect 27709 15855 27767 15861
rect 28534 15852 28540 15864
rect 28592 15852 28598 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 8389 15691 8447 15697
rect 8389 15657 8401 15691
rect 8435 15688 8447 15691
rect 9766 15688 9772 15700
rect 8435 15660 9772 15688
rect 8435 15657 8447 15660
rect 8389 15651 8447 15657
rect 9766 15648 9772 15660
rect 9824 15648 9830 15700
rect 12618 15688 12624 15700
rect 12579 15660 12624 15688
rect 12618 15648 12624 15660
rect 12676 15648 12682 15700
rect 12802 15688 12808 15700
rect 12763 15660 12808 15688
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 15654 15688 15660 15700
rect 14673 15660 15660 15688
rect 10318 15552 10324 15564
rect 10279 15524 10324 15552
rect 10318 15512 10324 15524
rect 10376 15512 10382 15564
rect 14673 15552 14701 15660
rect 15654 15648 15660 15660
rect 15712 15648 15718 15700
rect 17494 15648 17500 15700
rect 17552 15688 17558 15700
rect 17678 15688 17684 15700
rect 17552 15660 17597 15688
rect 17639 15660 17684 15688
rect 17552 15648 17558 15660
rect 17678 15648 17684 15660
rect 17736 15648 17742 15700
rect 18325 15691 18383 15697
rect 18325 15657 18337 15691
rect 18371 15688 18383 15691
rect 18690 15688 18696 15700
rect 18371 15660 18696 15688
rect 18371 15657 18383 15660
rect 18325 15651 18383 15657
rect 18690 15648 18696 15660
rect 18748 15648 18754 15700
rect 20438 15648 20444 15700
rect 20496 15688 20502 15700
rect 21913 15691 21971 15697
rect 21913 15688 21925 15691
rect 20496 15660 21925 15688
rect 20496 15648 20502 15660
rect 21913 15657 21925 15660
rect 21959 15657 21971 15691
rect 21913 15651 21971 15657
rect 22557 15691 22615 15697
rect 22557 15657 22569 15691
rect 22603 15688 22615 15691
rect 22646 15688 22652 15700
rect 22603 15660 22652 15688
rect 22603 15657 22615 15660
rect 22557 15651 22615 15657
rect 22646 15648 22652 15660
rect 22704 15648 22710 15700
rect 22925 15691 22983 15697
rect 22925 15657 22937 15691
rect 22971 15688 22983 15691
rect 23290 15688 23296 15700
rect 22971 15660 23296 15688
rect 22971 15657 22983 15660
rect 22925 15651 22983 15657
rect 23290 15648 23296 15660
rect 23348 15648 23354 15700
rect 23566 15688 23572 15700
rect 23527 15660 23572 15688
rect 23566 15648 23572 15660
rect 23624 15648 23630 15700
rect 16853 15623 16911 15629
rect 16853 15589 16865 15623
rect 16899 15589 16911 15623
rect 16853 15583 16911 15589
rect 14660 15524 14701 15552
rect 16868 15552 16896 15583
rect 16942 15580 16948 15632
rect 17000 15620 17006 15632
rect 19613 15623 19671 15629
rect 19613 15620 19625 15623
rect 17000 15592 19625 15620
rect 17000 15580 17006 15592
rect 19613 15589 19625 15592
rect 19659 15589 19671 15623
rect 19613 15583 19671 15589
rect 21453 15623 21511 15629
rect 21453 15589 21465 15623
rect 21499 15620 21511 15623
rect 21634 15620 21640 15632
rect 21499 15592 21640 15620
rect 21499 15589 21511 15592
rect 21453 15583 21511 15589
rect 17310 15552 17316 15564
rect 16868 15524 17316 15552
rect 7009 15487 7067 15493
rect 7009 15453 7021 15487
rect 7055 15484 7067 15487
rect 7834 15484 7840 15496
rect 7055 15456 7840 15484
rect 7055 15453 7067 15456
rect 7009 15447 7067 15453
rect 7834 15444 7840 15456
rect 7892 15444 7898 15496
rect 8941 15487 8999 15493
rect 8941 15453 8953 15487
rect 8987 15484 8999 15487
rect 9674 15484 9680 15496
rect 8987 15456 9680 15484
rect 8987 15453 8999 15456
rect 8941 15447 8999 15453
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 12526 15444 12532 15496
rect 12584 15484 12590 15496
rect 13354 15484 13360 15496
rect 12584 15456 13360 15484
rect 12584 15444 12590 15456
rect 13354 15444 13360 15456
rect 13412 15484 13418 15496
rect 14660 15493 14688 15524
rect 17310 15512 17316 15524
rect 17368 15552 17374 15564
rect 19518 15552 19524 15564
rect 17368 15524 19524 15552
rect 17368 15512 17374 15524
rect 19518 15512 19524 15524
rect 19576 15512 19582 15564
rect 13449 15487 13507 15493
rect 13449 15484 13461 15487
rect 13412 15456 13461 15484
rect 13412 15444 13418 15456
rect 13449 15453 13461 15456
rect 13495 15453 13507 15487
rect 13449 15447 13507 15453
rect 14625 15487 14688 15493
rect 14625 15453 14637 15487
rect 14671 15456 14688 15487
rect 14718 15484 14776 15490
rect 14671 15453 14683 15456
rect 14625 15447 14683 15453
rect 14718 15450 14730 15484
rect 14764 15481 14776 15484
rect 14764 15480 14777 15481
rect 14764 15450 14780 15480
rect 14718 15444 14780 15450
rect 14826 15444 14832 15496
rect 14884 15484 14890 15496
rect 15013 15487 15071 15493
rect 14884 15456 14929 15484
rect 14884 15444 14890 15456
rect 15013 15453 15025 15487
rect 15059 15484 15071 15487
rect 15286 15484 15292 15496
rect 15059 15456 15292 15484
rect 15059 15453 15071 15456
rect 15013 15447 15071 15453
rect 15286 15444 15292 15456
rect 15344 15444 15350 15496
rect 15470 15484 15476 15496
rect 15431 15456 15476 15484
rect 15470 15444 15476 15456
rect 15528 15484 15534 15496
rect 17218 15484 17224 15496
rect 15528 15456 17224 15484
rect 15528 15444 15534 15456
rect 17218 15444 17224 15456
rect 17276 15444 17282 15496
rect 19058 15484 19064 15496
rect 18616 15456 19064 15484
rect 7282 15425 7288 15428
rect 7276 15379 7288 15425
rect 7340 15416 7346 15428
rect 9122 15416 9128 15428
rect 7340 15388 7376 15416
rect 9083 15388 9128 15416
rect 7282 15376 7288 15379
rect 7340 15376 7346 15388
rect 9122 15376 9128 15388
rect 9180 15376 9186 15428
rect 10588 15419 10646 15425
rect 10588 15385 10600 15419
rect 10634 15416 10646 15419
rect 10778 15416 10784 15428
rect 10634 15388 10784 15416
rect 10634 15385 10646 15388
rect 10588 15379 10646 15385
rect 10778 15376 10784 15388
rect 10836 15376 10842 15428
rect 12434 15416 12440 15428
rect 12395 15388 12440 15416
rect 12434 15376 12440 15388
rect 12492 15376 12498 15428
rect 14752 15360 14780 15444
rect 15102 15376 15108 15428
rect 15160 15416 15166 15428
rect 15718 15419 15776 15425
rect 15718 15416 15730 15419
rect 15160 15388 15730 15416
rect 15160 15376 15166 15388
rect 15718 15385 15730 15388
rect 15764 15385 15776 15419
rect 15718 15379 15776 15385
rect 16022 15376 16028 15428
rect 16080 15416 16086 15428
rect 17313 15419 17371 15425
rect 17313 15416 17325 15419
rect 16080 15388 17325 15416
rect 16080 15376 16086 15388
rect 17313 15385 17325 15388
rect 17359 15385 17371 15419
rect 18233 15419 18291 15425
rect 17313 15379 17371 15385
rect 17420 15388 18000 15416
rect 9306 15348 9312 15360
rect 9267 15320 9312 15348
rect 9306 15308 9312 15320
rect 9364 15308 9370 15360
rect 11698 15348 11704 15360
rect 11659 15320 11704 15348
rect 11698 15308 11704 15320
rect 11756 15308 11762 15360
rect 12250 15308 12256 15360
rect 12308 15348 12314 15360
rect 12637 15351 12695 15357
rect 12637 15348 12649 15351
rect 12308 15320 12649 15348
rect 12308 15308 12314 15320
rect 12637 15317 12649 15320
rect 12683 15317 12695 15351
rect 13262 15348 13268 15360
rect 13223 15320 13268 15348
rect 12637 15311 12695 15317
rect 13262 15308 13268 15320
rect 13320 15308 13326 15360
rect 14274 15308 14280 15360
rect 14332 15348 14338 15360
rect 14369 15351 14427 15357
rect 14369 15348 14381 15351
rect 14332 15320 14381 15348
rect 14332 15308 14338 15320
rect 14369 15317 14381 15320
rect 14415 15317 14427 15351
rect 14369 15311 14427 15317
rect 14734 15308 14740 15360
rect 14792 15308 14798 15360
rect 16574 15308 16580 15360
rect 16632 15348 16638 15360
rect 17420 15348 17448 15388
rect 16632 15320 17448 15348
rect 17523 15351 17581 15357
rect 16632 15308 16638 15320
rect 17523 15317 17535 15351
rect 17569 15348 17581 15351
rect 17678 15348 17684 15360
rect 17569 15320 17684 15348
rect 17569 15317 17581 15320
rect 17523 15311 17581 15317
rect 17678 15308 17684 15320
rect 17736 15308 17742 15360
rect 17972 15348 18000 15388
rect 18233 15385 18245 15419
rect 18279 15416 18291 15419
rect 18616 15416 18644 15456
rect 19058 15444 19064 15456
rect 19116 15444 19122 15496
rect 18279 15388 18644 15416
rect 18279 15385 18291 15388
rect 18233 15379 18291 15385
rect 18690 15376 18696 15428
rect 18748 15416 18754 15428
rect 19429 15419 19487 15425
rect 19429 15416 19441 15419
rect 18748 15388 19441 15416
rect 18748 15376 18754 15388
rect 19429 15385 19441 15388
rect 19475 15385 19487 15419
rect 19429 15379 19487 15385
rect 19518 15376 19524 15428
rect 19576 15376 19582 15428
rect 19536 15348 19564 15376
rect 17972 15320 19564 15348
rect 19628 15348 19656 15583
rect 21634 15580 21640 15592
rect 21692 15580 21698 15632
rect 22094 15620 22100 15632
rect 22066 15580 22100 15620
rect 22152 15580 22158 15632
rect 22278 15580 22284 15632
rect 22336 15620 22342 15632
rect 25590 15620 25596 15632
rect 22336 15592 25596 15620
rect 22336 15580 22342 15592
rect 25590 15580 25596 15592
rect 25648 15580 25654 15632
rect 27801 15623 27859 15629
rect 27801 15620 27813 15623
rect 26436 15592 27813 15620
rect 21082 15512 21088 15564
rect 21140 15552 21146 15564
rect 21542 15552 21548 15564
rect 21140 15524 21548 15552
rect 21140 15512 21146 15524
rect 21542 15512 21548 15524
rect 21600 15552 21606 15564
rect 22066 15552 22094 15580
rect 21600 15524 22094 15552
rect 21600 15512 21606 15524
rect 22462 15512 22468 15564
rect 22520 15552 22526 15564
rect 23017 15555 23075 15561
rect 23017 15552 23029 15555
rect 22520 15524 23029 15552
rect 22520 15512 22526 15524
rect 23017 15521 23029 15524
rect 23063 15552 23075 15555
rect 23382 15552 23388 15564
rect 23063 15524 23388 15552
rect 23063 15521 23075 15524
rect 23017 15515 23075 15521
rect 23382 15512 23388 15524
rect 23440 15512 23446 15564
rect 24765 15555 24823 15561
rect 23584 15524 24532 15552
rect 20073 15487 20131 15493
rect 20073 15453 20085 15487
rect 20119 15484 20131 15487
rect 21910 15484 21916 15496
rect 20119 15456 21916 15484
rect 20119 15453 20131 15456
rect 20073 15447 20131 15453
rect 21910 15444 21916 15456
rect 21968 15444 21974 15496
rect 22097 15487 22155 15493
rect 22097 15453 22109 15487
rect 22143 15453 22155 15487
rect 22738 15484 22744 15496
rect 22699 15456 22744 15484
rect 22097 15447 22155 15453
rect 20162 15376 20168 15428
rect 20220 15416 20226 15428
rect 20318 15419 20376 15425
rect 20318 15416 20330 15419
rect 20220 15388 20330 15416
rect 20220 15376 20226 15388
rect 20318 15385 20330 15388
rect 20364 15385 20376 15419
rect 20318 15379 20376 15385
rect 21542 15376 21548 15428
rect 21600 15416 21606 15428
rect 22112 15416 22140 15447
rect 22738 15444 22744 15456
rect 22796 15444 22802 15496
rect 23474 15484 23480 15496
rect 23435 15456 23480 15484
rect 23474 15444 23480 15456
rect 23532 15444 23538 15496
rect 21600 15388 22140 15416
rect 21600 15376 21606 15388
rect 22554 15376 22560 15428
rect 22612 15416 22618 15428
rect 23584 15416 23612 15524
rect 24397 15487 24455 15493
rect 24397 15453 24409 15487
rect 24443 15453 24455 15487
rect 24504 15484 24532 15524
rect 24765 15521 24777 15555
rect 24811 15552 24823 15555
rect 24854 15552 24860 15564
rect 24811 15524 24860 15552
rect 24811 15521 24823 15524
rect 24765 15515 24823 15521
rect 24854 15512 24860 15524
rect 24912 15512 24918 15564
rect 25038 15512 25044 15564
rect 25096 15552 25102 15564
rect 26436 15561 26464 15592
rect 27801 15589 27813 15592
rect 27847 15620 27859 15623
rect 28534 15620 28540 15632
rect 27847 15592 28540 15620
rect 27847 15589 27859 15592
rect 27801 15583 27859 15589
rect 28534 15580 28540 15592
rect 28592 15620 28598 15632
rect 28721 15623 28779 15629
rect 28721 15620 28733 15623
rect 28592 15592 28733 15620
rect 28592 15580 28598 15592
rect 28721 15589 28733 15592
rect 28767 15589 28779 15623
rect 28721 15583 28779 15589
rect 26145 15555 26203 15561
rect 26145 15552 26157 15555
rect 25096 15524 26157 15552
rect 25096 15512 25102 15524
rect 26145 15521 26157 15524
rect 26191 15521 26203 15555
rect 26145 15515 26203 15521
rect 26421 15555 26479 15561
rect 26421 15521 26433 15555
rect 26467 15521 26479 15555
rect 27890 15552 27896 15564
rect 27851 15524 27896 15552
rect 26421 15515 26479 15521
rect 27890 15512 27896 15524
rect 27948 15512 27954 15564
rect 28442 15512 28448 15564
rect 28500 15552 28506 15564
rect 28813 15555 28871 15561
rect 28813 15552 28825 15555
rect 28500 15524 28825 15552
rect 28500 15512 28506 15524
rect 28813 15521 28825 15524
rect 28859 15521 28871 15555
rect 28813 15515 28871 15521
rect 24578 15493 24584 15496
rect 24569 15487 24584 15493
rect 24569 15484 24581 15487
rect 24491 15456 24581 15484
rect 24397 15447 24455 15453
rect 24569 15453 24581 15456
rect 24569 15447 24584 15453
rect 22612 15388 23612 15416
rect 24412 15416 24440 15447
rect 24578 15444 24584 15447
rect 24636 15444 24642 15496
rect 24670 15444 24676 15496
rect 24728 15484 24734 15496
rect 24949 15487 25007 15493
rect 24728 15456 24773 15484
rect 24728 15444 24734 15456
rect 24949 15453 24961 15487
rect 24995 15484 25007 15487
rect 25222 15484 25228 15496
rect 24995 15456 25228 15484
rect 24995 15453 25007 15456
rect 24949 15447 25007 15453
rect 25222 15444 25228 15456
rect 25280 15444 25286 15496
rect 27614 15484 27620 15496
rect 27575 15456 27620 15484
rect 27614 15444 27620 15456
rect 27672 15444 27678 15496
rect 28074 15444 28080 15496
rect 28132 15484 28138 15496
rect 28537 15487 28595 15493
rect 28537 15484 28549 15487
rect 28132 15456 28549 15484
rect 28132 15444 28138 15456
rect 28537 15453 28549 15456
rect 28583 15453 28595 15487
rect 28537 15447 28595 15453
rect 26234 15416 26240 15428
rect 24412 15388 26240 15416
rect 22612 15376 22618 15388
rect 24412 15348 24440 15388
rect 26234 15376 26240 15388
rect 26292 15376 26298 15428
rect 19628 15320 24440 15348
rect 25038 15308 25044 15360
rect 25096 15348 25102 15360
rect 25133 15351 25191 15357
rect 25133 15348 25145 15351
rect 25096 15320 25145 15348
rect 25096 15308 25102 15320
rect 25133 15317 25145 15320
rect 25179 15317 25191 15351
rect 27430 15348 27436 15360
rect 27391 15320 27436 15348
rect 25133 15311 25191 15317
rect 27430 15308 27436 15320
rect 27488 15308 27494 15360
rect 28350 15348 28356 15360
rect 28311 15320 28356 15348
rect 28350 15308 28356 15320
rect 28408 15308 28414 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 7193 15147 7251 15153
rect 7193 15113 7205 15147
rect 7239 15144 7251 15147
rect 7282 15144 7288 15156
rect 7239 15116 7288 15144
rect 7239 15113 7251 15116
rect 7193 15107 7251 15113
rect 7282 15104 7288 15116
rect 7340 15104 7346 15156
rect 9122 15104 9128 15156
rect 9180 15144 9186 15156
rect 9217 15147 9275 15153
rect 9217 15144 9229 15147
rect 9180 15116 9229 15144
rect 9180 15104 9186 15116
rect 9217 15113 9229 15116
rect 9263 15113 9275 15147
rect 10042 15144 10048 15156
rect 10003 15116 10048 15144
rect 9217 15107 9275 15113
rect 10042 15104 10048 15116
rect 10100 15104 10106 15156
rect 10778 15144 10784 15156
rect 10739 15116 10784 15144
rect 10778 15104 10784 15116
rect 10836 15104 10842 15156
rect 11727 15147 11785 15153
rect 11727 15113 11739 15147
rect 11773 15144 11785 15147
rect 12250 15144 12256 15156
rect 11773 15116 12256 15144
rect 11773 15113 11785 15116
rect 11727 15107 11785 15113
rect 12250 15104 12256 15116
rect 12308 15104 12314 15156
rect 12342 15104 12348 15156
rect 12400 15144 12406 15156
rect 17402 15144 17408 15156
rect 12400 15116 17408 15144
rect 12400 15104 12406 15116
rect 17402 15104 17408 15116
rect 17460 15104 17466 15156
rect 18414 15104 18420 15156
rect 18472 15104 18478 15156
rect 20530 15144 20536 15156
rect 18708 15116 20536 15144
rect 8846 15076 8852 15088
rect 7392 15048 8852 15076
rect 7392 15017 7420 15048
rect 8846 15036 8852 15048
rect 8904 15036 8910 15088
rect 9858 15076 9864 15088
rect 9819 15048 9864 15076
rect 9858 15036 9864 15048
rect 9916 15036 9922 15088
rect 11514 15076 11520 15088
rect 11475 15048 11520 15076
rect 11514 15036 11520 15048
rect 11572 15036 11578 15088
rect 12980 15079 13038 15085
rect 12980 15045 12992 15079
rect 13026 15076 13038 15079
rect 13078 15076 13084 15088
rect 13026 15048 13084 15076
rect 13026 15045 13038 15048
rect 12980 15039 13038 15045
rect 13078 15036 13084 15048
rect 13136 15036 13142 15088
rect 15470 15076 15476 15088
rect 14568 15048 15476 15076
rect 8110 15017 8116 15020
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 14977 7435 15011
rect 7377 14971 7435 14977
rect 8104 14971 8116 15017
rect 8168 15008 8174 15020
rect 9674 15008 9680 15020
rect 8168 14980 8204 15008
rect 9587 14980 9680 15008
rect 8110 14968 8116 14971
rect 8168 14968 8174 14980
rect 9674 14968 9680 14980
rect 9732 15008 9738 15020
rect 10502 15008 10508 15020
rect 9732 14980 10508 15008
rect 9732 14968 9738 14980
rect 10502 14968 10508 14980
rect 10560 14968 10566 15020
rect 14568 15017 14596 15048
rect 15470 15036 15476 15048
rect 15528 15036 15534 15088
rect 17497 15079 17555 15085
rect 17497 15076 17509 15079
rect 15580 15048 17509 15076
rect 10965 15011 11023 15017
rect 10965 14977 10977 15011
rect 11011 15008 11023 15011
rect 14553 15011 14611 15017
rect 11011 14980 11928 15008
rect 11011 14977 11023 14980
rect 10965 14971 11023 14977
rect 7834 14940 7840 14952
rect 7795 14912 7840 14940
rect 7834 14900 7840 14912
rect 7892 14900 7898 14952
rect 11900 14881 11928 14980
rect 14553 14977 14565 15011
rect 14599 14977 14611 15011
rect 14809 15011 14867 15017
rect 14809 15008 14821 15011
rect 14553 14971 14611 14977
rect 14660 14980 14821 15008
rect 12710 14940 12716 14952
rect 12671 14912 12716 14940
rect 12710 14900 12716 14912
rect 12768 14900 12774 14952
rect 14274 14900 14280 14952
rect 14332 14940 14338 14952
rect 14660 14940 14688 14980
rect 14809 14977 14821 14980
rect 14855 14977 14867 15011
rect 14809 14971 14867 14977
rect 14332 14912 14688 14940
rect 14332 14900 14338 14912
rect 11885 14875 11943 14881
rect 11885 14841 11897 14875
rect 11931 14841 11943 14875
rect 11885 14835 11943 14841
rect 13998 14832 14004 14884
rect 14056 14872 14062 14884
rect 14093 14875 14151 14881
rect 14093 14872 14105 14875
rect 14056 14844 14105 14872
rect 14056 14832 14062 14844
rect 14093 14841 14105 14844
rect 14139 14841 14151 14875
rect 14093 14835 14151 14841
rect 11698 14804 11704 14816
rect 11659 14776 11704 14804
rect 11698 14764 11704 14776
rect 11756 14764 11762 14816
rect 14108 14804 14136 14835
rect 15580 14804 15608 15048
rect 17497 15045 17509 15048
rect 17543 15045 17555 15079
rect 17497 15039 17555 15045
rect 17129 15011 17187 15017
rect 17129 14977 17141 15011
rect 17175 14977 17187 15011
rect 17129 14971 17187 14977
rect 15933 14875 15991 14881
rect 15933 14841 15945 14875
rect 15979 14872 15991 14875
rect 16022 14872 16028 14884
rect 15979 14844 16028 14872
rect 15979 14841 15991 14844
rect 15933 14835 15991 14841
rect 16022 14832 16028 14844
rect 16080 14832 16086 14884
rect 14108 14776 15608 14804
rect 16574 14764 16580 14816
rect 16632 14804 16638 14816
rect 17144 14804 17172 14971
rect 17218 14968 17224 15020
rect 17276 15008 17282 15020
rect 17678 15017 17684 15020
rect 17405 15011 17463 15017
rect 17276 14980 17321 15008
rect 17276 14968 17282 14980
rect 17405 14977 17417 15011
rect 17451 14977 17463 15011
rect 17405 14971 17463 14977
rect 17635 15011 17684 15017
rect 17635 14977 17647 15011
rect 17681 14977 17684 15011
rect 17635 14971 17684 14977
rect 17218 14832 17224 14884
rect 17276 14872 17282 14884
rect 17420 14872 17448 14971
rect 17678 14968 17684 14971
rect 17736 15008 17742 15020
rect 18138 15008 18144 15020
rect 17736 14980 18144 15008
rect 17736 14968 17742 14980
rect 18138 14968 18144 14980
rect 18196 14968 18202 15020
rect 18230 14968 18236 15020
rect 18288 15008 18294 15020
rect 18433 15017 18461 15104
rect 18325 15011 18383 15017
rect 18325 15008 18337 15011
rect 18288 14980 18337 15008
rect 18288 14968 18294 14980
rect 18325 14977 18337 14980
rect 18371 14977 18383 15011
rect 18325 14971 18383 14977
rect 18418 15011 18476 15017
rect 18418 14977 18430 15011
rect 18464 14977 18476 15011
rect 18598 15008 18604 15020
rect 18559 14980 18604 15008
rect 18418 14971 18476 14977
rect 18598 14968 18604 14980
rect 18656 14968 18662 15020
rect 18708 15017 18736 15116
rect 20530 15104 20536 15116
rect 20588 15104 20594 15156
rect 22186 15144 22192 15156
rect 22147 15116 22192 15144
rect 22186 15104 22192 15116
rect 22244 15104 22250 15156
rect 25961 15147 26019 15153
rect 25961 15113 25973 15147
rect 26007 15144 26019 15147
rect 26050 15144 26056 15156
rect 26007 15116 26056 15144
rect 26007 15113 26019 15116
rect 25961 15107 26019 15113
rect 26050 15104 26056 15116
rect 26108 15104 26114 15156
rect 27890 15104 27896 15156
rect 27948 15144 27954 15156
rect 28353 15147 28411 15153
rect 28353 15144 28365 15147
rect 27948 15116 28365 15144
rect 27948 15104 27954 15116
rect 28353 15113 28365 15116
rect 28399 15113 28411 15147
rect 28353 15107 28411 15113
rect 21358 15076 21364 15088
rect 19536 15048 21364 15076
rect 19536 15017 19564 15048
rect 21358 15036 21364 15048
rect 21416 15036 21422 15088
rect 27240 15079 27298 15085
rect 27240 15045 27252 15079
rect 27286 15076 27298 15079
rect 27430 15076 27436 15088
rect 27286 15048 27436 15076
rect 27286 15045 27298 15048
rect 27240 15039 27298 15045
rect 27430 15036 27436 15048
rect 27488 15036 27494 15088
rect 18693 15011 18751 15017
rect 18693 14977 18705 15011
rect 18739 14977 18751 15011
rect 18693 14971 18751 14977
rect 18790 15011 18848 15017
rect 18790 14977 18802 15011
rect 18836 14977 18848 15011
rect 18790 14971 18848 14977
rect 19521 15011 19579 15017
rect 19521 14977 19533 15011
rect 19567 14977 19579 15011
rect 19521 14971 19579 14977
rect 19628 14980 20300 15008
rect 18248 14940 18276 14968
rect 17276 14844 17448 14872
rect 17512 14912 18276 14940
rect 17276 14832 17282 14844
rect 17512 14804 17540 14912
rect 17862 14832 17868 14884
rect 17920 14872 17926 14884
rect 18805 14872 18833 14971
rect 19242 14900 19248 14952
rect 19300 14940 19306 14952
rect 19628 14940 19656 14980
rect 19300 14912 19656 14940
rect 19797 14943 19855 14949
rect 19300 14900 19306 14912
rect 19797 14909 19809 14943
rect 19843 14940 19855 14943
rect 20162 14940 20168 14952
rect 19843 14912 20168 14940
rect 19843 14909 19855 14912
rect 19797 14903 19855 14909
rect 20162 14900 20168 14912
rect 20220 14900 20226 14952
rect 20272 14940 20300 14980
rect 20714 14968 20720 15020
rect 20772 15008 20778 15020
rect 20993 15011 21051 15017
rect 20993 15008 21005 15011
rect 20772 14980 21005 15008
rect 20772 14968 20778 14980
rect 20993 14977 21005 14980
rect 21039 14977 21051 15011
rect 22370 15008 22376 15020
rect 22331 14980 22376 15008
rect 20993 14971 21051 14977
rect 22370 14968 22376 14980
rect 22428 14968 22434 15020
rect 22649 15011 22707 15017
rect 22649 14977 22661 15011
rect 22695 15008 22707 15011
rect 23014 15008 23020 15020
rect 22695 14980 23020 15008
rect 22695 14977 22707 14980
rect 22649 14971 22707 14977
rect 23014 14968 23020 14980
rect 23072 14968 23078 15020
rect 23477 15011 23535 15017
rect 23477 14977 23489 15011
rect 23523 15008 23535 15011
rect 23566 15008 23572 15020
rect 23523 14980 23572 15008
rect 23523 14977 23535 14980
rect 23477 14971 23535 14977
rect 23566 14968 23572 14980
rect 23624 14968 23630 15020
rect 24118 15008 24124 15020
rect 24079 14980 24124 15008
rect 24118 14968 24124 14980
rect 24176 14968 24182 15020
rect 24854 15017 24860 15020
rect 24848 14971 24860 15017
rect 24912 15008 24918 15020
rect 26970 15008 26976 15020
rect 24912 14980 24948 15008
rect 26931 14980 26976 15008
rect 24854 14968 24860 14971
rect 24912 14968 24918 14980
rect 26970 14968 26976 14980
rect 27028 14968 27034 15020
rect 21818 14940 21824 14952
rect 20272 14912 21824 14940
rect 21818 14900 21824 14912
rect 21876 14900 21882 14952
rect 22557 14943 22615 14949
rect 22557 14909 22569 14943
rect 22603 14940 22615 14943
rect 23290 14940 23296 14952
rect 22603 14912 23296 14940
rect 22603 14909 22615 14912
rect 22557 14903 22615 14909
rect 23290 14900 23296 14912
rect 23348 14900 23354 14952
rect 24578 14940 24584 14952
rect 24539 14912 24584 14940
rect 24578 14900 24584 14912
rect 24636 14900 24642 14952
rect 18874 14872 18880 14884
rect 17920 14844 18880 14872
rect 17920 14832 17926 14844
rect 18874 14832 18880 14844
rect 18932 14832 18938 14884
rect 18969 14875 19027 14881
rect 18969 14841 18981 14875
rect 19015 14872 19027 14875
rect 22094 14872 22100 14884
rect 19015 14844 22100 14872
rect 19015 14841 19027 14844
rect 18969 14835 19027 14841
rect 22094 14832 22100 14844
rect 22152 14832 22158 14884
rect 16632 14776 17540 14804
rect 17773 14807 17831 14813
rect 16632 14764 16638 14776
rect 17773 14773 17785 14807
rect 17819 14804 17831 14807
rect 19242 14804 19248 14816
rect 17819 14776 19248 14804
rect 17819 14773 17831 14776
rect 17773 14767 17831 14773
rect 19242 14764 19248 14776
rect 19300 14764 19306 14816
rect 20806 14804 20812 14816
rect 20767 14776 20812 14804
rect 20806 14764 20812 14776
rect 20864 14764 20870 14816
rect 23290 14804 23296 14816
rect 23251 14776 23296 14804
rect 23290 14764 23296 14776
rect 23348 14764 23354 14816
rect 23934 14804 23940 14816
rect 23895 14776 23940 14804
rect 23934 14764 23940 14776
rect 23992 14764 23998 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 7561 14603 7619 14609
rect 7561 14569 7573 14603
rect 7607 14600 7619 14603
rect 7926 14600 7932 14612
rect 7607 14572 7932 14600
rect 7607 14569 7619 14572
rect 7561 14563 7619 14569
rect 7926 14560 7932 14572
rect 7984 14560 7990 14612
rect 8110 14560 8116 14612
rect 8168 14600 8174 14612
rect 8205 14603 8263 14609
rect 8205 14600 8217 14603
rect 8168 14572 8217 14600
rect 8168 14560 8174 14572
rect 8205 14569 8217 14572
rect 8251 14569 8263 14603
rect 8205 14563 8263 14569
rect 9214 14560 9220 14612
rect 9272 14600 9278 14612
rect 9309 14603 9367 14609
rect 9309 14600 9321 14603
rect 9272 14572 9321 14600
rect 9272 14560 9278 14572
rect 9309 14569 9321 14572
rect 9355 14569 9367 14603
rect 9309 14563 9367 14569
rect 10686 14560 10692 14612
rect 10744 14600 10750 14612
rect 12621 14603 12679 14609
rect 12621 14600 12633 14603
rect 10744 14572 12633 14600
rect 10744 14560 10750 14572
rect 12621 14569 12633 14572
rect 12667 14569 12679 14603
rect 13538 14600 13544 14612
rect 13499 14572 13544 14600
rect 12621 14563 12679 14569
rect 13538 14560 13544 14572
rect 13596 14560 13602 14612
rect 17310 14600 17316 14612
rect 13832 14572 17316 14600
rect 13170 14492 13176 14544
rect 13228 14532 13234 14544
rect 13832 14532 13860 14572
rect 17310 14560 17316 14572
rect 17368 14560 17374 14612
rect 17402 14560 17408 14612
rect 17460 14600 17466 14612
rect 17865 14603 17923 14609
rect 17865 14600 17877 14603
rect 17460 14572 17877 14600
rect 17460 14560 17466 14572
rect 17865 14569 17877 14572
rect 17911 14569 17923 14603
rect 22002 14600 22008 14612
rect 17865 14563 17923 14569
rect 19260 14572 22008 14600
rect 13228 14504 13860 14532
rect 17221 14535 17279 14541
rect 13228 14492 13234 14504
rect 17221 14501 17233 14535
rect 17267 14532 17279 14535
rect 18782 14532 18788 14544
rect 17267 14504 18788 14532
rect 17267 14501 17279 14504
rect 17221 14495 17279 14501
rect 18782 14492 18788 14504
rect 18840 14492 18846 14544
rect 10318 14424 10324 14476
rect 10376 14464 10382 14476
rect 10413 14467 10471 14473
rect 10413 14464 10425 14467
rect 10376 14436 10425 14464
rect 10376 14424 10382 14436
rect 10413 14433 10425 14436
rect 10459 14433 10471 14467
rect 13188 14464 13216 14492
rect 14090 14464 14096 14476
rect 10413 14427 10471 14433
rect 12728 14436 13216 14464
rect 14051 14436 14096 14464
rect 7742 14396 7748 14408
rect 7703 14368 7748 14396
rect 7742 14356 7748 14368
rect 7800 14356 7806 14408
rect 8389 14399 8447 14405
rect 8389 14365 8401 14399
rect 8435 14396 8447 14399
rect 9306 14396 9312 14408
rect 8435 14368 9312 14396
rect 8435 14365 8447 14368
rect 8389 14359 8447 14365
rect 9306 14356 9312 14368
rect 9364 14356 9370 14408
rect 9953 14399 10011 14405
rect 9953 14365 9965 14399
rect 9999 14396 10011 14399
rect 11606 14396 11612 14408
rect 9999 14368 11612 14396
rect 9999 14365 10011 14368
rect 9953 14359 10011 14365
rect 11606 14356 11612 14368
rect 11664 14356 11670 14408
rect 12526 14396 12532 14408
rect 12487 14368 12532 14396
rect 12526 14356 12532 14368
rect 12584 14356 12590 14408
rect 12728 14405 12756 14436
rect 14090 14424 14096 14436
rect 14148 14424 14154 14476
rect 16206 14424 16212 14476
rect 16264 14464 16270 14476
rect 16264 14436 16804 14464
rect 16264 14424 16270 14436
rect 12713 14399 12771 14405
rect 12713 14365 12725 14399
rect 12759 14365 12771 14399
rect 12713 14359 12771 14365
rect 13173 14399 13231 14405
rect 13173 14365 13185 14399
rect 13219 14396 13231 14399
rect 13262 14396 13268 14408
rect 13219 14368 13268 14396
rect 13219 14365 13231 14368
rect 13173 14359 13231 14365
rect 13262 14356 13268 14368
rect 13320 14356 13326 14408
rect 13354 14356 13360 14408
rect 13412 14396 13418 14408
rect 14182 14396 14188 14408
rect 13412 14368 14188 14396
rect 13412 14356 13418 14368
rect 14182 14356 14188 14368
rect 14240 14356 14246 14408
rect 14366 14405 14372 14408
rect 14360 14396 14372 14405
rect 14327 14368 14372 14396
rect 14360 14359 14372 14368
rect 14366 14356 14372 14359
rect 14424 14356 14430 14408
rect 15933 14399 15991 14405
rect 15933 14396 15945 14399
rect 15488 14368 15945 14396
rect 8941 14331 8999 14337
rect 8941 14297 8953 14331
rect 8987 14297 8999 14331
rect 8941 14291 8999 14297
rect 9125 14331 9183 14337
rect 9125 14297 9137 14331
rect 9171 14328 9183 14331
rect 9214 14328 9220 14340
rect 9171 14300 9220 14328
rect 9171 14297 9183 14300
rect 9125 14291 9183 14297
rect 8956 14260 8984 14291
rect 9214 14288 9220 14300
rect 9272 14288 9278 14340
rect 10502 14328 10508 14340
rect 9324 14300 10508 14328
rect 9324 14260 9352 14300
rect 10502 14288 10508 14300
rect 10560 14288 10566 14340
rect 10680 14331 10738 14337
rect 10680 14297 10692 14331
rect 10726 14328 10738 14331
rect 10870 14328 10876 14340
rect 10726 14300 10876 14328
rect 10726 14297 10738 14300
rect 10680 14291 10738 14297
rect 10870 14288 10876 14300
rect 10928 14288 10934 14340
rect 13722 14288 13728 14340
rect 13780 14328 13786 14340
rect 15102 14328 15108 14340
rect 13780 14300 15108 14328
rect 13780 14288 13786 14300
rect 15102 14288 15108 14300
rect 15160 14288 15166 14340
rect 15488 14272 15516 14368
rect 15933 14365 15945 14368
rect 15979 14365 15991 14399
rect 16574 14396 16580 14408
rect 16535 14368 16580 14396
rect 15933 14359 15991 14365
rect 16574 14356 16580 14368
rect 16632 14356 16638 14408
rect 16670 14399 16728 14405
rect 16670 14365 16682 14399
rect 16716 14365 16728 14399
rect 16776 14396 16804 14436
rect 16850 14424 16856 14476
rect 16908 14464 16914 14476
rect 19260 14473 19288 14572
rect 22002 14560 22008 14572
rect 22060 14600 22066 14612
rect 23477 14603 23535 14609
rect 23477 14600 23489 14603
rect 22060 14572 23489 14600
rect 22060 14560 22066 14572
rect 23477 14569 23489 14572
rect 23523 14569 23535 14603
rect 24854 14600 24860 14612
rect 24815 14572 24860 14600
rect 23477 14563 23535 14569
rect 24854 14560 24860 14572
rect 24912 14560 24918 14612
rect 24946 14560 24952 14612
rect 25004 14600 25010 14612
rect 25225 14603 25283 14609
rect 25225 14600 25237 14603
rect 25004 14572 25237 14600
rect 25004 14560 25010 14572
rect 25225 14569 25237 14572
rect 25271 14569 25283 14603
rect 26970 14600 26976 14612
rect 25225 14563 25283 14569
rect 26712 14572 26976 14600
rect 21269 14535 21327 14541
rect 21269 14501 21281 14535
rect 21315 14532 21327 14535
rect 21358 14532 21364 14544
rect 21315 14504 21364 14532
rect 21315 14501 21327 14504
rect 21269 14495 21327 14501
rect 21358 14492 21364 14504
rect 21416 14492 21422 14544
rect 19245 14467 19303 14473
rect 16908 14436 17724 14464
rect 16908 14424 16914 14436
rect 17126 14405 17132 14408
rect 16945 14399 17003 14405
rect 16945 14396 16957 14399
rect 16776 14368 16957 14396
rect 16670 14359 16728 14365
rect 16945 14365 16957 14368
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 17083 14399 17132 14405
rect 17083 14365 17095 14399
rect 17129 14365 17132 14399
rect 17083 14359 17132 14365
rect 15562 14288 15568 14340
rect 15620 14328 15626 14340
rect 16685 14328 16713 14359
rect 17126 14356 17132 14359
rect 17184 14396 17190 14408
rect 17184 14368 17637 14396
rect 17184 14356 17190 14368
rect 15620 14300 16713 14328
rect 16853 14331 16911 14337
rect 15620 14288 15626 14300
rect 16853 14297 16865 14331
rect 16899 14328 16911 14331
rect 17218 14328 17224 14340
rect 16899 14300 17224 14328
rect 16899 14297 16911 14300
rect 16853 14291 16911 14297
rect 17218 14288 17224 14300
rect 17276 14288 17282 14340
rect 8956 14232 9352 14260
rect 9769 14263 9827 14269
rect 9769 14229 9781 14263
rect 9815 14260 9827 14263
rect 10594 14260 10600 14272
rect 9815 14232 10600 14260
rect 9815 14229 9827 14232
rect 9769 14223 9827 14229
rect 10594 14220 10600 14232
rect 10652 14220 10658 14272
rect 11698 14220 11704 14272
rect 11756 14260 11762 14272
rect 11793 14263 11851 14269
rect 11793 14260 11805 14263
rect 11756 14232 11805 14260
rect 11756 14220 11762 14232
rect 11793 14229 11805 14232
rect 11839 14229 11851 14263
rect 15470 14260 15476 14272
rect 15431 14232 15476 14260
rect 11793 14223 11851 14229
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 16022 14260 16028 14272
rect 15983 14232 16028 14260
rect 16022 14220 16028 14232
rect 16080 14220 16086 14272
rect 17609 14260 17637 14368
rect 17696 14337 17724 14436
rect 19245 14433 19257 14467
rect 19291 14433 19303 14467
rect 19245 14427 19303 14433
rect 20346 14424 20352 14476
rect 20404 14464 20410 14476
rect 22462 14464 22468 14476
rect 20404 14436 22048 14464
rect 22423 14436 22468 14464
rect 20404 14424 20410 14436
rect 17770 14356 17776 14408
rect 17828 14396 17834 14408
rect 18693 14399 18751 14405
rect 18693 14396 18705 14399
rect 17828 14368 18705 14396
rect 17828 14356 17834 14368
rect 18693 14365 18705 14368
rect 18739 14365 18751 14399
rect 18693 14359 18751 14365
rect 19512 14399 19570 14405
rect 19512 14365 19524 14399
rect 19558 14396 19570 14399
rect 20806 14396 20812 14408
rect 19558 14368 20812 14396
rect 19558 14365 19570 14368
rect 19512 14359 19570 14365
rect 20806 14356 20812 14368
rect 20864 14356 20870 14408
rect 21100 14405 21128 14436
rect 21085 14399 21143 14405
rect 21085 14365 21097 14399
rect 21131 14365 21143 14399
rect 21818 14396 21824 14408
rect 21779 14368 21824 14396
rect 21085 14359 21143 14365
rect 21818 14356 21824 14368
rect 21876 14356 21882 14408
rect 22020 14405 22048 14436
rect 22462 14424 22468 14436
rect 22520 14424 22526 14476
rect 25317 14467 25375 14473
rect 25317 14433 25329 14467
rect 25363 14464 25375 14467
rect 25682 14464 25688 14476
rect 25363 14436 25688 14464
rect 25363 14433 25375 14436
rect 25317 14427 25375 14433
rect 25682 14424 25688 14436
rect 25740 14464 25746 14476
rect 26050 14464 26056 14476
rect 25740 14436 26056 14464
rect 25740 14424 25746 14436
rect 26050 14424 26056 14436
rect 26108 14424 26114 14476
rect 26712 14473 26740 14572
rect 26970 14560 26976 14572
rect 27028 14560 27034 14612
rect 28074 14600 28080 14612
rect 27987 14572 28080 14600
rect 28074 14560 28080 14572
rect 28132 14600 28138 14612
rect 28442 14600 28448 14612
rect 28132 14572 28448 14600
rect 28132 14560 28138 14572
rect 28442 14560 28448 14572
rect 28500 14560 28506 14612
rect 26697 14467 26755 14473
rect 26697 14433 26709 14467
rect 26743 14433 26755 14467
rect 26697 14427 26755 14433
rect 22005 14399 22063 14405
rect 22005 14365 22017 14399
rect 22051 14365 22063 14399
rect 22646 14396 22652 14408
rect 22607 14368 22652 14396
rect 22005 14359 22063 14365
rect 22646 14356 22652 14368
rect 22704 14356 22710 14408
rect 23385 14399 23443 14405
rect 23385 14365 23397 14399
rect 23431 14396 23443 14399
rect 23474 14396 23480 14408
rect 23431 14368 23480 14396
rect 23431 14365 23443 14368
rect 23385 14359 23443 14365
rect 23474 14356 23480 14368
rect 23532 14356 23538 14408
rect 25038 14396 25044 14408
rect 24999 14368 25044 14396
rect 25038 14356 25044 14368
rect 25096 14356 25102 14408
rect 26964 14399 27022 14405
rect 26964 14365 26976 14399
rect 27010 14396 27022 14399
rect 28350 14396 28356 14408
rect 27010 14368 28356 14396
rect 27010 14365 27022 14368
rect 26964 14359 27022 14365
rect 28350 14356 28356 14368
rect 28408 14356 28414 14408
rect 17681 14331 17739 14337
rect 17681 14297 17693 14331
rect 17727 14297 17739 14331
rect 17681 14291 17739 14297
rect 17862 14288 17868 14340
rect 17920 14337 17926 14340
rect 17920 14331 17939 14337
rect 17927 14297 17939 14331
rect 21726 14328 21732 14340
rect 17920 14291 17939 14297
rect 18064 14300 21732 14328
rect 17920 14288 17926 14291
rect 17880 14260 17908 14288
rect 18064 14269 18092 14300
rect 21726 14288 21732 14300
rect 21784 14288 21790 14340
rect 21913 14331 21971 14337
rect 21913 14297 21925 14331
rect 21959 14328 21971 14331
rect 23842 14328 23848 14340
rect 21959 14300 23848 14328
rect 21959 14297 21971 14300
rect 21913 14291 21971 14297
rect 23842 14288 23848 14300
rect 23900 14288 23906 14340
rect 17609 14232 17908 14260
rect 18049 14263 18107 14269
rect 18049 14229 18061 14263
rect 18095 14229 18107 14263
rect 18506 14260 18512 14272
rect 18467 14232 18512 14260
rect 18049 14223 18107 14229
rect 18506 14220 18512 14232
rect 18564 14220 18570 14272
rect 20070 14220 20076 14272
rect 20128 14260 20134 14272
rect 20625 14263 20683 14269
rect 20625 14260 20637 14263
rect 20128 14232 20637 14260
rect 20128 14220 20134 14232
rect 20625 14229 20637 14232
rect 20671 14229 20683 14263
rect 20625 14223 20683 14229
rect 22462 14220 22468 14272
rect 22520 14260 22526 14272
rect 22833 14263 22891 14269
rect 22833 14260 22845 14263
rect 22520 14232 22845 14260
rect 22520 14220 22526 14232
rect 22833 14229 22845 14232
rect 22879 14229 22891 14263
rect 22833 14223 22891 14229
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 9214 14056 9220 14068
rect 9175 14028 9220 14056
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 10318 14056 10324 14068
rect 10279 14028 10324 14056
rect 10318 14016 10324 14028
rect 10376 14016 10382 14068
rect 14093 14059 14151 14065
rect 14093 14025 14105 14059
rect 14139 14056 14151 14059
rect 14826 14056 14832 14068
rect 14139 14028 14832 14056
rect 14139 14025 14151 14028
rect 14093 14019 14151 14025
rect 14826 14016 14832 14028
rect 14884 14016 14890 14068
rect 14918 14016 14924 14068
rect 14976 14056 14982 14068
rect 15565 14059 15623 14065
rect 14976 14028 15056 14056
rect 14976 14016 14982 14028
rect 8202 13988 8208 14000
rect 7944 13960 8208 13988
rect 7834 13920 7840 13932
rect 7747 13892 7840 13920
rect 7834 13880 7840 13892
rect 7892 13920 7898 13932
rect 7944 13920 7972 13960
rect 8202 13948 8208 13960
rect 8260 13948 8266 14000
rect 11514 13988 11520 14000
rect 11475 13960 11520 13988
rect 11514 13948 11520 13960
rect 11572 13948 11578 14000
rect 11733 13991 11791 13997
rect 11733 13957 11745 13991
rect 11779 13988 11791 13991
rect 12434 13988 12440 14000
rect 11779 13960 12440 13988
rect 11779 13957 11791 13960
rect 11733 13951 11791 13957
rect 12434 13948 12440 13960
rect 12492 13988 12498 14000
rect 13262 13988 13268 14000
rect 12492 13960 13268 13988
rect 12492 13948 12498 13960
rect 13262 13948 13268 13960
rect 13320 13988 13326 14000
rect 13725 13991 13783 13997
rect 13725 13988 13737 13991
rect 13320 13960 13737 13988
rect 13320 13948 13326 13960
rect 13725 13957 13737 13960
rect 13771 13957 13783 13991
rect 13725 13951 13783 13957
rect 14642 13948 14648 14000
rect 14700 13988 14706 14000
rect 14700 13960 14852 13988
rect 14700 13948 14706 13960
rect 8110 13929 8116 13932
rect 8104 13920 8116 13929
rect 7892 13892 7972 13920
rect 8071 13892 8116 13920
rect 7892 13880 7898 13892
rect 8104 13883 8116 13892
rect 8110 13880 8116 13883
rect 8168 13880 8174 13932
rect 10229 13923 10287 13929
rect 10229 13889 10241 13923
rect 10275 13920 10287 13923
rect 10962 13920 10968 13932
rect 10275 13892 10968 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 10962 13880 10968 13892
rect 11020 13880 11026 13932
rect 12618 13920 12624 13932
rect 12579 13892 12624 13920
rect 12618 13880 12624 13892
rect 12676 13880 12682 13932
rect 12802 13920 12808 13932
rect 12763 13892 12808 13920
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 13909 13923 13967 13929
rect 13909 13889 13921 13923
rect 13955 13920 13967 13923
rect 14458 13920 14464 13932
rect 13955 13892 14464 13920
rect 13955 13889 13967 13892
rect 13909 13883 13967 13889
rect 14458 13880 14464 13892
rect 14516 13880 14522 13932
rect 14824 13929 14852 13960
rect 14818 13923 14876 13929
rect 14818 13889 14830 13923
rect 14864 13889 14876 13923
rect 15028 13920 15056 14028
rect 15565 14025 15577 14059
rect 15611 14056 15623 14059
rect 16574 14056 16580 14068
rect 15611 14028 16580 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 16574 14016 16580 14028
rect 16632 14016 16638 14068
rect 17037 14059 17095 14065
rect 17037 14025 17049 14059
rect 17083 14056 17095 14059
rect 25314 14056 25320 14068
rect 17083 14028 25320 14056
rect 17083 14025 17095 14028
rect 17037 14019 17095 14025
rect 25314 14016 25320 14028
rect 25372 14016 25378 14068
rect 26237 14059 26295 14065
rect 26237 14025 26249 14059
rect 26283 14056 26295 14059
rect 26418 14056 26424 14068
rect 26283 14028 26424 14056
rect 26283 14025 26295 14028
rect 26237 14019 26295 14025
rect 26418 14016 26424 14028
rect 26476 14016 26482 14068
rect 16669 13991 16727 13997
rect 16669 13957 16681 13991
rect 16715 13957 16727 13991
rect 16669 13951 16727 13957
rect 16885 13991 16943 13997
rect 16885 13957 16897 13991
rect 16931 13988 16943 13991
rect 16931 13960 17448 13988
rect 16931 13957 16943 13960
rect 16885 13951 16943 13957
rect 14366 13812 14372 13864
rect 14424 13852 14430 13864
rect 14568 13858 14701 13886
rect 14818 13883 14876 13889
rect 14936 13892 15056 13920
rect 14936 13861 14964 13892
rect 15654 13880 15660 13932
rect 15712 13920 15718 13932
rect 15841 13923 15899 13929
rect 15841 13920 15853 13923
rect 15712 13892 15853 13920
rect 15712 13880 15718 13892
rect 15841 13889 15853 13892
rect 15887 13889 15899 13923
rect 15841 13883 15899 13889
rect 16025 13923 16083 13929
rect 16025 13889 16037 13923
rect 16071 13920 16083 13923
rect 16114 13920 16120 13932
rect 16071 13892 16120 13920
rect 16071 13889 16083 13892
rect 16025 13883 16083 13889
rect 16114 13880 16120 13892
rect 16172 13880 16178 13932
rect 16684 13920 16712 13951
rect 17034 13920 17040 13932
rect 16684 13892 17040 13920
rect 17034 13880 17040 13892
rect 17092 13880 17098 13932
rect 17420 13920 17448 13960
rect 17494 13948 17500 14000
rect 17552 13988 17558 14000
rect 17713 13991 17771 13997
rect 17552 13960 17597 13988
rect 17552 13948 17558 13960
rect 17713 13957 17725 13991
rect 17759 13988 17771 13991
rect 18138 13988 18144 14000
rect 17759 13960 18144 13988
rect 17759 13957 17771 13960
rect 17713 13951 17771 13957
rect 17728 13920 17756 13951
rect 18138 13948 18144 13960
rect 18196 13948 18202 14000
rect 20349 13991 20407 13997
rect 20349 13988 20361 13991
rect 19168 13960 20361 13988
rect 17420 13892 17756 13920
rect 18046 13880 18052 13932
rect 18104 13920 18110 13932
rect 19168 13929 19196 13960
rect 20349 13957 20361 13960
rect 20395 13957 20407 13991
rect 20349 13951 20407 13957
rect 20530 13948 20536 14000
rect 20588 13988 20594 14000
rect 21177 13991 21235 13997
rect 21177 13988 21189 13991
rect 20588 13960 21189 13988
rect 20588 13948 20594 13960
rect 21177 13957 21189 13960
rect 21223 13957 21235 13991
rect 22088 13991 22146 13997
rect 21177 13951 21235 13957
rect 21744 13960 22048 13988
rect 18509 13923 18567 13929
rect 18509 13920 18521 13923
rect 18104 13892 18521 13920
rect 18104 13880 18110 13892
rect 18509 13889 18521 13892
rect 18555 13889 18567 13923
rect 18509 13883 18567 13889
rect 19153 13923 19211 13929
rect 19153 13889 19165 13923
rect 19199 13889 19211 13923
rect 19153 13883 19211 13889
rect 19242 13880 19248 13932
rect 19300 13920 19306 13932
rect 19521 13923 19579 13929
rect 19300 13892 19345 13920
rect 19300 13880 19306 13892
rect 19521 13889 19533 13923
rect 19567 13920 19579 13923
rect 20070 13920 20076 13932
rect 19567 13892 20076 13920
rect 19567 13889 19579 13892
rect 19521 13883 19579 13889
rect 20070 13880 20076 13892
rect 20128 13880 20134 13932
rect 20165 13923 20223 13929
rect 20165 13889 20177 13923
rect 20211 13920 20223 13923
rect 20993 13923 21051 13929
rect 20993 13920 21005 13923
rect 20211 13892 21005 13920
rect 20211 13889 20223 13892
rect 20165 13883 20223 13889
rect 14568 13852 14596 13858
rect 14424 13824 14596 13852
rect 14673 13852 14701 13858
rect 14738 13855 14796 13861
rect 14738 13852 14750 13855
rect 14673 13824 14750 13852
rect 14424 13812 14430 13824
rect 14738 13821 14750 13824
rect 14784 13821 14796 13855
rect 14738 13815 14796 13821
rect 14912 13855 14970 13861
rect 14912 13821 14924 13855
rect 14958 13821 14970 13855
rect 14912 13815 14970 13821
rect 15013 13855 15071 13861
rect 15013 13821 15025 13855
rect 15059 13852 15071 13855
rect 15470 13852 15476 13864
rect 15059 13824 15476 13852
rect 15059 13821 15071 13824
rect 15013 13815 15071 13821
rect 15470 13812 15476 13824
rect 15528 13812 15534 13864
rect 15749 13855 15807 13861
rect 15749 13821 15761 13855
rect 15795 13821 15807 13855
rect 15749 13815 15807 13821
rect 15933 13855 15991 13861
rect 15933 13821 15945 13855
rect 15979 13852 15991 13855
rect 16298 13852 16304 13864
rect 15979 13824 16304 13852
rect 15979 13821 15991 13824
rect 15933 13815 15991 13821
rect 14553 13787 14611 13793
rect 14553 13753 14565 13787
rect 14599 13784 14611 13787
rect 15194 13784 15200 13796
rect 14599 13756 15200 13784
rect 14599 13753 14611 13756
rect 14553 13747 14611 13753
rect 15194 13744 15200 13756
rect 15252 13744 15258 13796
rect 15764 13784 15792 13815
rect 16298 13812 16304 13824
rect 16356 13812 16362 13864
rect 17494 13852 17500 13864
rect 16685 13824 17500 13852
rect 16685 13784 16713 13824
rect 17494 13812 17500 13824
rect 17552 13852 17558 13864
rect 18414 13852 18420 13864
rect 17552 13824 18420 13852
rect 17552 13812 17558 13824
rect 18414 13812 18420 13824
rect 18472 13812 18478 13864
rect 18969 13855 19027 13861
rect 18969 13821 18981 13855
rect 19015 13852 19027 13855
rect 19334 13852 19340 13864
rect 19015 13824 19340 13852
rect 19015 13821 19027 13824
rect 18969 13815 19027 13821
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 19981 13855 20039 13861
rect 19981 13821 19993 13855
rect 20027 13852 20039 13855
rect 20622 13852 20628 13864
rect 20027 13824 20628 13852
rect 20027 13821 20039 13824
rect 19981 13815 20039 13821
rect 20622 13812 20628 13824
rect 20680 13812 20686 13864
rect 20732 13784 20760 13892
rect 20993 13889 21005 13892
rect 21039 13920 21051 13923
rect 21744 13920 21772 13960
rect 21039 13892 21772 13920
rect 21821 13923 21879 13929
rect 21039 13889 21051 13892
rect 20993 13883 21051 13889
rect 21821 13889 21833 13923
rect 21867 13920 21879 13923
rect 21910 13920 21916 13932
rect 21867 13892 21916 13920
rect 21867 13889 21879 13892
rect 21821 13883 21879 13889
rect 21910 13880 21916 13892
rect 21968 13880 21974 13932
rect 22020 13920 22048 13960
rect 22088 13957 22100 13991
rect 22134 13988 22146 13991
rect 23290 13988 23296 14000
rect 22134 13960 23296 13988
rect 22134 13957 22146 13960
rect 22088 13951 22146 13957
rect 23290 13948 23296 13960
rect 23348 13948 23354 14000
rect 24578 13988 24584 14000
rect 23676 13960 24584 13988
rect 22646 13920 22652 13932
rect 22020 13892 22652 13920
rect 22646 13880 22652 13892
rect 22704 13880 22710 13932
rect 23676 13929 23704 13960
rect 24578 13948 24584 13960
rect 24636 13948 24642 14000
rect 25961 13991 26019 13997
rect 25961 13957 25973 13991
rect 26007 13988 26019 13991
rect 27522 13988 27528 14000
rect 26007 13960 27528 13988
rect 26007 13957 26019 13960
rect 25961 13951 26019 13957
rect 27522 13948 27528 13960
rect 27580 13948 27586 14000
rect 23934 13929 23940 13932
rect 23661 13923 23719 13929
rect 23661 13889 23673 13923
rect 23707 13889 23719 13923
rect 23928 13920 23940 13929
rect 23895 13892 23940 13920
rect 23661 13883 23719 13889
rect 23928 13883 23940 13892
rect 23934 13880 23940 13883
rect 23992 13880 23998 13932
rect 25590 13920 25596 13932
rect 25551 13892 25596 13920
rect 25590 13880 25596 13892
rect 25648 13880 25654 13932
rect 25682 13880 25688 13932
rect 25740 13920 25746 13932
rect 25740 13892 25785 13920
rect 25740 13880 25746 13892
rect 25866 13880 25872 13932
rect 25924 13920 25930 13932
rect 25924 13892 25969 13920
rect 25924 13880 25930 13892
rect 26050 13880 26056 13932
rect 26108 13929 26114 13932
rect 26108 13920 26116 13929
rect 27157 13923 27215 13929
rect 26108 13892 26153 13920
rect 26108 13883 26116 13892
rect 27157 13889 27169 13923
rect 27203 13889 27215 13923
rect 27157 13883 27215 13889
rect 26108 13880 26114 13883
rect 20809 13855 20867 13861
rect 20809 13821 20821 13855
rect 20855 13852 20867 13855
rect 20898 13852 20904 13864
rect 20855 13824 20904 13852
rect 20855 13821 20867 13824
rect 20809 13815 20867 13821
rect 20898 13812 20904 13824
rect 20956 13812 20962 13864
rect 27172 13852 27200 13883
rect 25792 13824 27200 13852
rect 25792 13796 25820 13824
rect 15764 13756 16713 13784
rect 16776 13756 20760 13784
rect 11698 13716 11704 13728
rect 11659 13688 11704 13716
rect 11698 13676 11704 13688
rect 11756 13676 11762 13728
rect 11882 13716 11888 13728
rect 11843 13688 11888 13716
rect 11882 13676 11888 13688
rect 11940 13676 11946 13728
rect 12621 13719 12679 13725
rect 12621 13685 12633 13719
rect 12667 13716 12679 13719
rect 13906 13716 13912 13728
rect 12667 13688 13912 13716
rect 12667 13685 12679 13688
rect 12621 13679 12679 13685
rect 13906 13676 13912 13688
rect 13964 13676 13970 13728
rect 14274 13676 14280 13728
rect 14332 13716 14338 13728
rect 16776 13716 16804 13756
rect 25774 13744 25780 13796
rect 25832 13744 25838 13796
rect 14332 13688 16804 13716
rect 16853 13719 16911 13725
rect 14332 13676 14338 13688
rect 16853 13685 16865 13719
rect 16899 13716 16911 13719
rect 17034 13716 17040 13728
rect 16899 13688 17040 13716
rect 16899 13685 16911 13688
rect 16853 13679 16911 13685
rect 17034 13676 17040 13688
rect 17092 13676 17098 13728
rect 17494 13676 17500 13728
rect 17552 13716 17558 13728
rect 17681 13719 17739 13725
rect 17681 13716 17693 13719
rect 17552 13688 17693 13716
rect 17552 13676 17558 13688
rect 17681 13685 17693 13688
rect 17727 13685 17739 13719
rect 17862 13716 17868 13728
rect 17823 13688 17868 13716
rect 17681 13679 17739 13685
rect 17862 13676 17868 13688
rect 17920 13676 17926 13728
rect 18138 13676 18144 13728
rect 18196 13716 18202 13728
rect 18325 13719 18383 13725
rect 18325 13716 18337 13719
rect 18196 13688 18337 13716
rect 18196 13676 18202 13688
rect 18325 13685 18337 13688
rect 18371 13685 18383 13719
rect 18325 13679 18383 13685
rect 18414 13676 18420 13728
rect 18472 13716 18478 13728
rect 19429 13719 19487 13725
rect 19429 13716 19441 13719
rect 18472 13688 19441 13716
rect 18472 13676 18478 13688
rect 19429 13685 19441 13688
rect 19475 13685 19487 13719
rect 19429 13679 19487 13685
rect 19518 13676 19524 13728
rect 19576 13716 19582 13728
rect 21082 13716 21088 13728
rect 19576 13688 21088 13716
rect 19576 13676 19582 13688
rect 21082 13676 21088 13688
rect 21140 13716 21146 13728
rect 21818 13716 21824 13728
rect 21140 13688 21824 13716
rect 21140 13676 21146 13688
rect 21818 13676 21824 13688
rect 21876 13676 21882 13728
rect 22186 13676 22192 13728
rect 22244 13716 22250 13728
rect 23201 13719 23259 13725
rect 23201 13716 23213 13719
rect 22244 13688 23213 13716
rect 22244 13676 22250 13688
rect 23201 13685 23213 13688
rect 23247 13685 23259 13719
rect 23201 13679 23259 13685
rect 24946 13676 24952 13728
rect 25004 13716 25010 13728
rect 25041 13719 25099 13725
rect 25041 13716 25053 13719
rect 25004 13688 25053 13716
rect 25004 13676 25010 13688
rect 25041 13685 25053 13688
rect 25087 13685 25099 13719
rect 25041 13679 25099 13685
rect 26234 13676 26240 13728
rect 26292 13716 26298 13728
rect 26973 13719 27031 13725
rect 26973 13716 26985 13719
rect 26292 13688 26985 13716
rect 26292 13676 26298 13688
rect 26973 13685 26985 13688
rect 27019 13685 27031 13719
rect 26973 13679 27031 13685
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 11793 13515 11851 13521
rect 11793 13481 11805 13515
rect 11839 13512 11851 13515
rect 12437 13515 12495 13521
rect 12437 13512 12449 13515
rect 11839 13484 12449 13512
rect 11839 13481 11851 13484
rect 11793 13475 11851 13481
rect 12437 13481 12449 13484
rect 12483 13481 12495 13515
rect 12437 13475 12495 13481
rect 12526 13472 12532 13524
rect 12584 13512 12590 13524
rect 14274 13512 14280 13524
rect 12584 13484 12756 13512
rect 14235 13484 14280 13512
rect 12584 13472 12590 13484
rect 11422 13404 11428 13456
rect 11480 13444 11486 13456
rect 12621 13447 12679 13453
rect 12621 13444 12633 13447
rect 11480 13416 12633 13444
rect 11480 13404 11486 13416
rect 12621 13413 12633 13416
rect 12667 13413 12679 13447
rect 12728 13444 12756 13484
rect 14274 13472 14280 13484
rect 14332 13472 14338 13524
rect 14642 13472 14648 13524
rect 14700 13512 14706 13524
rect 15838 13512 15844 13524
rect 14700 13484 15844 13512
rect 14700 13472 14706 13484
rect 15838 13472 15844 13484
rect 15896 13512 15902 13524
rect 16209 13515 16267 13521
rect 16209 13512 16221 13515
rect 15896 13484 16221 13512
rect 15896 13472 15902 13484
rect 16209 13481 16221 13484
rect 16255 13481 16267 13515
rect 16209 13475 16267 13481
rect 16393 13515 16451 13521
rect 16393 13481 16405 13515
rect 16439 13512 16451 13515
rect 16666 13512 16672 13524
rect 16439 13484 16672 13512
rect 16439 13481 16451 13484
rect 16393 13475 16451 13481
rect 16666 13472 16672 13484
rect 16724 13472 16730 13524
rect 17034 13512 17040 13524
rect 16995 13484 17040 13512
rect 17034 13472 17040 13484
rect 17092 13512 17098 13524
rect 17586 13512 17592 13524
rect 17092 13484 17592 13512
rect 17092 13472 17098 13484
rect 17586 13472 17592 13484
rect 17644 13512 17650 13524
rect 18141 13515 18199 13521
rect 18141 13512 18153 13515
rect 17644 13484 18153 13512
rect 17644 13472 17650 13484
rect 18141 13481 18153 13484
rect 18187 13512 18199 13515
rect 18506 13512 18512 13524
rect 18187 13484 18512 13512
rect 18187 13481 18199 13484
rect 18141 13475 18199 13481
rect 18506 13472 18512 13484
rect 18564 13472 18570 13524
rect 19429 13515 19487 13521
rect 19429 13481 19441 13515
rect 19475 13512 19487 13515
rect 19518 13512 19524 13524
rect 19475 13484 19524 13512
rect 19475 13481 19487 13484
rect 19429 13475 19487 13481
rect 19518 13472 19524 13484
rect 19576 13472 19582 13524
rect 19613 13515 19671 13521
rect 19613 13481 19625 13515
rect 19659 13512 19671 13515
rect 20622 13512 20628 13524
rect 19659 13484 20628 13512
rect 19659 13481 19671 13484
rect 19613 13475 19671 13481
rect 20622 13472 20628 13484
rect 20680 13472 20686 13524
rect 22554 13512 22560 13524
rect 20916 13484 22560 13512
rect 14461 13447 14519 13453
rect 14461 13444 14473 13447
rect 12728 13416 14473 13444
rect 12621 13407 12679 13413
rect 14461 13413 14473 13416
rect 14507 13413 14519 13447
rect 14461 13407 14519 13413
rect 15102 13404 15108 13456
rect 15160 13444 15166 13456
rect 15160 13416 16436 13444
rect 15160 13404 15166 13416
rect 9398 13336 9404 13388
rect 9456 13376 9462 13388
rect 10318 13376 10324 13388
rect 9456 13348 10324 13376
rect 9456 13336 9462 13348
rect 10318 13336 10324 13348
rect 10376 13376 10382 13388
rect 10413 13379 10471 13385
rect 10413 13376 10425 13379
rect 10376 13348 10425 13376
rect 10376 13336 10382 13348
rect 10413 13345 10425 13348
rect 10459 13345 10471 13379
rect 10413 13339 10471 13345
rect 12802 13336 12808 13388
rect 12860 13376 12866 13388
rect 12860 13348 14320 13376
rect 12860 13336 12866 13348
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13308 8447 13311
rect 12158 13308 12164 13320
rect 8435 13280 12164 13308
rect 8435 13277 8447 13280
rect 8389 13271 8447 13277
rect 12158 13268 12164 13280
rect 12216 13268 12222 13320
rect 13170 13308 13176 13320
rect 13131 13280 13176 13308
rect 13170 13268 13176 13280
rect 13228 13268 13234 13320
rect 14090 13308 14096 13320
rect 14051 13280 14096 13308
rect 14090 13268 14096 13280
rect 14148 13268 14154 13320
rect 14292 13317 14320 13348
rect 16298 13336 16304 13388
rect 16356 13336 16362 13388
rect 14277 13311 14335 13317
rect 14277 13277 14289 13311
rect 14323 13308 14335 13311
rect 14458 13308 14464 13320
rect 14323 13280 14464 13308
rect 14323 13277 14335 13280
rect 14277 13271 14335 13277
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 15378 13308 15384 13320
rect 15339 13280 15384 13308
rect 15378 13268 15384 13280
rect 15436 13268 15442 13320
rect 16316 13308 16344 13336
rect 16040 13280 16344 13308
rect 9306 13240 9312 13252
rect 9267 13212 9312 13240
rect 9306 13200 9312 13212
rect 9364 13200 9370 13252
rect 9493 13243 9551 13249
rect 9493 13209 9505 13243
rect 9539 13240 9551 13243
rect 9858 13240 9864 13252
rect 9539 13212 9864 13240
rect 9539 13209 9551 13212
rect 9493 13203 9551 13209
rect 9858 13200 9864 13212
rect 9916 13200 9922 13252
rect 10680 13243 10738 13249
rect 10680 13209 10692 13243
rect 10726 13240 10738 13243
rect 10778 13240 10784 13252
rect 10726 13212 10784 13240
rect 10726 13209 10738 13212
rect 10680 13203 10738 13209
rect 10778 13200 10784 13212
rect 10836 13200 10842 13252
rect 11514 13200 11520 13252
rect 11572 13240 11578 13252
rect 12250 13240 12256 13252
rect 11572 13212 12256 13240
rect 11572 13200 11578 13212
rect 12250 13200 12256 13212
rect 12308 13200 12314 13252
rect 12434 13200 12440 13252
rect 12492 13249 12498 13252
rect 12492 13243 12511 13249
rect 12499 13209 12511 13243
rect 12492 13203 12511 13209
rect 12492 13200 12498 13203
rect 13262 13200 13268 13252
rect 13320 13240 13326 13252
rect 13541 13243 13599 13249
rect 13541 13240 13553 13243
rect 13320 13212 13553 13240
rect 13320 13200 13326 13212
rect 13541 13209 13553 13212
rect 13587 13240 13599 13243
rect 14550 13240 14556 13252
rect 13587 13212 14556 13240
rect 13587 13209 13599 13212
rect 13541 13203 13599 13209
rect 14550 13200 14556 13212
rect 14608 13200 14614 13252
rect 14918 13200 14924 13252
rect 14976 13240 14982 13252
rect 16040 13249 16068 13280
rect 16025 13243 16083 13249
rect 16025 13240 16037 13243
rect 14976 13212 16037 13240
rect 14976 13200 14982 13212
rect 16025 13209 16037 13212
rect 16071 13209 16083 13243
rect 16408 13240 16436 13416
rect 17862 13404 17868 13456
rect 17920 13444 17926 13456
rect 20916 13444 20944 13484
rect 22554 13472 22560 13484
rect 22612 13472 22618 13524
rect 24578 13472 24584 13524
rect 24636 13512 24642 13524
rect 26970 13512 26976 13524
rect 24636 13484 26976 13512
rect 24636 13472 24642 13484
rect 21174 13444 21180 13456
rect 17920 13416 20944 13444
rect 21008 13416 21180 13444
rect 17920 13404 17926 13416
rect 16574 13336 16580 13388
rect 16632 13376 16638 13388
rect 17126 13376 17132 13388
rect 16632 13348 17132 13376
rect 16632 13336 16638 13348
rect 17126 13336 17132 13348
rect 17184 13336 17190 13388
rect 20162 13376 20168 13388
rect 19306 13348 20168 13376
rect 18046 13308 18052 13320
rect 17068 13280 18052 13308
rect 16853 13243 16911 13249
rect 16853 13240 16865 13243
rect 16408 13212 16865 13240
rect 16025 13203 16083 13209
rect 16853 13209 16865 13212
rect 16899 13209 16911 13243
rect 16853 13203 16911 13209
rect 8018 13132 8024 13184
rect 8076 13172 8082 13184
rect 8205 13175 8263 13181
rect 8205 13172 8217 13175
rect 8076 13144 8217 13172
rect 8076 13132 8082 13144
rect 8205 13141 8217 13144
rect 8251 13141 8263 13175
rect 9674 13172 9680 13184
rect 9635 13144 9680 13172
rect 8205 13135 8263 13141
rect 9674 13132 9680 13144
rect 9732 13132 9738 13184
rect 15470 13172 15476 13184
rect 15431 13144 15476 13172
rect 15470 13132 15476 13144
rect 15528 13132 15534 13184
rect 16225 13175 16283 13181
rect 16225 13141 16237 13175
rect 16271 13172 16283 13175
rect 16574 13172 16580 13184
rect 16271 13144 16580 13172
rect 16271 13141 16283 13144
rect 16225 13135 16283 13141
rect 16574 13132 16580 13144
rect 16632 13132 16638 13184
rect 16942 13132 16948 13184
rect 17000 13172 17006 13184
rect 17068 13181 17096 13280
rect 18046 13268 18052 13280
rect 18104 13268 18110 13320
rect 19306 13308 19334 13348
rect 20162 13336 20168 13348
rect 20220 13336 20226 13388
rect 19260 13280 19334 13308
rect 19260 13252 19288 13280
rect 19978 13268 19984 13320
rect 20036 13308 20042 13320
rect 20625 13311 20683 13317
rect 20036 13280 20208 13308
rect 20036 13268 20042 13280
rect 20180 13252 20208 13280
rect 20625 13277 20637 13311
rect 20671 13277 20683 13311
rect 20625 13271 20683 13277
rect 20773 13311 20831 13317
rect 20773 13277 20785 13311
rect 20819 13308 20831 13311
rect 21008 13308 21036 13416
rect 21174 13404 21180 13416
rect 21232 13404 21238 13456
rect 21634 13336 21640 13388
rect 21692 13376 21698 13388
rect 24872 13385 24900 13484
rect 26970 13472 26976 13484
rect 27028 13512 27034 13524
rect 27617 13515 27675 13521
rect 27617 13512 27629 13515
rect 27028 13484 27629 13512
rect 27028 13472 27034 13484
rect 27617 13481 27629 13484
rect 27663 13481 27675 13515
rect 27617 13475 27675 13481
rect 27430 13404 27436 13456
rect 27488 13444 27494 13456
rect 28258 13444 28264 13456
rect 27488 13416 28264 13444
rect 27488 13404 27494 13416
rect 28258 13404 28264 13416
rect 28316 13404 28322 13456
rect 24857 13379 24915 13385
rect 21692 13348 21956 13376
rect 21692 13336 21698 13348
rect 21174 13317 21180 13320
rect 20819 13280 21036 13308
rect 21131 13311 21180 13317
rect 20819 13277 20831 13280
rect 20773 13271 20831 13277
rect 21131 13277 21143 13311
rect 21177 13277 21180 13311
rect 21131 13271 21180 13277
rect 17954 13240 17960 13252
rect 17915 13212 17960 13240
rect 17954 13200 17960 13212
rect 18012 13200 18018 13252
rect 18138 13200 18144 13252
rect 18196 13249 18202 13252
rect 18196 13243 18215 13249
rect 18203 13209 18215 13243
rect 19242 13240 19248 13252
rect 19155 13212 19248 13240
rect 18196 13203 18215 13209
rect 18196 13200 18202 13203
rect 19242 13200 19248 13212
rect 19300 13200 19306 13252
rect 19334 13200 19340 13252
rect 19392 13240 19398 13252
rect 19461 13243 19519 13249
rect 19461 13240 19473 13243
rect 19392 13212 19473 13240
rect 19392 13200 19398 13212
rect 19461 13209 19473 13212
rect 19507 13240 19519 13243
rect 20070 13240 20076 13252
rect 19507 13212 20076 13240
rect 19507 13209 19519 13212
rect 19461 13203 19519 13209
rect 20070 13200 20076 13212
rect 20128 13200 20134 13252
rect 20162 13200 20168 13252
rect 20220 13200 20226 13252
rect 17053 13175 17111 13181
rect 17053 13172 17065 13175
rect 17000 13144 17065 13172
rect 17000 13132 17006 13144
rect 17053 13141 17065 13144
rect 17099 13141 17111 13175
rect 17053 13135 17111 13141
rect 17221 13175 17279 13181
rect 17221 13141 17233 13175
rect 17267 13172 17279 13175
rect 18046 13172 18052 13184
rect 17267 13144 18052 13172
rect 17267 13141 17279 13144
rect 17221 13135 17279 13141
rect 18046 13132 18052 13144
rect 18104 13132 18110 13184
rect 18325 13175 18383 13181
rect 18325 13141 18337 13175
rect 18371 13172 18383 13175
rect 20640 13172 20668 13271
rect 21174 13268 21180 13271
rect 21232 13268 21238 13320
rect 21726 13268 21732 13320
rect 21784 13308 21790 13320
rect 21928 13317 21956 13348
rect 22342 13348 23709 13376
rect 21821 13311 21879 13317
rect 21821 13308 21833 13311
rect 21784 13280 21833 13308
rect 21784 13268 21790 13280
rect 21821 13277 21833 13280
rect 21867 13277 21879 13311
rect 21821 13271 21879 13277
rect 21914 13311 21972 13317
rect 21914 13277 21926 13311
rect 21960 13277 21972 13311
rect 22186 13308 22192 13320
rect 22147 13280 22192 13308
rect 21914 13271 21972 13277
rect 22186 13268 22192 13280
rect 22244 13268 22250 13320
rect 22342 13317 22370 13348
rect 22327 13311 22385 13317
rect 22327 13277 22339 13311
rect 22373 13277 22385 13311
rect 22327 13271 22385 13277
rect 22554 13268 22560 13320
rect 22612 13308 22618 13320
rect 23201 13311 23259 13317
rect 23201 13308 23213 13311
rect 22612 13280 23213 13308
rect 22612 13268 22618 13280
rect 23201 13277 23213 13280
rect 23247 13277 23259 13311
rect 23201 13271 23259 13277
rect 23290 13268 23296 13320
rect 23348 13308 23354 13320
rect 23681 13317 23709 13348
rect 24857 13345 24869 13379
rect 24903 13345 24915 13379
rect 24857 13339 24915 13345
rect 27062 13336 27068 13388
rect 27120 13376 27126 13388
rect 27120 13348 28396 13376
rect 27120 13336 27126 13348
rect 23666 13311 23724 13317
rect 23348 13280 23393 13308
rect 23348 13268 23354 13280
rect 23666 13277 23678 13311
rect 23712 13308 23724 13311
rect 25124 13311 25182 13317
rect 23712 13280 25084 13308
rect 23712 13277 23724 13280
rect 23666 13271 23724 13277
rect 20901 13243 20959 13249
rect 20901 13209 20913 13243
rect 20947 13209 20959 13243
rect 20901 13203 20959 13209
rect 18371 13144 20668 13172
rect 20916 13172 20944 13203
rect 20990 13200 20996 13252
rect 21048 13240 21054 13252
rect 22097 13243 22155 13249
rect 22097 13240 22109 13243
rect 21048 13212 21093 13240
rect 21192 13212 22109 13240
rect 21048 13200 21054 13212
rect 21192 13172 21220 13212
rect 22097 13209 22109 13212
rect 22143 13240 22155 13243
rect 23477 13243 23535 13249
rect 22143 13212 22600 13240
rect 22143 13209 22155 13212
rect 22097 13203 22155 13209
rect 20916 13144 21220 13172
rect 21269 13175 21327 13181
rect 18371 13141 18383 13144
rect 18325 13135 18383 13141
rect 21269 13141 21281 13175
rect 21315 13172 21327 13175
rect 21450 13172 21456 13184
rect 21315 13144 21456 13172
rect 21315 13141 21327 13144
rect 21269 13135 21327 13141
rect 21450 13132 21456 13144
rect 21508 13132 21514 13184
rect 22002 13132 22008 13184
rect 22060 13172 22066 13184
rect 22465 13175 22523 13181
rect 22465 13172 22477 13175
rect 22060 13144 22477 13172
rect 22060 13132 22066 13144
rect 22465 13141 22477 13144
rect 22511 13141 22523 13175
rect 22572 13172 22600 13212
rect 23477 13209 23489 13243
rect 23523 13209 23535 13243
rect 23477 13203 23535 13209
rect 23569 13243 23627 13249
rect 23569 13209 23581 13243
rect 23615 13240 23627 13243
rect 24946 13240 24952 13252
rect 23615 13212 24952 13240
rect 23615 13209 23627 13212
rect 23569 13203 23627 13209
rect 23492 13172 23520 13203
rect 24946 13200 24952 13212
rect 25004 13200 25010 13252
rect 25056 13240 25084 13280
rect 25124 13277 25136 13311
rect 25170 13308 25182 13311
rect 26234 13308 26240 13320
rect 25170 13280 26240 13308
rect 25170 13277 25182 13280
rect 25124 13271 25182 13277
rect 26234 13268 26240 13280
rect 26292 13268 26298 13320
rect 26694 13268 26700 13320
rect 26752 13308 26758 13320
rect 26789 13311 26847 13317
rect 26789 13308 26801 13311
rect 26752 13280 26801 13308
rect 26752 13268 26758 13280
rect 26789 13277 26801 13280
rect 26835 13277 26847 13311
rect 26789 13271 26847 13277
rect 27614 13268 27620 13320
rect 27672 13268 27678 13320
rect 28368 13317 28396 13348
rect 28353 13311 28411 13317
rect 28353 13277 28365 13311
rect 28399 13277 28411 13311
rect 28353 13271 28411 13277
rect 25958 13240 25964 13252
rect 25056 13212 25964 13240
rect 25958 13200 25964 13212
rect 26016 13200 26022 13252
rect 26973 13243 27031 13249
rect 26973 13209 26985 13243
rect 27019 13240 27031 13243
rect 27525 13243 27583 13249
rect 27525 13240 27537 13243
rect 27019 13212 27537 13240
rect 27019 13209 27031 13212
rect 26973 13203 27031 13209
rect 27525 13209 27537 13212
rect 27571 13240 27583 13243
rect 27632 13240 27660 13268
rect 27571 13212 27660 13240
rect 27571 13209 27583 13212
rect 27525 13203 27583 13209
rect 23658 13172 23664 13184
rect 22572 13144 23664 13172
rect 22465 13135 22523 13141
rect 23658 13132 23664 13144
rect 23716 13132 23722 13184
rect 23845 13175 23903 13181
rect 23845 13141 23857 13175
rect 23891 13172 23903 13175
rect 24026 13172 24032 13184
rect 23891 13144 24032 13172
rect 23891 13141 23903 13144
rect 23845 13135 23903 13141
rect 24026 13132 24032 13144
rect 24084 13132 24090 13184
rect 25682 13132 25688 13184
rect 25740 13172 25746 13184
rect 26237 13175 26295 13181
rect 26237 13172 26249 13175
rect 25740 13144 26249 13172
rect 25740 13132 25746 13144
rect 26237 13141 26249 13144
rect 26283 13141 26295 13175
rect 26237 13135 26295 13141
rect 27246 13132 27252 13184
rect 27304 13172 27310 13184
rect 28169 13175 28227 13181
rect 28169 13172 28181 13175
rect 27304 13144 28181 13172
rect 27304 13132 27310 13144
rect 28169 13141 28181 13144
rect 28215 13141 28227 13175
rect 28169 13135 28227 13141
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 7837 12971 7895 12977
rect 7837 12937 7849 12971
rect 7883 12968 7895 12971
rect 9858 12968 9864 12980
rect 7883 12940 9674 12968
rect 9819 12940 9864 12968
rect 7883 12937 7895 12940
rect 7837 12931 7895 12937
rect 8294 12860 8300 12912
rect 8352 12900 8358 12912
rect 8662 12900 8668 12912
rect 8352 12872 8668 12900
rect 8352 12860 8358 12872
rect 8496 12841 8524 12872
rect 8662 12860 8668 12872
rect 8720 12900 8726 12912
rect 9398 12900 9404 12912
rect 8720 12872 9404 12900
rect 8720 12860 8726 12872
rect 9398 12860 9404 12872
rect 9456 12860 9462 12912
rect 9646 12900 9674 12940
rect 9858 12928 9864 12940
rect 9916 12928 9922 12980
rect 10502 12968 10508 12980
rect 10463 12940 10508 12968
rect 10502 12928 10508 12940
rect 10560 12928 10566 12980
rect 11606 12928 11612 12980
rect 11664 12968 11670 12980
rect 11885 12971 11943 12977
rect 11885 12968 11897 12971
rect 11664 12940 11897 12968
rect 11664 12928 11670 12940
rect 11885 12937 11897 12940
rect 11931 12937 11943 12971
rect 11885 12931 11943 12937
rect 13081 12971 13139 12977
rect 13081 12937 13093 12971
rect 13127 12968 13139 12971
rect 13170 12968 13176 12980
rect 13127 12940 13176 12968
rect 13127 12937 13139 12940
rect 13081 12931 13139 12937
rect 13170 12928 13176 12940
rect 13228 12928 13234 12980
rect 13906 12928 13912 12980
rect 13964 12968 13970 12980
rect 15949 12971 16007 12977
rect 15949 12968 15961 12971
rect 13964 12940 15961 12968
rect 13964 12928 13970 12940
rect 15949 12937 15961 12940
rect 15995 12937 16007 12971
rect 15949 12931 16007 12937
rect 16117 12971 16175 12977
rect 16117 12937 16129 12971
rect 16163 12968 16175 12971
rect 16163 12940 20944 12968
rect 16163 12937 16175 12940
rect 16117 12931 16175 12937
rect 11054 12900 11060 12912
rect 9646 12872 11060 12900
rect 11054 12860 11060 12872
rect 11112 12860 11118 12912
rect 11514 12900 11520 12912
rect 11475 12872 11520 12900
rect 11514 12860 11520 12872
rect 11572 12860 11578 12912
rect 11733 12903 11791 12909
rect 11733 12869 11745 12903
rect 11779 12900 11791 12903
rect 12434 12900 12440 12912
rect 11779 12872 12440 12900
rect 11779 12869 11791 12872
rect 11733 12863 11791 12869
rect 12434 12860 12440 12872
rect 12492 12860 12498 12912
rect 12618 12860 12624 12912
rect 12676 12900 12682 12912
rect 15746 12900 15752 12912
rect 12676 12872 14044 12900
rect 15707 12872 15752 12900
rect 12676 12860 12682 12872
rect 8021 12835 8079 12841
rect 8021 12801 8033 12835
rect 8067 12801 8079 12835
rect 8021 12795 8079 12801
rect 8481 12835 8539 12841
rect 8481 12801 8493 12835
rect 8527 12801 8539 12835
rect 8481 12795 8539 12801
rect 8748 12835 8806 12841
rect 8748 12801 8760 12835
rect 8794 12832 8806 12835
rect 9122 12832 9128 12844
rect 8794 12804 9128 12832
rect 8794 12801 8806 12804
rect 8748 12795 8806 12801
rect 8036 12628 8064 12795
rect 9122 12792 9128 12804
rect 9180 12792 9186 12844
rect 9306 12792 9312 12844
rect 9364 12832 9370 12844
rect 10686 12832 10692 12844
rect 9364 12804 10692 12832
rect 9364 12792 9370 12804
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 14016 12841 14044 12872
rect 15746 12860 15752 12872
rect 15804 12860 15810 12912
rect 15964 12900 15992 12931
rect 16942 12900 16948 12912
rect 15964 12872 16948 12900
rect 16942 12860 16948 12872
rect 17000 12860 17006 12912
rect 17218 12860 17224 12912
rect 17276 12900 17282 12912
rect 18601 12903 18659 12909
rect 18601 12900 18613 12903
rect 17276 12872 18613 12900
rect 17276 12860 17282 12872
rect 18601 12869 18613 12872
rect 18647 12869 18659 12903
rect 18601 12863 18659 12869
rect 18690 12860 18696 12912
rect 18748 12900 18754 12912
rect 20916 12900 20944 12940
rect 20990 12928 20996 12980
rect 21048 12968 21054 12980
rect 21269 12971 21327 12977
rect 21269 12968 21281 12971
rect 21048 12940 21281 12968
rect 21048 12928 21054 12940
rect 21269 12937 21281 12940
rect 21315 12937 21327 12971
rect 21269 12931 21327 12937
rect 23477 12971 23535 12977
rect 23477 12937 23489 12971
rect 23523 12968 23535 12971
rect 23566 12968 23572 12980
rect 23523 12940 23572 12968
rect 23523 12937 23535 12940
rect 23477 12931 23535 12937
rect 23566 12928 23572 12940
rect 23624 12928 23630 12980
rect 24118 12928 24124 12980
rect 24176 12968 24182 12980
rect 24305 12971 24363 12977
rect 24305 12968 24317 12971
rect 24176 12940 24317 12968
rect 24176 12928 24182 12940
rect 24305 12937 24317 12940
rect 24351 12937 24363 12971
rect 27430 12968 27436 12980
rect 24305 12931 24363 12937
rect 25516 12940 27436 12968
rect 21358 12900 21364 12912
rect 18748 12872 18793 12900
rect 19904 12872 20760 12900
rect 20916 12872 21364 12900
rect 18748 12860 18754 12872
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 14001 12835 14059 12841
rect 14001 12801 14013 12835
rect 14047 12832 14059 12835
rect 14274 12832 14280 12844
rect 14047 12804 14136 12832
rect 14235 12804 14280 12832
rect 14047 12801 14059 12804
rect 14001 12795 14059 12801
rect 13004 12764 13032 12795
rect 14108 12764 14136 12804
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 15470 12792 15476 12844
rect 15528 12832 15534 12844
rect 16669 12835 16727 12841
rect 16669 12832 16681 12835
rect 15528 12804 16681 12832
rect 15528 12792 15534 12804
rect 16669 12801 16681 12804
rect 16715 12832 16727 12835
rect 17678 12832 17684 12844
rect 16715 12804 17684 12832
rect 16715 12801 16727 12804
rect 16669 12795 16727 12801
rect 17678 12792 17684 12804
rect 17736 12792 17742 12844
rect 18230 12792 18236 12844
rect 18288 12832 18294 12844
rect 18506 12841 18512 12844
rect 18325 12835 18383 12841
rect 18325 12832 18337 12835
rect 18288 12804 18337 12832
rect 18288 12792 18294 12804
rect 18325 12801 18337 12804
rect 18371 12801 18383 12835
rect 18325 12795 18383 12801
rect 18473 12835 18512 12841
rect 18473 12801 18485 12835
rect 18473 12795 18512 12801
rect 18506 12792 18512 12795
rect 18564 12792 18570 12844
rect 18874 12841 18880 12844
rect 18831 12835 18880 12841
rect 18831 12801 18843 12835
rect 18877 12801 18880 12835
rect 18831 12795 18880 12801
rect 18874 12792 18880 12795
rect 18932 12792 18938 12844
rect 19904 12841 19932 12872
rect 20732 12844 20760 12872
rect 21358 12860 21364 12872
rect 21416 12860 21422 12912
rect 23293 12903 23351 12909
rect 23293 12900 23305 12903
rect 22066 12872 23305 12900
rect 19889 12835 19947 12841
rect 19889 12801 19901 12835
rect 19935 12801 19947 12835
rect 19889 12795 19947 12801
rect 20156 12835 20214 12841
rect 20156 12801 20168 12835
rect 20202 12832 20214 12835
rect 20438 12832 20444 12844
rect 20202 12804 20444 12832
rect 20202 12801 20214 12804
rect 20156 12795 20214 12801
rect 20438 12792 20444 12804
rect 20496 12792 20502 12844
rect 20714 12792 20720 12844
rect 20772 12832 20778 12844
rect 21910 12832 21916 12844
rect 20772 12804 21916 12832
rect 20772 12792 20778 12804
rect 21910 12792 21916 12804
rect 21968 12792 21974 12844
rect 22066 12776 22094 12872
rect 23293 12869 23305 12872
rect 23339 12869 23351 12903
rect 23293 12863 23351 12869
rect 23658 12860 23664 12912
rect 23716 12900 23722 12912
rect 23716 12872 24716 12900
rect 23716 12860 23722 12872
rect 22465 12835 22523 12841
rect 22465 12801 22477 12835
rect 22511 12832 22523 12835
rect 22646 12832 22652 12844
rect 22511 12804 22652 12832
rect 22511 12801 22523 12804
rect 22465 12795 22523 12801
rect 22646 12792 22652 12804
rect 22704 12792 22710 12844
rect 23109 12835 23167 12841
rect 23109 12801 23121 12835
rect 23155 12832 23167 12835
rect 23937 12835 23995 12841
rect 23937 12832 23949 12835
rect 23155 12804 23949 12832
rect 23155 12801 23167 12804
rect 23109 12795 23167 12801
rect 23937 12801 23949 12804
rect 23983 12801 23995 12835
rect 23937 12795 23995 12801
rect 16850 12764 16856 12776
rect 13004 12736 14044 12764
rect 14108 12736 16856 12764
rect 13906 12696 13912 12708
rect 9646 12668 13912 12696
rect 9646 12628 9674 12668
rect 13906 12656 13912 12668
rect 13964 12656 13970 12708
rect 14016 12696 14044 12736
rect 16850 12724 16856 12736
rect 16908 12724 16914 12776
rect 16945 12767 17003 12773
rect 16945 12733 16957 12767
rect 16991 12764 17003 12767
rect 17494 12764 17500 12776
rect 16991 12736 17500 12764
rect 16991 12733 17003 12736
rect 16945 12727 17003 12733
rect 17494 12724 17500 12736
rect 17552 12724 17558 12776
rect 20898 12724 20904 12776
rect 20956 12764 20962 12776
rect 21174 12764 21180 12776
rect 20956 12736 21180 12764
rect 20956 12724 20962 12736
rect 21174 12724 21180 12736
rect 21232 12724 21238 12776
rect 22002 12724 22008 12776
rect 22060 12736 22094 12776
rect 22281 12767 22339 12773
rect 22060 12724 22066 12736
rect 22281 12733 22293 12767
rect 22327 12764 22339 12767
rect 23014 12764 23020 12776
rect 22327 12736 23020 12764
rect 22327 12733 22339 12736
rect 22281 12727 22339 12733
rect 23014 12724 23020 12736
rect 23072 12724 23078 12776
rect 23952 12764 23980 12795
rect 24026 12792 24032 12844
rect 24084 12832 24090 12844
rect 24121 12835 24179 12841
rect 24121 12832 24133 12835
rect 24084 12804 24133 12832
rect 24084 12792 24090 12804
rect 24121 12801 24133 12804
rect 24167 12832 24179 12835
rect 24578 12832 24584 12844
rect 24167 12804 24584 12832
rect 24167 12801 24179 12804
rect 24121 12795 24179 12801
rect 24578 12792 24584 12804
rect 24636 12792 24642 12844
rect 24688 12764 24716 12872
rect 25314 12832 25320 12844
rect 25275 12804 25320 12832
rect 25314 12792 25320 12804
rect 25372 12792 25378 12844
rect 25516 12841 25544 12940
rect 27430 12928 27436 12940
rect 27488 12928 27494 12980
rect 27522 12928 27528 12980
rect 27580 12968 27586 12980
rect 28353 12971 28411 12977
rect 28353 12968 28365 12971
rect 27580 12940 28365 12968
rect 27580 12928 27586 12940
rect 28353 12937 28365 12940
rect 28399 12937 28411 12971
rect 28353 12931 28411 12937
rect 28813 12971 28871 12977
rect 28813 12937 28825 12971
rect 28859 12937 28871 12971
rect 28813 12931 28871 12937
rect 25682 12900 25688 12912
rect 25643 12872 25688 12900
rect 25682 12860 25688 12872
rect 25740 12860 25746 12912
rect 27240 12903 27298 12909
rect 27240 12869 27252 12903
rect 27286 12900 27298 12903
rect 28828 12900 28856 12931
rect 27286 12872 28856 12900
rect 27286 12869 27298 12872
rect 27240 12863 27298 12869
rect 25465 12835 25544 12841
rect 25465 12801 25477 12835
rect 25511 12804 25544 12835
rect 25593 12835 25651 12841
rect 25511 12801 25523 12804
rect 25465 12795 25523 12801
rect 25593 12801 25605 12835
rect 25639 12801 25651 12835
rect 25593 12795 25651 12801
rect 25782 12835 25840 12841
rect 25782 12801 25794 12835
rect 25828 12832 25840 12835
rect 25958 12832 25964 12844
rect 25828 12804 25964 12832
rect 25828 12801 25840 12804
rect 25782 12795 25840 12801
rect 25608 12764 25636 12795
rect 25958 12792 25964 12804
rect 26016 12792 26022 12844
rect 26970 12832 26976 12844
rect 26931 12804 26976 12832
rect 26970 12792 26976 12804
rect 27028 12792 27034 12844
rect 27706 12792 27712 12844
rect 27764 12832 27770 12844
rect 28997 12835 29055 12841
rect 28997 12832 29009 12835
rect 27764 12804 29009 12832
rect 27764 12792 27770 12804
rect 28997 12801 29009 12804
rect 29043 12801 29055 12835
rect 28997 12795 29055 12801
rect 23952 12736 24164 12764
rect 24688 12736 25636 12764
rect 24136 12708 24164 12736
rect 19058 12696 19064 12708
rect 14016 12668 19064 12696
rect 19058 12656 19064 12668
rect 19116 12656 19122 12708
rect 24118 12656 24124 12708
rect 24176 12656 24182 12708
rect 25608 12696 25636 12736
rect 25866 12724 25872 12776
rect 25924 12724 25930 12776
rect 25884 12696 25912 12724
rect 25608 12668 25912 12696
rect 11698 12628 11704 12640
rect 8036 12600 9674 12628
rect 11659 12600 11704 12628
rect 11698 12588 11704 12600
rect 11756 12588 11762 12640
rect 13446 12588 13452 12640
rect 13504 12628 13510 12640
rect 14366 12628 14372 12640
rect 13504 12600 14372 12628
rect 13504 12588 13510 12600
rect 14366 12588 14372 12600
rect 14424 12628 14430 12640
rect 15654 12628 15660 12640
rect 14424 12600 15660 12628
rect 14424 12588 14430 12600
rect 15654 12588 15660 12600
rect 15712 12588 15718 12640
rect 15933 12631 15991 12637
rect 15933 12597 15945 12631
rect 15979 12628 15991 12631
rect 17034 12628 17040 12640
rect 15979 12600 17040 12628
rect 15979 12597 15991 12600
rect 15933 12591 15991 12597
rect 17034 12588 17040 12600
rect 17092 12588 17098 12640
rect 18969 12631 19027 12637
rect 18969 12597 18981 12631
rect 19015 12628 19027 12631
rect 20622 12628 20628 12640
rect 19015 12600 20628 12628
rect 19015 12597 19027 12600
rect 18969 12591 19027 12597
rect 20622 12588 20628 12600
rect 20680 12588 20686 12640
rect 22370 12588 22376 12640
rect 22428 12628 22434 12640
rect 22649 12631 22707 12637
rect 22649 12628 22661 12631
rect 22428 12600 22661 12628
rect 22428 12588 22434 12600
rect 22649 12597 22661 12600
rect 22695 12597 22707 12631
rect 22649 12591 22707 12597
rect 25866 12588 25872 12640
rect 25924 12628 25930 12640
rect 25961 12631 26019 12637
rect 25961 12628 25973 12631
rect 25924 12600 25973 12628
rect 25924 12588 25930 12600
rect 25961 12597 25973 12600
rect 26007 12597 26019 12631
rect 25961 12591 26019 12597
rect 26786 12588 26792 12640
rect 26844 12628 26850 12640
rect 26970 12628 26976 12640
rect 26844 12600 26976 12628
rect 26844 12588 26850 12600
rect 26970 12588 26976 12600
rect 27028 12588 27034 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 5994 12384 6000 12436
rect 6052 12424 6058 12436
rect 8846 12424 8852 12436
rect 6052 12396 8852 12424
rect 6052 12384 6058 12396
rect 8846 12384 8852 12396
rect 8904 12384 8910 12436
rect 9122 12424 9128 12436
rect 9083 12396 9128 12424
rect 9122 12384 9128 12396
rect 9180 12384 9186 12436
rect 11698 12384 11704 12436
rect 11756 12424 11762 12436
rect 11793 12427 11851 12433
rect 11793 12424 11805 12427
rect 11756 12396 11805 12424
rect 11756 12384 11762 12396
rect 11793 12393 11805 12396
rect 11839 12393 11851 12427
rect 13446 12424 13452 12436
rect 13407 12396 13452 12424
rect 11793 12387 11851 12393
rect 13446 12384 13452 12396
rect 13504 12384 13510 12436
rect 14369 12427 14427 12433
rect 14369 12424 14381 12427
rect 13648 12396 14381 12424
rect 7561 12359 7619 12365
rect 7561 12325 7573 12359
rect 7607 12356 7619 12359
rect 10134 12356 10140 12368
rect 7607 12328 10140 12356
rect 7607 12325 7619 12328
rect 7561 12319 7619 12325
rect 10134 12316 10140 12328
rect 10192 12316 10198 12368
rect 10226 12288 10232 12300
rect 7760 12260 10232 12288
rect 7760 12229 7788 12260
rect 10226 12248 10232 12260
rect 10284 12248 10290 12300
rect 13078 12248 13084 12300
rect 13136 12288 13142 12300
rect 13357 12291 13415 12297
rect 13357 12288 13369 12291
rect 13136 12260 13369 12288
rect 13136 12248 13142 12260
rect 13357 12257 13369 12260
rect 13403 12288 13415 12291
rect 13648 12288 13676 12396
rect 14369 12393 14381 12396
rect 14415 12393 14427 12427
rect 14369 12387 14427 12393
rect 14737 12427 14795 12433
rect 14737 12393 14749 12427
rect 14783 12424 14795 12427
rect 15010 12424 15016 12436
rect 14783 12396 15016 12424
rect 14783 12393 14795 12396
rect 14737 12387 14795 12393
rect 15010 12384 15016 12396
rect 15068 12384 15074 12436
rect 15286 12384 15292 12436
rect 15344 12424 15350 12436
rect 15749 12427 15807 12433
rect 15749 12424 15761 12427
rect 15344 12396 15761 12424
rect 15344 12384 15350 12396
rect 15749 12393 15761 12396
rect 15795 12424 15807 12427
rect 16482 12424 16488 12436
rect 15795 12396 16488 12424
rect 15795 12393 15807 12396
rect 15749 12387 15807 12393
rect 16482 12384 16488 12396
rect 16540 12384 16546 12436
rect 18230 12384 18236 12436
rect 18288 12424 18294 12436
rect 20898 12424 20904 12436
rect 18288 12396 20904 12424
rect 18288 12384 18294 12396
rect 20898 12384 20904 12396
rect 20956 12384 20962 12436
rect 21082 12384 21088 12436
rect 21140 12424 21146 12436
rect 21269 12427 21327 12433
rect 21269 12424 21281 12427
rect 21140 12396 21281 12424
rect 21140 12384 21146 12396
rect 21269 12393 21281 12396
rect 21315 12393 21327 12427
rect 21269 12387 21327 12393
rect 21453 12427 21511 12433
rect 21453 12393 21465 12427
rect 21499 12424 21511 12427
rect 21542 12424 21548 12436
rect 21499 12396 21548 12424
rect 21499 12393 21511 12396
rect 21453 12387 21511 12393
rect 21542 12384 21548 12396
rect 21600 12384 21606 12436
rect 23658 12384 23664 12436
rect 23716 12424 23722 12436
rect 23753 12427 23811 12433
rect 23753 12424 23765 12427
rect 23716 12396 23765 12424
rect 23716 12384 23722 12396
rect 23753 12393 23765 12396
rect 23799 12393 23811 12427
rect 23753 12387 23811 12393
rect 25593 12427 25651 12433
rect 25593 12393 25605 12427
rect 25639 12424 25651 12427
rect 25774 12424 25780 12436
rect 25639 12396 25780 12424
rect 25639 12393 25651 12396
rect 25593 12387 25651 12393
rect 25774 12384 25780 12396
rect 25832 12384 25838 12436
rect 26142 12384 26148 12436
rect 26200 12424 26206 12436
rect 28537 12427 28595 12433
rect 28537 12424 28549 12427
rect 26200 12396 28549 12424
rect 26200 12384 26206 12396
rect 28537 12393 28549 12396
rect 28583 12393 28595 12427
rect 28537 12387 28595 12393
rect 13722 12316 13728 12368
rect 13780 12356 13786 12368
rect 14231 12359 14289 12365
rect 14231 12356 14243 12359
rect 13780 12328 14243 12356
rect 13780 12316 13786 12328
rect 14231 12325 14243 12328
rect 14277 12325 14289 12359
rect 14231 12319 14289 12325
rect 14550 12316 14556 12368
rect 14608 12356 14614 12368
rect 21634 12356 21640 12368
rect 14608 12328 21640 12356
rect 14608 12316 14614 12328
rect 21634 12316 21640 12328
rect 21692 12316 21698 12368
rect 22649 12359 22707 12365
rect 22649 12356 22661 12359
rect 21744 12328 22661 12356
rect 13403 12260 13676 12288
rect 13403 12257 13415 12260
rect 13357 12251 13415 12257
rect 13814 12248 13820 12300
rect 13872 12288 13878 12300
rect 14461 12291 14519 12297
rect 14461 12288 14473 12291
rect 13872 12260 14473 12288
rect 13872 12248 13878 12260
rect 14461 12257 14473 12260
rect 14507 12257 14519 12291
rect 15654 12288 15660 12300
rect 15567 12260 15660 12288
rect 14461 12251 14519 12257
rect 15654 12248 15660 12260
rect 15712 12288 15718 12300
rect 16022 12288 16028 12300
rect 15712 12260 16028 12288
rect 15712 12248 15718 12260
rect 16022 12248 16028 12260
rect 16080 12248 16086 12300
rect 16853 12291 16911 12297
rect 16853 12257 16865 12291
rect 16899 12288 16911 12291
rect 16942 12288 16948 12300
rect 16899 12260 16948 12288
rect 16899 12257 16911 12260
rect 16853 12251 16911 12257
rect 16942 12248 16948 12260
rect 17000 12248 17006 12300
rect 17126 12288 17132 12300
rect 17087 12260 17132 12288
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 19797 12291 19855 12297
rect 19797 12257 19809 12291
rect 19843 12288 19855 12291
rect 20346 12288 20352 12300
rect 19843 12260 20352 12288
rect 19843 12257 19855 12260
rect 19797 12251 19855 12257
rect 20346 12248 20352 12260
rect 20404 12248 20410 12300
rect 20438 12248 20444 12300
rect 20496 12288 20502 12300
rect 21744 12288 21772 12328
rect 22649 12325 22661 12328
rect 22695 12325 22707 12359
rect 22649 12319 22707 12325
rect 24302 12316 24308 12368
rect 24360 12356 24366 12368
rect 28074 12356 28080 12368
rect 24360 12328 28080 12356
rect 24360 12316 24366 12328
rect 28074 12316 28080 12328
rect 28132 12316 28138 12368
rect 20496 12260 21772 12288
rect 20496 12248 20502 12260
rect 22094 12248 22100 12300
rect 22152 12288 22158 12300
rect 22152 12260 22508 12288
rect 22152 12248 22158 12260
rect 7745 12223 7803 12229
rect 7745 12189 7757 12223
rect 7791 12189 7803 12223
rect 7745 12183 7803 12189
rect 8389 12223 8447 12229
rect 8389 12189 8401 12223
rect 8435 12189 8447 12223
rect 8389 12183 8447 12189
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12220 9367 12223
rect 9674 12220 9680 12232
rect 9355 12192 9680 12220
rect 9355 12189 9367 12192
rect 9309 12183 9367 12189
rect 8404 12152 8432 12183
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 9950 12220 9956 12232
rect 9911 12192 9956 12220
rect 9950 12180 9956 12192
rect 10008 12180 10014 12232
rect 10410 12220 10416 12232
rect 10371 12192 10416 12220
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 10686 12229 10692 12232
rect 10680 12183 10692 12229
rect 10744 12220 10750 12232
rect 10744 12192 10780 12220
rect 10686 12180 10692 12183
rect 10744 12180 10750 12192
rect 10962 12180 10968 12232
rect 11020 12220 11026 12232
rect 12529 12223 12587 12229
rect 12529 12220 12541 12223
rect 11020 12192 12541 12220
rect 11020 12180 11026 12192
rect 12529 12189 12541 12192
rect 12575 12189 12587 12223
rect 12529 12183 12587 12189
rect 12802 12180 12808 12232
rect 12860 12220 12866 12232
rect 13265 12223 13323 12229
rect 13265 12220 13277 12223
rect 12860 12192 13277 12220
rect 12860 12180 12866 12192
rect 13265 12189 13277 12192
rect 13311 12189 13323 12223
rect 15470 12220 15476 12232
rect 15431 12192 15476 12220
rect 13265 12183 13323 12189
rect 15470 12180 15476 12192
rect 15528 12180 15534 12232
rect 15838 12220 15844 12232
rect 15799 12192 15844 12220
rect 15838 12180 15844 12192
rect 15896 12180 15902 12232
rect 17494 12180 17500 12232
rect 17552 12220 17558 12232
rect 18509 12223 18567 12229
rect 18509 12220 18521 12223
rect 17552 12192 18521 12220
rect 17552 12180 17558 12192
rect 18509 12189 18521 12192
rect 18555 12189 18567 12223
rect 18509 12183 18567 12189
rect 19978 12180 19984 12232
rect 20036 12220 20042 12232
rect 20073 12223 20131 12229
rect 20073 12220 20085 12223
rect 20036 12192 20085 12220
rect 20036 12180 20042 12192
rect 20073 12189 20085 12192
rect 20119 12220 20131 12223
rect 22370 12220 22376 12232
rect 20119 12216 20944 12220
rect 20119 12192 21036 12216
rect 22331 12192 22376 12220
rect 20119 12189 20131 12192
rect 20073 12183 20131 12189
rect 20916 12188 21036 12192
rect 10318 12152 10324 12164
rect 8404 12124 10324 12152
rect 10318 12112 10324 12124
rect 10376 12112 10382 12164
rect 12345 12155 12403 12161
rect 12345 12121 12357 12155
rect 12391 12152 12403 12155
rect 12434 12152 12440 12164
rect 12391 12124 12440 12152
rect 12391 12121 12403 12124
rect 12345 12115 12403 12121
rect 12434 12112 12440 12124
rect 12492 12152 12498 12164
rect 12986 12152 12992 12164
rect 12492 12124 12992 12152
rect 12492 12112 12498 12124
rect 12986 12112 12992 12124
rect 13044 12112 13050 12164
rect 13541 12155 13599 12161
rect 13541 12121 13553 12155
rect 13587 12121 13599 12155
rect 13541 12115 13599 12121
rect 14093 12155 14151 12161
rect 14093 12121 14105 12155
rect 14139 12152 14151 12155
rect 14182 12152 14188 12164
rect 14139 12124 14188 12152
rect 14139 12121 14151 12124
rect 14093 12115 14151 12121
rect 8205 12087 8263 12093
rect 8205 12053 8217 12087
rect 8251 12084 8263 12087
rect 8938 12084 8944 12096
rect 8251 12056 8944 12084
rect 8251 12053 8263 12056
rect 8205 12047 8263 12053
rect 8938 12044 8944 12056
rect 8996 12044 9002 12096
rect 9766 12084 9772 12096
rect 9727 12056 9772 12084
rect 9766 12044 9772 12056
rect 9824 12044 9830 12096
rect 12526 12044 12532 12096
rect 12584 12084 12590 12096
rect 13556 12084 13584 12115
rect 14182 12112 14188 12124
rect 14240 12112 14246 12164
rect 18693 12155 18751 12161
rect 18693 12121 18705 12155
rect 18739 12152 18751 12155
rect 18966 12152 18972 12164
rect 18739 12124 18972 12152
rect 18739 12121 18751 12124
rect 18693 12115 18751 12121
rect 18966 12112 18972 12124
rect 19024 12152 19030 12164
rect 20438 12152 20444 12164
rect 19024 12124 20444 12152
rect 19024 12112 19030 12124
rect 20438 12112 20444 12124
rect 20496 12112 20502 12164
rect 21008 12152 21036 12188
rect 22370 12180 22376 12192
rect 22428 12180 22434 12232
rect 22480 12229 22508 12260
rect 23658 12248 23664 12300
rect 23716 12288 23722 12300
rect 24210 12288 24216 12300
rect 23716 12260 24216 12288
rect 23716 12248 23722 12260
rect 24210 12248 24216 12260
rect 24268 12248 24274 12300
rect 25406 12288 25412 12300
rect 24596 12260 25412 12288
rect 22465 12223 22523 12229
rect 22465 12189 22477 12223
rect 22511 12189 22523 12223
rect 22465 12183 22523 12189
rect 22741 12223 22799 12229
rect 22741 12189 22753 12223
rect 22787 12220 22799 12223
rect 23290 12220 23296 12232
rect 22787 12192 23296 12220
rect 22787 12189 22799 12192
rect 22741 12183 22799 12189
rect 23290 12180 23296 12192
rect 23348 12180 23354 12232
rect 21111 12155 21169 12161
rect 21111 12152 21123 12155
rect 21008 12124 21123 12152
rect 21111 12121 21123 12124
rect 21157 12121 21169 12155
rect 21111 12115 21169 12121
rect 23106 12112 23112 12164
rect 23164 12152 23170 12164
rect 23661 12155 23719 12161
rect 23661 12152 23673 12155
rect 23164 12124 23673 12152
rect 23164 12112 23170 12124
rect 23661 12121 23673 12124
rect 23707 12121 23719 12155
rect 23661 12115 23719 12121
rect 24210 12112 24216 12164
rect 24268 12152 24274 12164
rect 24596 12161 24624 12260
rect 25406 12248 25412 12260
rect 25464 12248 25470 12300
rect 25958 12248 25964 12300
rect 26016 12288 26022 12300
rect 26973 12291 27031 12297
rect 26973 12288 26985 12291
rect 26016 12260 26985 12288
rect 26016 12248 26022 12260
rect 26973 12257 26985 12260
rect 27019 12288 27031 12291
rect 27019 12260 28396 12288
rect 27019 12257 27031 12260
rect 26973 12251 27031 12257
rect 24765 12223 24823 12229
rect 24765 12189 24777 12223
rect 24811 12220 24823 12223
rect 24811 12192 26188 12220
rect 24811 12189 24823 12192
rect 24765 12183 24823 12189
rect 24397 12155 24455 12161
rect 24397 12152 24409 12155
rect 24268 12124 24409 12152
rect 24268 12112 24274 12124
rect 24397 12121 24409 12124
rect 24443 12121 24455 12155
rect 24397 12115 24455 12121
rect 24581 12155 24639 12161
rect 24581 12121 24593 12155
rect 24627 12121 24639 12155
rect 25225 12155 25283 12161
rect 25225 12152 25237 12155
rect 24581 12115 24639 12121
rect 24688 12124 25237 12152
rect 13814 12084 13820 12096
rect 12584 12056 13820 12084
rect 12584 12044 12590 12056
rect 13814 12044 13820 12056
rect 13872 12044 13878 12096
rect 19334 12044 19340 12096
rect 19392 12084 19398 12096
rect 20254 12084 20260 12096
rect 19392 12056 20260 12084
rect 19392 12044 19398 12056
rect 20254 12044 20260 12056
rect 20312 12044 20318 12096
rect 20806 12044 20812 12096
rect 20864 12084 20870 12096
rect 21285 12087 21343 12093
rect 21285 12084 21297 12087
rect 20864 12056 21297 12084
rect 20864 12044 20870 12056
rect 21285 12053 21297 12056
rect 21331 12084 21343 12087
rect 21450 12084 21456 12096
rect 21331 12056 21456 12084
rect 21331 12053 21343 12056
rect 21285 12047 21343 12053
rect 21450 12044 21456 12056
rect 21508 12044 21514 12096
rect 22189 12087 22247 12093
rect 22189 12053 22201 12087
rect 22235 12084 22247 12087
rect 22646 12084 22652 12096
rect 22235 12056 22652 12084
rect 22235 12053 22247 12056
rect 22189 12047 22247 12053
rect 22646 12044 22652 12056
rect 22704 12044 22710 12096
rect 24412 12084 24440 12115
rect 24688 12084 24716 12124
rect 25225 12121 25237 12124
rect 25271 12121 25283 12155
rect 25225 12115 25283 12121
rect 25409 12155 25467 12161
rect 25409 12121 25421 12155
rect 25455 12152 25467 12155
rect 25682 12152 25688 12164
rect 25455 12124 25688 12152
rect 25455 12121 25467 12124
rect 25409 12115 25467 12121
rect 25682 12112 25688 12124
rect 25740 12152 25746 12164
rect 25866 12152 25872 12164
rect 25740 12124 25872 12152
rect 25740 12112 25746 12124
rect 25866 12112 25872 12124
rect 25924 12112 25930 12164
rect 26160 12152 26188 12192
rect 26234 12180 26240 12232
rect 26292 12220 26298 12232
rect 26697 12223 26755 12229
rect 26292 12192 26337 12220
rect 26292 12180 26298 12192
rect 26697 12189 26709 12223
rect 26743 12220 26755 12223
rect 27430 12220 27436 12232
rect 26743 12192 27436 12220
rect 26743 12189 26755 12192
rect 26697 12183 26755 12189
rect 27430 12180 27436 12192
rect 27488 12180 27494 12232
rect 27982 12220 27988 12232
rect 27943 12192 27988 12220
rect 27982 12180 27988 12192
rect 28040 12180 28046 12232
rect 28368 12229 28396 12260
rect 28353 12223 28411 12229
rect 28353 12189 28365 12223
rect 28399 12189 28411 12223
rect 28353 12183 28411 12189
rect 26160 12124 28028 12152
rect 24412 12056 24716 12084
rect 24854 12044 24860 12096
rect 24912 12084 24918 12096
rect 26053 12087 26111 12093
rect 26053 12084 26065 12087
rect 24912 12056 26065 12084
rect 24912 12044 24918 12056
rect 26053 12053 26065 12056
rect 26099 12053 26111 12087
rect 26053 12047 26111 12053
rect 27154 12044 27160 12096
rect 27212 12084 27218 12096
rect 27522 12084 27528 12096
rect 27212 12056 27528 12084
rect 27212 12044 27218 12056
rect 27522 12044 27528 12056
rect 27580 12044 27586 12096
rect 28000 12084 28028 12124
rect 28074 12112 28080 12164
rect 28132 12152 28138 12164
rect 28169 12155 28227 12161
rect 28169 12152 28181 12155
rect 28132 12124 28181 12152
rect 28132 12112 28138 12124
rect 28169 12121 28181 12124
rect 28215 12121 28227 12155
rect 28169 12115 28227 12121
rect 28258 12112 28264 12164
rect 28316 12152 28322 12164
rect 28316 12124 28361 12152
rect 28316 12112 28322 12124
rect 28442 12084 28448 12096
rect 28000 12056 28448 12084
rect 28442 12044 28448 12056
rect 28500 12044 28506 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 5902 11840 5908 11892
rect 5960 11880 5966 11892
rect 10778 11880 10784 11892
rect 5960 11852 10640 11880
rect 10739 11852 10784 11880
rect 5960 11840 5966 11852
rect 8754 11812 8760 11824
rect 6380 11784 8760 11812
rect 6380 11753 6408 11784
rect 8754 11772 8760 11784
rect 8812 11772 8818 11824
rect 10612 11812 10640 11852
rect 10778 11840 10784 11852
rect 10836 11840 10842 11892
rect 10870 11840 10876 11892
rect 10928 11880 10934 11892
rect 11517 11883 11575 11889
rect 11517 11880 11529 11883
rect 10928 11852 11529 11880
rect 10928 11840 10934 11852
rect 11517 11849 11529 11852
rect 11563 11849 11575 11883
rect 11517 11843 11575 11849
rect 12437 11883 12495 11889
rect 12437 11849 12449 11883
rect 12483 11880 12495 11883
rect 12526 11880 12532 11892
rect 12483 11852 12532 11880
rect 12483 11849 12495 11852
rect 12437 11843 12495 11849
rect 12526 11840 12532 11852
rect 12584 11840 12590 11892
rect 15013 11883 15071 11889
rect 12636 11852 14504 11880
rect 12161 11815 12219 11821
rect 12161 11812 12173 11815
rect 10612 11784 12173 11812
rect 12161 11781 12173 11784
rect 12207 11812 12219 11815
rect 12250 11812 12256 11824
rect 12207 11784 12256 11812
rect 12207 11781 12219 11784
rect 12161 11775 12219 11781
rect 12250 11772 12256 11784
rect 12308 11772 12314 11824
rect 12342 11772 12348 11824
rect 12400 11812 12406 11824
rect 12636 11812 12664 11852
rect 14476 11824 14504 11852
rect 15013 11849 15025 11883
rect 15059 11880 15071 11883
rect 15378 11880 15384 11892
rect 15059 11852 15384 11880
rect 15059 11849 15071 11852
rect 15013 11843 15071 11849
rect 15378 11840 15384 11852
rect 15436 11840 15442 11892
rect 15930 11840 15936 11892
rect 15988 11880 15994 11892
rect 15988 11852 18460 11880
rect 15988 11840 15994 11852
rect 13722 11812 13728 11824
rect 12400 11784 12445 11812
rect 12544 11784 12664 11812
rect 12912 11784 13728 11812
rect 12400 11772 12406 11784
rect 6365 11747 6423 11753
rect 6365 11713 6377 11747
rect 6411 11713 6423 11747
rect 6365 11707 6423 11713
rect 6454 11704 6460 11756
rect 6512 11744 6518 11756
rect 6621 11747 6679 11753
rect 6621 11744 6633 11747
rect 6512 11716 6633 11744
rect 6512 11704 6518 11716
rect 6621 11713 6633 11716
rect 6667 11713 6679 11747
rect 6621 11707 6679 11713
rect 8564 11747 8622 11753
rect 8564 11713 8576 11747
rect 8610 11744 8622 11747
rect 9766 11744 9772 11756
rect 8610 11716 9772 11744
rect 8610 11713 8622 11716
rect 8564 11707 8622 11713
rect 9766 11704 9772 11716
rect 9824 11704 9830 11756
rect 10965 11747 11023 11753
rect 10965 11713 10977 11747
rect 11011 11744 11023 11747
rect 11422 11744 11428 11756
rect 11011 11716 11428 11744
rect 11011 11713 11023 11716
rect 10965 11707 11023 11713
rect 11422 11704 11428 11716
rect 11480 11704 11486 11756
rect 11701 11747 11759 11753
rect 11701 11713 11713 11747
rect 11747 11744 11759 11747
rect 11882 11744 11888 11756
rect 11747 11716 11888 11744
rect 11747 11713 11759 11716
rect 11701 11707 11759 11713
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 12437 11747 12495 11753
rect 12437 11713 12449 11747
rect 12483 11746 12495 11747
rect 12483 11744 12496 11746
rect 12544 11744 12572 11784
rect 12483 11716 12572 11744
rect 12483 11713 12495 11716
rect 12437 11707 12495 11713
rect 8297 11679 8355 11685
rect 8297 11645 8309 11679
rect 8343 11645 8355 11679
rect 8297 11639 8355 11645
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 7524 11512 7757 11540
rect 7524 11500 7530 11512
rect 7745 11509 7757 11512
rect 7791 11509 7803 11543
rect 8312 11540 8340 11639
rect 10410 11608 10416 11620
rect 9232 11580 10416 11608
rect 9232 11540 9260 11580
rect 10410 11568 10416 11580
rect 10468 11568 10474 11620
rect 12544 11608 12572 11716
rect 12802 11704 12808 11756
rect 12860 11744 12866 11756
rect 12912 11753 12940 11784
rect 13722 11772 13728 11784
rect 13780 11812 13786 11824
rect 13817 11815 13875 11821
rect 13817 11812 13829 11815
rect 13780 11784 13829 11812
rect 13780 11772 13786 11784
rect 13817 11781 13829 11784
rect 13863 11781 13875 11815
rect 13817 11775 13875 11781
rect 14458 11772 14464 11824
rect 14516 11812 14522 11824
rect 16025 11815 16083 11821
rect 14516 11784 15976 11812
rect 14516 11772 14522 11784
rect 12897 11747 12955 11753
rect 12897 11744 12909 11747
rect 12860 11716 12909 11744
rect 12860 11704 12866 11716
rect 12897 11713 12909 11716
rect 12943 11713 12955 11747
rect 13078 11744 13084 11756
rect 13039 11716 13084 11744
rect 12897 11707 12955 11713
rect 13078 11704 13084 11716
rect 13136 11744 13142 11756
rect 14001 11747 14059 11753
rect 14001 11744 14013 11747
rect 13136 11716 14013 11744
rect 13136 11704 13142 11716
rect 14001 11713 14013 11716
rect 14047 11713 14059 11747
rect 14001 11707 14059 11713
rect 14093 11747 14151 11753
rect 14093 11713 14105 11747
rect 14139 11744 14151 11747
rect 14826 11744 14832 11756
rect 14139 11716 14832 11744
rect 14139 11713 14151 11716
rect 14093 11707 14151 11713
rect 14826 11704 14832 11716
rect 14884 11704 14890 11756
rect 15197 11747 15255 11753
rect 15197 11713 15209 11747
rect 15243 11713 15255 11747
rect 15197 11707 15255 11713
rect 15473 11747 15531 11753
rect 15473 11713 15485 11747
rect 15519 11744 15531 11747
rect 15654 11744 15660 11756
rect 15519 11716 15660 11744
rect 15519 11713 15531 11716
rect 15473 11707 15531 11713
rect 15212 11676 15240 11707
rect 15654 11704 15660 11716
rect 15712 11704 15718 11756
rect 15948 11753 15976 11784
rect 16025 11781 16037 11815
rect 16071 11812 16083 11815
rect 16574 11812 16580 11824
rect 16071 11784 16580 11812
rect 16071 11781 16083 11784
rect 16025 11775 16083 11781
rect 16574 11772 16580 11784
rect 16632 11812 16638 11824
rect 17037 11815 17095 11821
rect 17037 11812 17049 11815
rect 16632 11784 17049 11812
rect 16632 11772 16638 11784
rect 17037 11781 17049 11784
rect 17083 11781 17095 11815
rect 18432 11812 18460 11852
rect 18506 11840 18512 11892
rect 18564 11880 18570 11892
rect 19245 11883 19303 11889
rect 19245 11880 19257 11883
rect 18564 11852 19257 11880
rect 18564 11840 18570 11852
rect 19245 11849 19257 11852
rect 19291 11880 19303 11883
rect 22922 11880 22928 11892
rect 19291 11852 19840 11880
rect 19291 11849 19303 11852
rect 19245 11843 19303 11849
rect 19518 11812 19524 11824
rect 18432 11784 19524 11812
rect 17037 11775 17095 11781
rect 19518 11772 19524 11784
rect 19576 11812 19582 11824
rect 19576 11784 19748 11812
rect 19576 11772 19582 11784
rect 15933 11747 15991 11753
rect 15933 11713 15945 11747
rect 15979 11713 15991 11747
rect 16850 11744 16856 11756
rect 16811 11716 16856 11744
rect 15933 11707 15991 11713
rect 16850 11704 16856 11716
rect 16908 11704 16914 11756
rect 19720 11753 19748 11784
rect 17129 11747 17187 11753
rect 17129 11713 17141 11747
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 17865 11747 17923 11753
rect 17865 11713 17877 11747
rect 17911 11713 17923 11747
rect 17865 11707 17923 11713
rect 18132 11747 18190 11753
rect 18132 11713 18144 11747
rect 18178 11744 18190 11747
rect 19705 11747 19763 11753
rect 18178 11716 19288 11744
rect 18178 11713 18190 11716
rect 18132 11707 18190 11713
rect 15212 11648 15700 11676
rect 15672 11620 15700 11648
rect 12360 11580 12572 11608
rect 14277 11611 14335 11617
rect 8312 11512 9260 11540
rect 7745 11503 7803 11509
rect 9582 11500 9588 11552
rect 9640 11540 9646 11552
rect 9677 11543 9735 11549
rect 9677 11540 9689 11543
rect 9640 11512 9689 11540
rect 9640 11500 9646 11512
rect 9677 11509 9689 11512
rect 9723 11540 9735 11543
rect 12360 11540 12388 11580
rect 14277 11577 14289 11611
rect 14323 11608 14335 11611
rect 15381 11611 15439 11617
rect 15381 11608 15393 11611
rect 14323 11580 15393 11608
rect 14323 11577 14335 11580
rect 14277 11571 14335 11577
rect 15381 11577 15393 11580
rect 15427 11608 15439 11611
rect 15470 11608 15476 11620
rect 15427 11580 15476 11608
rect 15427 11577 15439 11580
rect 15381 11571 15439 11577
rect 15470 11568 15476 11580
rect 15528 11568 15534 11620
rect 15654 11568 15660 11620
rect 15712 11568 15718 11620
rect 17144 11608 17172 11707
rect 15764 11580 17172 11608
rect 9723 11512 12388 11540
rect 9723 11509 9735 11512
rect 9677 11503 9735 11509
rect 12894 11500 12900 11552
rect 12952 11540 12958 11552
rect 13265 11543 13323 11549
rect 13265 11540 13277 11543
rect 12952 11512 13277 11540
rect 12952 11500 12958 11512
rect 13265 11509 13277 11512
rect 13311 11509 13323 11543
rect 13814 11540 13820 11552
rect 13775 11512 13820 11540
rect 13265 11503 13323 11509
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 14826 11500 14832 11552
rect 14884 11540 14890 11552
rect 15764 11540 15792 11580
rect 16666 11540 16672 11552
rect 14884 11512 15792 11540
rect 16627 11512 16672 11540
rect 14884 11500 14890 11512
rect 16666 11500 16672 11512
rect 16724 11500 16730 11552
rect 17880 11540 17908 11707
rect 19260 11608 19288 11716
rect 19705 11713 19717 11747
rect 19751 11713 19763 11747
rect 19705 11707 19763 11713
rect 19812 11676 19840 11852
rect 19904 11852 22928 11880
rect 19904 11753 19932 11852
rect 22922 11840 22928 11852
rect 22980 11840 22986 11892
rect 23290 11880 23296 11892
rect 23251 11852 23296 11880
rect 23290 11840 23296 11852
rect 23348 11840 23354 11892
rect 23842 11840 23848 11892
rect 23900 11880 23906 11892
rect 26421 11883 26479 11889
rect 23900 11852 26096 11880
rect 23900 11840 23906 11852
rect 22180 11815 22238 11821
rect 22180 11781 22192 11815
rect 22226 11812 22238 11815
rect 24854 11812 24860 11824
rect 22226 11784 24860 11812
rect 22226 11781 22238 11784
rect 22180 11775 22238 11781
rect 24854 11772 24860 11784
rect 24912 11772 24918 11824
rect 26068 11821 26096 11852
rect 26421 11849 26433 11883
rect 26467 11880 26479 11883
rect 27706 11880 27712 11892
rect 26467 11852 27712 11880
rect 26467 11849 26479 11852
rect 26421 11843 26479 11849
rect 27706 11840 27712 11852
rect 27764 11840 27770 11892
rect 28258 11840 28264 11892
rect 28316 11880 28322 11892
rect 28353 11883 28411 11889
rect 28353 11880 28365 11883
rect 28316 11852 28365 11880
rect 28316 11840 28322 11852
rect 28353 11849 28365 11852
rect 28399 11849 28411 11883
rect 28353 11843 28411 11849
rect 26053 11815 26111 11821
rect 26053 11781 26065 11815
rect 26099 11812 26111 11815
rect 26510 11812 26516 11824
rect 26099 11784 26516 11812
rect 26099 11781 26111 11784
rect 26053 11775 26111 11781
rect 26510 11772 26516 11784
rect 26568 11772 26574 11824
rect 27246 11821 27252 11824
rect 27240 11812 27252 11821
rect 27207 11784 27252 11812
rect 27240 11775 27252 11784
rect 27246 11772 27252 11775
rect 27304 11772 27310 11824
rect 19889 11747 19947 11753
rect 19889 11713 19901 11747
rect 19935 11713 19947 11747
rect 19889 11707 19947 11713
rect 20257 11747 20315 11753
rect 20257 11713 20269 11747
rect 20303 11744 20315 11747
rect 20346 11744 20352 11756
rect 20303 11716 20352 11744
rect 20303 11713 20315 11716
rect 20257 11707 20315 11713
rect 20346 11704 20352 11716
rect 20404 11704 20410 11756
rect 21269 11747 21327 11753
rect 21269 11713 21281 11747
rect 21315 11744 21327 11747
rect 21450 11744 21456 11756
rect 21315 11716 21456 11744
rect 21315 11713 21327 11716
rect 21269 11707 21327 11713
rect 21450 11704 21456 11716
rect 21508 11704 21514 11756
rect 21910 11744 21916 11756
rect 21871 11716 21916 11744
rect 21910 11704 21916 11716
rect 21968 11704 21974 11756
rect 23750 11744 23756 11756
rect 22020 11716 23756 11744
rect 19981 11679 20039 11685
rect 19981 11676 19993 11679
rect 19812 11648 19993 11676
rect 19981 11645 19993 11648
rect 20027 11645 20039 11679
rect 19981 11639 20039 11645
rect 20073 11679 20131 11685
rect 20073 11645 20085 11679
rect 20119 11676 20131 11679
rect 22020 11676 22048 11716
rect 23750 11704 23756 11716
rect 23808 11704 23814 11756
rect 25317 11747 25375 11753
rect 25317 11744 25329 11747
rect 23860 11716 25329 11744
rect 20119 11648 22048 11676
rect 20119 11645 20131 11648
rect 20073 11639 20131 11645
rect 23106 11636 23112 11688
rect 23164 11676 23170 11688
rect 23860 11676 23888 11716
rect 25317 11713 25329 11716
rect 25363 11713 25375 11747
rect 25317 11707 25375 11713
rect 26237 11747 26295 11753
rect 26237 11713 26249 11747
rect 26283 11744 26295 11747
rect 26418 11744 26424 11756
rect 26283 11716 26424 11744
rect 26283 11713 26295 11716
rect 26237 11707 26295 11713
rect 26418 11704 26424 11716
rect 26476 11744 26482 11756
rect 26786 11744 26792 11756
rect 26476 11716 26792 11744
rect 26476 11704 26482 11716
rect 26786 11704 26792 11716
rect 26844 11704 26850 11756
rect 28074 11744 28080 11756
rect 26896 11716 28080 11744
rect 23164 11648 23888 11676
rect 23164 11636 23170 11648
rect 23934 11636 23940 11688
rect 23992 11676 23998 11688
rect 24210 11676 24216 11688
rect 23992 11648 24037 11676
rect 24171 11648 24216 11676
rect 23992 11636 23998 11648
rect 24210 11636 24216 11648
rect 24268 11636 24274 11688
rect 25038 11636 25044 11688
rect 25096 11676 25102 11688
rect 25501 11679 25559 11685
rect 25501 11676 25513 11679
rect 25096 11648 25513 11676
rect 25096 11636 25102 11648
rect 25501 11645 25513 11648
rect 25547 11676 25559 11679
rect 26896 11676 26924 11716
rect 28074 11704 28080 11716
rect 28132 11704 28138 11756
rect 28994 11744 29000 11756
rect 28955 11716 29000 11744
rect 28994 11704 29000 11716
rect 29052 11704 29058 11756
rect 25547 11648 26924 11676
rect 26973 11679 27031 11685
rect 25547 11645 25559 11648
rect 25501 11639 25559 11645
rect 26973 11645 26985 11679
rect 27019 11645 27031 11679
rect 26973 11639 27031 11645
rect 20441 11611 20499 11617
rect 20441 11608 20453 11611
rect 19260 11580 20453 11608
rect 20441 11577 20453 11580
rect 20487 11577 20499 11611
rect 20441 11571 20499 11577
rect 21085 11611 21143 11617
rect 21085 11577 21097 11611
rect 21131 11608 21143 11611
rect 21726 11608 21732 11620
rect 21131 11580 21732 11608
rect 21131 11577 21143 11580
rect 21085 11571 21143 11577
rect 21726 11568 21732 11580
rect 21784 11568 21790 11620
rect 23492 11580 25544 11608
rect 20714 11540 20720 11552
rect 17880 11512 20720 11540
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 21542 11500 21548 11552
rect 21600 11540 21606 11552
rect 22186 11540 22192 11552
rect 21600 11512 22192 11540
rect 21600 11500 21606 11512
rect 22186 11500 22192 11512
rect 22244 11500 22250 11552
rect 22278 11500 22284 11552
rect 22336 11540 22342 11552
rect 23492 11540 23520 11580
rect 22336 11512 23520 11540
rect 25516 11540 25544 11580
rect 26878 11568 26884 11620
rect 26936 11608 26942 11620
rect 26988 11608 27016 11639
rect 26936 11580 27016 11608
rect 26936 11568 26942 11580
rect 28813 11543 28871 11549
rect 28813 11540 28825 11543
rect 25516 11512 28825 11540
rect 22336 11500 22342 11512
rect 28813 11509 28825 11512
rect 28859 11509 28871 11543
rect 28813 11503 28871 11509
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 7193 11339 7251 11345
rect 7193 11305 7205 11339
rect 7239 11305 7251 11339
rect 7193 11299 7251 11305
rect 8021 11339 8079 11345
rect 8021 11305 8033 11339
rect 8067 11336 8079 11339
rect 9950 11336 9956 11348
rect 8067 11308 9956 11336
rect 8067 11305 8079 11308
rect 8021 11299 8079 11305
rect 7208 11268 7236 11299
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 10152 11308 12296 11336
rect 8294 11268 8300 11280
rect 7208 11240 8300 11268
rect 8294 11228 8300 11240
rect 8352 11228 8358 11280
rect 9398 11228 9404 11280
rect 9456 11268 9462 11280
rect 10152 11268 10180 11308
rect 9456 11240 10180 11268
rect 10229 11271 10287 11277
rect 9456 11228 9462 11240
rect 10229 11237 10241 11271
rect 10275 11268 10287 11271
rect 11330 11268 11336 11280
rect 10275 11240 11336 11268
rect 10275 11237 10287 11240
rect 10229 11231 10287 11237
rect 11330 11228 11336 11240
rect 11388 11228 11394 11280
rect 12268 11268 12296 11308
rect 12342 11296 12348 11348
rect 12400 11336 12406 11348
rect 12897 11339 12955 11345
rect 12897 11336 12909 11339
rect 12400 11308 12909 11336
rect 12400 11296 12406 11308
rect 12897 11305 12909 11308
rect 12943 11305 12955 11339
rect 14182 11336 14188 11348
rect 14143 11308 14188 11336
rect 12897 11299 12955 11305
rect 14182 11296 14188 11308
rect 14240 11296 14246 11348
rect 14918 11336 14924 11348
rect 14879 11308 14924 11336
rect 14918 11296 14924 11308
rect 14976 11296 14982 11348
rect 15473 11339 15531 11345
rect 15473 11305 15485 11339
rect 15519 11336 15531 11339
rect 16758 11336 16764 11348
rect 15519 11308 16764 11336
rect 15519 11305 15531 11308
rect 15473 11299 15531 11305
rect 16758 11296 16764 11308
rect 16816 11336 16822 11348
rect 17218 11336 17224 11348
rect 16816 11308 17224 11336
rect 16816 11296 16822 11308
rect 17218 11296 17224 11308
rect 17276 11296 17282 11348
rect 18046 11296 18052 11348
rect 18104 11336 18110 11348
rect 20990 11336 20996 11348
rect 18104 11308 20116 11336
rect 18104 11296 18110 11308
rect 13078 11268 13084 11280
rect 12268 11240 13084 11268
rect 13078 11228 13084 11240
rect 13136 11228 13142 11280
rect 15838 11268 15844 11280
rect 14108 11240 15844 11268
rect 5813 11203 5871 11209
rect 5813 11200 5825 11203
rect 4816 11172 5825 11200
rect 4816 11141 4844 11172
rect 5813 11169 5825 11172
rect 5859 11169 5871 11203
rect 7190 11200 7196 11212
rect 5813 11163 5871 11169
rect 6748 11172 7196 11200
rect 4801 11135 4859 11141
rect 4801 11101 4813 11135
rect 4847 11101 4859 11135
rect 4801 11095 4859 11101
rect 5537 11135 5595 11141
rect 5537 11101 5549 11135
rect 5583 11101 5595 11135
rect 5537 11095 5595 11101
rect 5629 11135 5687 11141
rect 5629 11101 5641 11135
rect 5675 11132 5687 11135
rect 6748 11132 6776 11172
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 7653 11203 7711 11209
rect 7653 11169 7665 11203
rect 7699 11200 7711 11203
rect 7699 11172 7972 11200
rect 7699 11169 7711 11172
rect 7653 11163 7711 11169
rect 6914 11132 6920 11144
rect 5675 11104 6776 11132
rect 6875 11104 6920 11132
rect 5675 11101 5687 11104
rect 5629 11095 5687 11101
rect 5442 11024 5448 11076
rect 5500 11064 5506 11076
rect 5552 11064 5580 11095
rect 6914 11092 6920 11104
rect 6972 11092 6978 11144
rect 7012 11129 7070 11135
rect 7012 11095 7024 11129
rect 7058 11095 7070 11129
rect 6932 11064 6960 11092
rect 7012 11089 7070 11095
rect 7098 11092 7104 11144
rect 7156 11132 7162 11144
rect 7668 11132 7696 11163
rect 7834 11132 7840 11144
rect 7156 11104 7696 11132
rect 7795 11104 7840 11132
rect 7156 11092 7162 11104
rect 7834 11092 7840 11104
rect 7892 11092 7898 11144
rect 7944 11132 7972 11172
rect 8018 11160 8024 11212
rect 8076 11200 8082 11212
rect 12342 11200 12348 11212
rect 8076 11172 9168 11200
rect 8076 11160 8082 11172
rect 8110 11132 8116 11144
rect 7944 11104 8116 11132
rect 8110 11092 8116 11104
rect 8168 11132 8174 11144
rect 9140 11141 9168 11172
rect 10428 11172 12348 11200
rect 10428 11141 10456 11172
rect 12342 11160 12348 11172
rect 12400 11160 12406 11212
rect 12526 11160 12532 11212
rect 12584 11200 12590 11212
rect 12894 11200 12900 11212
rect 12584 11172 12629 11200
rect 12855 11172 12900 11200
rect 12584 11160 12590 11172
rect 12894 11160 12900 11172
rect 12952 11160 12958 11212
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 8168 11104 8953 11132
rect 8168 11092 8174 11104
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11101 9183 11135
rect 9125 11095 9183 11101
rect 10413 11135 10471 11141
rect 10413 11101 10425 11135
rect 10459 11101 10471 11135
rect 10962 11132 10968 11144
rect 10923 11104 10968 11132
rect 10413 11095 10471 11101
rect 10962 11092 10968 11104
rect 11020 11092 11026 11144
rect 11885 11135 11943 11141
rect 11885 11101 11897 11135
rect 11931 11132 11943 11135
rect 12084 11132 12296 11134
rect 12434 11132 12440 11144
rect 11931 11106 12440 11132
rect 11931 11104 12112 11106
rect 12268 11104 12440 11106
rect 11931 11101 11943 11104
rect 11885 11095 11943 11101
rect 12434 11092 12440 11104
rect 12492 11092 12498 11144
rect 14108 11141 14136 11240
rect 15838 11228 15844 11240
rect 15896 11228 15902 11280
rect 19429 11271 19487 11277
rect 19429 11237 19441 11271
rect 19475 11268 19487 11271
rect 19518 11268 19524 11280
rect 19475 11240 19524 11268
rect 19475 11237 19487 11240
rect 19429 11231 19487 11237
rect 19518 11228 19524 11240
rect 19576 11228 19582 11280
rect 16666 11200 16672 11212
rect 15672 11172 16672 11200
rect 14093 11135 14151 11141
rect 14093 11101 14105 11135
rect 14139 11101 14151 11135
rect 14093 11095 14151 11101
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11132 14335 11135
rect 14458 11132 14464 11144
rect 14323 11104 14464 11132
rect 14323 11101 14335 11104
rect 14277 11095 14335 11101
rect 14458 11092 14464 11104
rect 14516 11132 14522 11144
rect 14918 11132 14924 11144
rect 14516 11104 14924 11132
rect 14516 11092 14522 11104
rect 14918 11092 14924 11104
rect 14976 11092 14982 11144
rect 15470 11092 15476 11144
rect 15528 11092 15534 11144
rect 15672 11141 15700 11172
rect 16666 11160 16672 11172
rect 16724 11160 16730 11212
rect 16945 11203 17003 11209
rect 16945 11169 16957 11203
rect 16991 11200 17003 11203
rect 17126 11200 17132 11212
rect 16991 11172 17132 11200
rect 16991 11169 17003 11172
rect 16945 11163 17003 11169
rect 17126 11160 17132 11172
rect 17184 11160 17190 11212
rect 17310 11160 17316 11212
rect 17368 11200 17374 11212
rect 17405 11203 17463 11209
rect 17405 11200 17417 11203
rect 17368 11172 17417 11200
rect 17368 11160 17374 11172
rect 17405 11169 17417 11172
rect 17451 11200 17463 11203
rect 17678 11200 17684 11212
rect 17451 11172 17684 11200
rect 17451 11169 17463 11172
rect 17405 11163 17463 11169
rect 17678 11160 17684 11172
rect 17736 11160 17742 11212
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11101 15715 11135
rect 15838 11132 15844 11144
rect 15799 11104 15844 11132
rect 15657 11095 15715 11101
rect 15838 11092 15844 11104
rect 15896 11092 15902 11144
rect 16117 11135 16175 11141
rect 16117 11101 16129 11135
rect 16163 11101 16175 11135
rect 16574 11132 16580 11144
rect 16535 11104 16580 11132
rect 16117 11095 16175 11101
rect 5500 11036 6960 11064
rect 5500 11024 5506 11036
rect 7024 11008 7052 11089
rect 7282 11024 7288 11076
rect 7340 11064 7346 11076
rect 9309 11067 9367 11073
rect 9309 11064 9321 11067
rect 7340 11036 9321 11064
rect 7340 11024 7346 11036
rect 9309 11033 9321 11036
rect 9355 11033 9367 11067
rect 9309 11027 9367 11033
rect 9674 11024 9680 11076
rect 9732 11064 9738 11076
rect 11149 11067 11207 11073
rect 11149 11064 11161 11067
rect 9732 11036 11161 11064
rect 9732 11024 9738 11036
rect 11149 11033 11161 11036
rect 11195 11033 11207 11067
rect 11149 11027 11207 11033
rect 11790 11024 11796 11076
rect 11848 11064 11854 11076
rect 12069 11067 12127 11073
rect 12069 11064 12081 11067
rect 11848 11036 12081 11064
rect 11848 11024 11854 11036
rect 12069 11033 12081 11036
rect 12115 11033 12127 11067
rect 14826 11064 14832 11076
rect 14787 11036 14832 11064
rect 12069 11027 12127 11033
rect 14826 11024 14832 11036
rect 14884 11024 14890 11076
rect 15488 11064 15516 11092
rect 15749 11067 15807 11073
rect 15749 11064 15761 11067
rect 15488 11036 15761 11064
rect 15749 11033 15761 11036
rect 15795 11033 15807 11067
rect 15749 11027 15807 11033
rect 15979 11067 16037 11073
rect 15979 11033 15991 11067
rect 16025 11033 16037 11067
rect 16132 11064 16160 11095
rect 16574 11092 16580 11104
rect 16632 11092 16638 11144
rect 16850 11132 16856 11144
rect 16811 11104 16856 11132
rect 16850 11092 16856 11104
rect 16908 11132 16914 11144
rect 17589 11135 17647 11141
rect 17589 11132 17601 11135
rect 16908 11104 17601 11132
rect 16908 11092 16914 11104
rect 17589 11101 17601 11104
rect 17635 11101 17647 11135
rect 17589 11095 17647 11101
rect 17773 11135 17831 11141
rect 17773 11101 17785 11135
rect 17819 11132 17831 11135
rect 19245 11135 19303 11141
rect 17819 11104 19196 11132
rect 17819 11101 17831 11104
rect 17773 11095 17831 11101
rect 17862 11064 17868 11076
rect 16132 11036 17868 11064
rect 15979 11027 16037 11033
rect 4614 10996 4620 11008
rect 4575 10968 4620 10996
rect 4614 10956 4620 10968
rect 4672 10956 4678 11008
rect 7006 10956 7012 11008
rect 7064 10956 7070 11008
rect 7098 10956 7104 11008
rect 7156 10996 7162 11008
rect 9582 10996 9588 11008
rect 7156 10968 9588 10996
rect 7156 10956 7162 10968
rect 9582 10956 9588 10968
rect 9640 10956 9646 11008
rect 11054 10956 11060 11008
rect 11112 10996 11118 11008
rect 12526 10996 12532 11008
rect 11112 10968 12532 10996
rect 11112 10956 11118 10968
rect 12526 10956 12532 10968
rect 12584 10956 12590 11008
rect 12618 10956 12624 11008
rect 12676 10996 12682 11008
rect 12713 10999 12771 11005
rect 12713 10996 12725 10999
rect 12676 10968 12725 10996
rect 12676 10956 12682 10968
rect 12713 10965 12725 10968
rect 12759 10965 12771 10999
rect 15994 10996 16022 11027
rect 17862 11024 17868 11036
rect 17920 11024 17926 11076
rect 18325 11067 18383 11073
rect 18325 11033 18337 11067
rect 18371 11033 18383 11067
rect 18325 11027 18383 11033
rect 17126 10996 17132 11008
rect 15994 10968 17132 10996
rect 12713 10959 12771 10965
rect 17126 10956 17132 10968
rect 17184 10996 17190 11008
rect 18340 10996 18368 11027
rect 18414 11024 18420 11076
rect 18472 11064 18478 11076
rect 18509 11067 18567 11073
rect 18509 11064 18521 11067
rect 18472 11036 18521 11064
rect 18472 11024 18478 11036
rect 18509 11033 18521 11036
rect 18555 11033 18567 11067
rect 19168 11064 19196 11104
rect 19245 11101 19257 11135
rect 19291 11132 19303 11135
rect 19978 11132 19984 11144
rect 19291 11104 19984 11132
rect 19291 11101 19303 11104
rect 19245 11095 19303 11101
rect 19978 11092 19984 11104
rect 20036 11092 20042 11144
rect 20088 11141 20116 11308
rect 20272 11308 20996 11336
rect 20272 11141 20300 11308
rect 20990 11296 20996 11308
rect 21048 11296 21054 11348
rect 21177 11339 21235 11345
rect 21177 11305 21189 11339
rect 21223 11336 21235 11339
rect 21634 11336 21640 11348
rect 21223 11308 21640 11336
rect 21223 11305 21235 11308
rect 21177 11299 21235 11305
rect 21634 11296 21640 11308
rect 21692 11296 21698 11348
rect 22557 11339 22615 11345
rect 22557 11305 22569 11339
rect 22603 11336 22615 11339
rect 26234 11336 26240 11348
rect 22603 11308 26240 11336
rect 22603 11305 22615 11308
rect 22557 11299 22615 11305
rect 26234 11296 26240 11308
rect 26292 11296 26298 11348
rect 27062 11336 27068 11348
rect 27023 11308 27068 11336
rect 27062 11296 27068 11308
rect 27120 11296 27126 11348
rect 21358 11228 21364 11280
rect 21416 11268 21422 11280
rect 21416 11240 23244 11268
rect 21416 11228 21422 11240
rect 23106 11200 23112 11212
rect 20073 11135 20131 11141
rect 20073 11101 20085 11135
rect 20119 11101 20131 11135
rect 20073 11095 20131 11101
rect 20221 11135 20300 11141
rect 20221 11101 20233 11135
rect 20267 11104 20300 11135
rect 20364 11172 23112 11200
rect 20267 11101 20279 11104
rect 20221 11095 20279 11101
rect 20364 11073 20392 11172
rect 23106 11160 23112 11172
rect 23164 11160 23170 11212
rect 20579 11135 20637 11141
rect 20579 11101 20591 11135
rect 20625 11132 20637 11135
rect 20898 11132 20904 11144
rect 20625 11104 20904 11132
rect 20625 11101 20637 11104
rect 20579 11095 20637 11101
rect 20898 11092 20904 11104
rect 20956 11132 20962 11144
rect 21361 11135 21419 11141
rect 20956 11104 21328 11132
rect 20956 11092 20962 11104
rect 20349 11067 20407 11073
rect 20349 11064 20361 11067
rect 19168 11036 20361 11064
rect 18509 11027 18567 11033
rect 20349 11033 20361 11036
rect 20395 11033 20407 11067
rect 20349 11027 20407 11033
rect 20441 11067 20499 11073
rect 20441 11033 20453 11067
rect 20487 11064 20499 11067
rect 20990 11064 20996 11076
rect 20487 11036 20996 11064
rect 20487 11033 20499 11036
rect 20441 11027 20499 11033
rect 20990 11024 20996 11036
rect 21048 11024 21054 11076
rect 21300 11064 21328 11104
rect 21361 11101 21373 11135
rect 21407 11132 21419 11135
rect 21634 11132 21640 11144
rect 21407 11104 21640 11132
rect 21407 11101 21419 11104
rect 21361 11095 21419 11101
rect 21634 11092 21640 11104
rect 21692 11092 21698 11144
rect 21744 11104 23060 11132
rect 21744 11064 21772 11104
rect 21300 11036 21772 11064
rect 22189 11067 22247 11073
rect 22189 11033 22201 11067
rect 22235 11064 22247 11067
rect 22373 11067 22431 11073
rect 22235 11036 22324 11064
rect 22235 11033 22247 11036
rect 22189 11027 22247 11033
rect 17184 10968 18368 10996
rect 20717 10999 20775 11005
rect 17184 10956 17190 10968
rect 20717 10965 20729 10999
rect 20763 10996 20775 10999
rect 20898 10996 20904 11008
rect 20763 10968 20904 10996
rect 20763 10965 20775 10968
rect 20717 10959 20775 10965
rect 20898 10956 20904 10968
rect 20956 10956 20962 11008
rect 22296 10996 22324 11036
rect 22373 11033 22385 11067
rect 22419 11064 22431 11067
rect 22646 11064 22652 11076
rect 22419 11036 22652 11064
rect 22419 11033 22431 11036
rect 22373 11027 22431 11033
rect 22646 11024 22652 11036
rect 22704 11024 22710 11076
rect 22922 11064 22928 11076
rect 22756 11036 22928 11064
rect 22756 10996 22784 11036
rect 22922 11024 22928 11036
rect 22980 11024 22986 11076
rect 22296 10968 22784 10996
rect 23032 10996 23060 11104
rect 23124 11064 23152 11160
rect 23216 11141 23244 11240
rect 23290 11228 23296 11280
rect 23348 11268 23354 11280
rect 24210 11268 24216 11280
rect 23348 11240 24216 11268
rect 23348 11228 23354 11240
rect 24210 11228 24216 11240
rect 24268 11228 24274 11280
rect 28261 11271 28319 11277
rect 28261 11237 28273 11271
rect 28307 11237 28319 11271
rect 29546 11268 29552 11280
rect 29507 11240 29552 11268
rect 28261 11231 28319 11237
rect 24302 11200 24308 11212
rect 23308 11172 24308 11200
rect 23308 11141 23336 11172
rect 24302 11160 24308 11172
rect 24360 11160 24366 11212
rect 28276 11200 28304 11231
rect 29546 11228 29552 11240
rect 29604 11228 29610 11280
rect 26436 11172 28304 11200
rect 23201 11135 23259 11141
rect 23201 11101 23213 11135
rect 23247 11101 23259 11135
rect 23201 11095 23259 11101
rect 23294 11135 23352 11141
rect 23294 11101 23306 11135
rect 23340 11101 23352 11135
rect 23566 11132 23572 11144
rect 23527 11104 23572 11132
rect 23294 11095 23352 11101
rect 23566 11092 23572 11104
rect 23624 11092 23630 11144
rect 23666 11135 23724 11141
rect 23666 11101 23678 11135
rect 23712 11132 23724 11135
rect 24210 11132 24216 11144
rect 23712 11104 24216 11132
rect 23712 11101 23724 11104
rect 23666 11095 23724 11101
rect 23477 11067 23535 11073
rect 23477 11064 23489 11067
rect 23124 11036 23489 11064
rect 23477 11033 23489 11036
rect 23523 11033 23535 11067
rect 23477 11027 23535 11033
rect 23681 10996 23709 11095
rect 24210 11092 24216 11104
rect 24268 11092 24274 11144
rect 24394 11132 24400 11144
rect 24355 11104 24400 11132
rect 24394 11092 24400 11104
rect 24452 11092 24458 11144
rect 24664 11135 24722 11141
rect 24664 11101 24676 11135
rect 24710 11132 24722 11135
rect 26436 11132 26464 11172
rect 24710 11104 26464 11132
rect 24710 11101 24722 11104
rect 24664 11095 24722 11101
rect 26510 11092 26516 11144
rect 26568 11132 26574 11144
rect 26697 11135 26755 11141
rect 26697 11132 26709 11135
rect 26568 11104 26709 11132
rect 26568 11092 26574 11104
rect 26697 11101 26709 11104
rect 26743 11101 26755 11135
rect 27614 11132 27620 11144
rect 27575 11104 27620 11132
rect 26697 11095 26755 11101
rect 27614 11092 27620 11104
rect 27672 11092 27678 11144
rect 28442 11132 28448 11144
rect 28403 11104 28448 11132
rect 28442 11092 28448 11104
rect 28500 11092 28506 11144
rect 29730 11132 29736 11144
rect 29691 11104 29736 11132
rect 29730 11092 29736 11104
rect 29788 11092 29794 11144
rect 23750 11024 23756 11076
rect 23808 11064 23814 11076
rect 24118 11064 24124 11076
rect 23808 11036 24124 11064
rect 23808 11024 23814 11036
rect 23860 11005 23888 11036
rect 24118 11024 24124 11036
rect 24176 11024 24182 11076
rect 24302 11024 24308 11076
rect 24360 11064 24366 11076
rect 24360 11036 25900 11064
rect 24360 11024 24366 11036
rect 23032 10968 23709 10996
rect 23845 10999 23903 11005
rect 23845 10965 23857 10999
rect 23891 10965 23903 10999
rect 25774 10996 25780 11008
rect 25735 10968 25780 10996
rect 23845 10959 23903 10965
rect 25774 10956 25780 10968
rect 25832 10956 25838 11008
rect 25872 10996 25900 11036
rect 26142 11024 26148 11076
rect 26200 11064 26206 11076
rect 26881 11067 26939 11073
rect 26881 11064 26893 11067
rect 26200 11036 26893 11064
rect 26200 11024 26206 11036
rect 26881 11033 26893 11036
rect 26927 11033 26939 11067
rect 26881 11027 26939 11033
rect 27062 11024 27068 11076
rect 27120 11064 27126 11076
rect 27801 11067 27859 11073
rect 27801 11064 27813 11067
rect 27120 11036 27813 11064
rect 27120 11024 27126 11036
rect 27801 11033 27813 11036
rect 27847 11033 27859 11067
rect 27801 11027 27859 11033
rect 29472 11036 29776 11064
rect 29472 10996 29500 11036
rect 25872 10968 29500 10996
rect 29748 10996 29776 11036
rect 36262 10996 36268 11008
rect 29748 10968 36268 10996
rect 36262 10956 36268 10968
rect 36320 10956 36326 11008
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 198 10752 204 10804
rect 256 10792 262 10804
rect 6454 10792 6460 10804
rect 256 10764 2774 10792
rect 6415 10764 6460 10792
rect 256 10752 262 10764
rect 2746 10724 2774 10764
rect 6454 10752 6460 10764
rect 6512 10752 6518 10804
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7282 10792 7288 10804
rect 6972 10764 7288 10792
rect 6972 10752 6978 10764
rect 7282 10752 7288 10764
rect 7340 10752 7346 10804
rect 7653 10795 7711 10801
rect 7653 10761 7665 10795
rect 7699 10792 7711 10795
rect 7834 10792 7840 10804
rect 7699 10764 7840 10792
rect 7699 10761 7711 10764
rect 7653 10755 7711 10761
rect 7834 10752 7840 10764
rect 7892 10752 7898 10804
rect 11790 10752 11796 10804
rect 11848 10792 11854 10804
rect 23385 10795 23443 10801
rect 11848 10764 17908 10792
rect 11848 10752 11854 10764
rect 17880 10733 17908 10764
rect 23385 10761 23397 10795
rect 23431 10792 23443 10795
rect 23566 10792 23572 10804
rect 23431 10764 23572 10792
rect 23431 10761 23443 10764
rect 23385 10755 23443 10761
rect 23566 10752 23572 10764
rect 23624 10752 23630 10804
rect 23676 10764 28948 10792
rect 17865 10727 17923 10733
rect 2746 10696 17264 10724
rect 4893 10659 4951 10665
rect 4893 10625 4905 10659
rect 4939 10656 4951 10659
rect 5629 10659 5687 10665
rect 4939 10628 5580 10656
rect 4939 10625 4951 10628
rect 4893 10619 4951 10625
rect 1854 10548 1860 10600
rect 1912 10588 1918 10600
rect 5442 10588 5448 10600
rect 1912 10560 2774 10588
rect 5403 10560 5448 10588
rect 1912 10548 1918 10560
rect 2746 10520 2774 10560
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 5552 10588 5580 10628
rect 5629 10625 5641 10659
rect 5675 10656 5687 10659
rect 6362 10656 6368 10668
rect 5675 10628 6368 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 6362 10616 6368 10628
rect 6420 10616 6426 10668
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 6914 10656 6920 10668
rect 6687 10628 6920 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 7098 10656 7104 10668
rect 7059 10628 7104 10656
rect 7098 10616 7104 10628
rect 7156 10616 7162 10668
rect 7282 10656 7288 10668
rect 7243 10628 7288 10656
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 7377 10659 7435 10665
rect 7377 10625 7389 10659
rect 7423 10625 7435 10659
rect 7377 10619 7435 10625
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10656 7527 10659
rect 7558 10656 7564 10668
rect 7515 10628 7564 10656
rect 7515 10625 7527 10628
rect 7469 10619 7527 10625
rect 5813 10591 5871 10597
rect 5813 10588 5825 10591
rect 5552 10560 5825 10588
rect 5813 10557 5825 10560
rect 5859 10557 5871 10591
rect 5813 10551 5871 10557
rect 7392 10520 7420 10619
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 8386 10656 8392 10668
rect 8347 10628 8392 10656
rect 8386 10616 8392 10628
rect 8444 10616 8450 10668
rect 8938 10616 8944 10668
rect 8996 10656 9002 10668
rect 9105 10659 9163 10665
rect 9105 10656 9117 10659
rect 8996 10628 9117 10656
rect 8996 10616 9002 10628
rect 9105 10625 9117 10628
rect 9151 10625 9163 10659
rect 9105 10619 9163 10625
rect 10781 10659 10839 10665
rect 10781 10625 10793 10659
rect 10827 10656 10839 10659
rect 11790 10656 11796 10668
rect 10827 10628 11796 10656
rect 10827 10625 10839 10628
rect 10781 10619 10839 10625
rect 11790 10616 11796 10628
rect 11848 10616 11854 10668
rect 12066 10656 12072 10668
rect 12027 10628 12072 10656
rect 12066 10616 12072 10628
rect 12124 10656 12130 10668
rect 12894 10656 12900 10668
rect 12124 10628 12900 10656
rect 12124 10616 12130 10628
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 13429 10659 13487 10665
rect 13429 10656 13441 10659
rect 13096 10628 13441 10656
rect 8849 10591 8907 10597
rect 8849 10557 8861 10591
rect 8895 10557 8907 10591
rect 12710 10588 12716 10600
rect 8849 10551 8907 10557
rect 10980 10560 12716 10588
rect 2746 10492 7420 10520
rect 4706 10452 4712 10464
rect 4667 10424 4712 10452
rect 4706 10412 4712 10424
rect 4764 10412 4770 10464
rect 8202 10452 8208 10464
rect 8163 10424 8208 10452
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 8864 10452 8892 10551
rect 10980 10532 11008 10560
rect 12710 10548 12716 10560
rect 12768 10548 12774 10600
rect 10410 10520 10416 10532
rect 9784 10492 10416 10520
rect 9784 10452 9812 10492
rect 10410 10480 10416 10492
rect 10468 10520 10474 10532
rect 10962 10520 10968 10532
rect 10468 10492 10968 10520
rect 10468 10480 10474 10492
rect 10962 10480 10968 10492
rect 11020 10480 11026 10532
rect 11330 10480 11336 10532
rect 11388 10520 11394 10532
rect 13096 10520 13124 10628
rect 13429 10625 13441 10628
rect 13475 10625 13487 10659
rect 15654 10656 15660 10668
rect 15615 10628 15660 10656
rect 13429 10619 13487 10625
rect 15654 10616 15660 10628
rect 15712 10616 15718 10668
rect 15838 10656 15844 10668
rect 15799 10628 15844 10656
rect 15838 10616 15844 10628
rect 15896 10616 15902 10668
rect 17126 10656 17132 10668
rect 17087 10628 17132 10656
rect 17126 10616 17132 10628
rect 17184 10616 17190 10668
rect 17236 10656 17264 10696
rect 17865 10693 17877 10727
rect 17911 10693 17923 10727
rect 19426 10724 19432 10736
rect 17865 10687 17923 10693
rect 17972 10696 19432 10724
rect 17972 10656 18000 10696
rect 19426 10684 19432 10696
rect 19484 10684 19490 10736
rect 20714 10724 20720 10736
rect 19628 10696 20720 10724
rect 18506 10656 18512 10668
rect 17236 10628 18000 10656
rect 18467 10628 18512 10656
rect 18506 10616 18512 10628
rect 18564 10616 18570 10668
rect 19628 10665 19656 10696
rect 20714 10684 20720 10696
rect 20772 10724 20778 10736
rect 20772 10696 22048 10724
rect 20772 10684 20778 10696
rect 19886 10665 19892 10668
rect 19613 10659 19671 10665
rect 19613 10625 19625 10659
rect 19659 10625 19671 10659
rect 19880 10656 19892 10665
rect 19847 10628 19892 10656
rect 19613 10619 19671 10625
rect 19880 10619 19892 10628
rect 19886 10616 19892 10619
rect 19944 10616 19950 10668
rect 22020 10665 22048 10696
rect 23290 10684 23296 10736
rect 23348 10724 23354 10736
rect 23676 10724 23704 10764
rect 24210 10724 24216 10736
rect 23348 10696 23704 10724
rect 24171 10696 24216 10724
rect 23348 10684 23354 10696
rect 24210 10684 24216 10696
rect 24268 10684 24274 10736
rect 25041 10727 25099 10733
rect 25041 10693 25053 10727
rect 25087 10693 25099 10727
rect 25041 10687 25099 10693
rect 26237 10727 26295 10733
rect 26237 10693 26249 10727
rect 26283 10724 26295 10727
rect 26510 10724 26516 10736
rect 26283 10696 26516 10724
rect 26283 10693 26295 10696
rect 26237 10687 26295 10693
rect 22278 10665 22284 10668
rect 22005 10659 22063 10665
rect 22005 10625 22017 10659
rect 22051 10625 22063 10659
rect 22272 10656 22284 10665
rect 22239 10628 22284 10656
rect 22005 10619 22063 10625
rect 22272 10619 22284 10628
rect 22278 10616 22284 10619
rect 22336 10616 22342 10668
rect 24854 10616 24860 10668
rect 24912 10656 24918 10668
rect 24912 10628 24957 10656
rect 24912 10616 24918 10628
rect 25056 10600 25084 10687
rect 26510 10684 26516 10696
rect 26568 10684 26574 10736
rect 25314 10665 25320 10668
rect 25129 10659 25187 10665
rect 25129 10625 25141 10659
rect 25175 10625 25187 10659
rect 25129 10619 25187 10625
rect 25271 10659 25320 10665
rect 25271 10625 25283 10659
rect 25317 10625 25320 10659
rect 25271 10619 25320 10625
rect 13173 10591 13231 10597
rect 13173 10557 13185 10591
rect 13219 10557 13231 10591
rect 13173 10551 13231 10557
rect 11388 10492 13124 10520
rect 11388 10480 11394 10492
rect 8864 10424 9812 10452
rect 9950 10412 9956 10464
rect 10008 10452 10014 10464
rect 10229 10455 10287 10461
rect 10229 10452 10241 10455
rect 10008 10424 10241 10452
rect 10008 10412 10014 10424
rect 10229 10421 10241 10424
rect 10275 10421 10287 10455
rect 10229 10415 10287 10421
rect 12161 10455 12219 10461
rect 12161 10421 12173 10455
rect 12207 10452 12219 10455
rect 12434 10452 12440 10464
rect 12207 10424 12440 10452
rect 12207 10421 12219 10424
rect 12161 10415 12219 10421
rect 12434 10412 12440 10424
rect 12492 10412 12498 10464
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 13188 10452 13216 10551
rect 17862 10548 17868 10600
rect 17920 10588 17926 10600
rect 18601 10591 18659 10597
rect 18601 10588 18613 10591
rect 17920 10560 18613 10588
rect 17920 10548 17926 10560
rect 18601 10557 18613 10560
rect 18647 10557 18659 10591
rect 18601 10551 18659 10557
rect 24397 10591 24455 10597
rect 24397 10557 24409 10591
rect 24443 10588 24455 10591
rect 24486 10588 24492 10600
rect 24443 10560 24492 10588
rect 24443 10557 24455 10560
rect 24397 10551 24455 10557
rect 24486 10548 24492 10560
rect 24544 10548 24550 10600
rect 25038 10548 25044 10600
rect 25096 10548 25102 10600
rect 14553 10523 14611 10529
rect 14553 10489 14565 10523
rect 14599 10520 14611 10523
rect 14826 10520 14832 10532
rect 14599 10492 14832 10520
rect 14599 10489 14611 10492
rect 14553 10483 14611 10489
rect 14826 10480 14832 10492
rect 14884 10480 14890 10532
rect 17313 10523 17371 10529
rect 17313 10489 17325 10523
rect 17359 10520 17371 10523
rect 18138 10520 18144 10532
rect 17359 10492 18144 10520
rect 17359 10489 17371 10492
rect 17313 10483 17371 10489
rect 18138 10480 18144 10492
rect 18196 10520 18202 10532
rect 19610 10520 19616 10532
rect 18196 10492 19616 10520
rect 18196 10480 18202 10492
rect 19610 10480 19616 10492
rect 19668 10480 19674 10532
rect 20990 10520 20996 10532
rect 20951 10492 20996 10520
rect 20990 10480 20996 10492
rect 21048 10480 21054 10532
rect 25139 10520 25167 10619
rect 25314 10616 25320 10619
rect 25372 10616 25378 10668
rect 27430 10656 27436 10668
rect 27391 10628 27436 10656
rect 27430 10616 27436 10628
rect 27488 10616 27494 10668
rect 27706 10616 27712 10668
rect 27764 10656 27770 10668
rect 28261 10659 28319 10665
rect 28261 10656 28273 10659
rect 27764 10628 28273 10656
rect 27764 10616 27770 10628
rect 28261 10625 28273 10628
rect 28307 10625 28319 10659
rect 28261 10619 28319 10625
rect 28442 10616 28448 10668
rect 28500 10656 28506 10668
rect 28920 10665 28948 10764
rect 28994 10684 29000 10736
rect 29052 10724 29058 10736
rect 29052 10696 29592 10724
rect 29052 10684 29058 10696
rect 29564 10665 29592 10696
rect 28905 10659 28963 10665
rect 28500 10628 28764 10656
rect 28500 10616 28506 10628
rect 27617 10591 27675 10597
rect 27617 10557 27629 10591
rect 27663 10588 27675 10591
rect 28626 10588 28632 10600
rect 27663 10560 28632 10588
rect 27663 10557 27675 10560
rect 27617 10551 27675 10557
rect 28626 10548 28632 10560
rect 28684 10548 28690 10600
rect 28736 10588 28764 10628
rect 28905 10625 28917 10659
rect 28951 10625 28963 10659
rect 28905 10619 28963 10625
rect 29365 10659 29423 10665
rect 29365 10625 29377 10659
rect 29411 10625 29423 10659
rect 29365 10619 29423 10625
rect 29549 10659 29607 10665
rect 29549 10625 29561 10659
rect 29595 10625 29607 10659
rect 30190 10656 30196 10668
rect 30151 10628 30196 10656
rect 29549 10619 29607 10625
rect 29380 10588 29408 10619
rect 30190 10616 30196 10628
rect 30248 10616 30254 10668
rect 30282 10616 30288 10668
rect 30340 10656 30346 10668
rect 30837 10659 30895 10665
rect 30837 10656 30849 10659
rect 30340 10628 30849 10656
rect 30340 10616 30346 10628
rect 30837 10625 30849 10628
rect 30883 10625 30895 10659
rect 30837 10619 30895 10625
rect 28736 10560 29408 10588
rect 25774 10520 25780 10532
rect 25139 10492 25780 10520
rect 25774 10480 25780 10492
rect 25832 10480 25838 10532
rect 28718 10520 28724 10532
rect 28679 10492 28724 10520
rect 28718 10480 28724 10492
rect 28776 10480 28782 10532
rect 28810 10480 28816 10532
rect 28868 10520 28874 10532
rect 30009 10523 30067 10529
rect 30009 10520 30021 10523
rect 28868 10492 30021 10520
rect 28868 10480 28874 10492
rect 30009 10489 30021 10492
rect 30055 10489 30067 10523
rect 30009 10483 30067 10489
rect 12768 10424 13216 10452
rect 12768 10412 12774 10424
rect 17862 10412 17868 10464
rect 17920 10452 17926 10464
rect 17957 10455 18015 10461
rect 17957 10452 17969 10455
rect 17920 10424 17969 10452
rect 17920 10412 17926 10424
rect 17957 10421 17969 10424
rect 18003 10421 18015 10455
rect 17957 10415 18015 10421
rect 18598 10412 18604 10464
rect 18656 10452 18662 10464
rect 24302 10452 24308 10464
rect 18656 10424 24308 10452
rect 18656 10412 18662 10424
rect 24302 10412 24308 10424
rect 24360 10412 24366 10464
rect 25406 10452 25412 10464
rect 25319 10424 25412 10452
rect 25406 10412 25412 10424
rect 25464 10452 25470 10464
rect 25866 10452 25872 10464
rect 25464 10424 25872 10452
rect 25464 10412 25470 10424
rect 25866 10412 25872 10424
rect 25924 10412 25930 10464
rect 26234 10412 26240 10464
rect 26292 10452 26298 10464
rect 26329 10455 26387 10461
rect 26329 10452 26341 10455
rect 26292 10424 26341 10452
rect 26292 10412 26298 10424
rect 26329 10421 26341 10424
rect 26375 10421 26387 10455
rect 26329 10415 26387 10421
rect 27614 10412 27620 10464
rect 27672 10452 27678 10464
rect 28077 10455 28135 10461
rect 28077 10452 28089 10455
rect 27672 10424 28089 10452
rect 27672 10412 27678 10424
rect 28077 10421 28089 10424
rect 28123 10421 28135 10455
rect 29362 10452 29368 10464
rect 29323 10424 29368 10452
rect 28077 10415 28135 10421
rect 29362 10412 29368 10424
rect 29420 10412 29426 10464
rect 30650 10452 30656 10464
rect 30611 10424 30656 10452
rect 30650 10412 30656 10424
rect 30708 10412 30714 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 6362 10248 6368 10260
rect 6323 10220 6368 10248
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 7006 10208 7012 10260
rect 7064 10248 7070 10260
rect 7653 10251 7711 10257
rect 7653 10248 7665 10251
rect 7064 10220 7665 10248
rect 7064 10208 7070 10220
rect 7653 10217 7665 10220
rect 7699 10217 7711 10251
rect 8110 10248 8116 10260
rect 8071 10220 8116 10248
rect 7653 10211 7711 10217
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 8386 10208 8392 10260
rect 8444 10248 8450 10260
rect 12805 10251 12863 10257
rect 12805 10248 12817 10251
rect 8444 10220 12817 10248
rect 8444 10208 8450 10220
rect 12805 10217 12817 10220
rect 12851 10217 12863 10251
rect 17034 10248 17040 10260
rect 12805 10211 12863 10217
rect 14844 10220 17040 10248
rect 7282 10180 7288 10192
rect 6104 10152 7288 10180
rect 5000 10084 5948 10112
rect 3970 10044 3976 10056
rect 3931 10016 3976 10044
rect 3970 10004 3976 10016
rect 4028 10004 4034 10056
rect 4240 10047 4298 10053
rect 4240 10013 4252 10047
rect 4286 10044 4298 10047
rect 4706 10044 4712 10056
rect 4286 10016 4712 10044
rect 4286 10013 4298 10016
rect 4240 10007 4298 10013
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 2958 9936 2964 9988
rect 3016 9976 3022 9988
rect 5000 9976 5028 10084
rect 5534 10044 5540 10056
rect 3016 9948 5028 9976
rect 5368 10016 5540 10044
rect 3016 9936 3022 9948
rect 5368 9917 5396 10016
rect 5534 10004 5540 10016
rect 5592 10044 5598 10056
rect 5813 10047 5871 10053
rect 5813 10044 5825 10047
rect 5592 10016 5825 10044
rect 5592 10004 5598 10016
rect 5813 10013 5825 10016
rect 5859 10013 5871 10047
rect 5813 10007 5871 10013
rect 5920 9976 5948 10084
rect 5997 10047 6055 10053
rect 5997 10013 6009 10047
rect 6043 10044 6055 10047
rect 6104 10044 6132 10152
rect 7282 10140 7288 10152
rect 7340 10180 7346 10192
rect 9171 10183 9229 10189
rect 9171 10180 9183 10183
rect 7340 10152 9183 10180
rect 7340 10140 7346 10152
rect 9171 10149 9183 10152
rect 9217 10149 9229 10183
rect 9171 10143 9229 10149
rect 12158 10140 12164 10192
rect 12216 10180 12222 10192
rect 14844 10180 14872 10220
rect 17034 10208 17040 10220
rect 17092 10208 17098 10260
rect 17221 10251 17279 10257
rect 17221 10217 17233 10251
rect 17267 10248 17279 10251
rect 18506 10248 18512 10260
rect 17267 10220 18512 10248
rect 17267 10217 17279 10220
rect 17221 10211 17279 10217
rect 18506 10208 18512 10220
rect 18564 10208 18570 10260
rect 20073 10251 20131 10257
rect 20073 10217 20085 10251
rect 20119 10248 20131 10251
rect 20993 10251 21051 10257
rect 20993 10248 21005 10251
rect 20119 10220 21005 10248
rect 20119 10217 20131 10220
rect 20073 10211 20131 10217
rect 20993 10217 21005 10220
rect 21039 10248 21051 10251
rect 21082 10248 21088 10260
rect 21039 10220 21088 10248
rect 21039 10217 21051 10220
rect 20993 10211 21051 10217
rect 20088 10180 20116 10211
rect 21082 10208 21088 10220
rect 21140 10208 21146 10260
rect 23290 10248 23296 10260
rect 21192 10220 23296 10248
rect 12216 10152 14872 10180
rect 18156 10152 20116 10180
rect 20257 10183 20315 10189
rect 12216 10140 12222 10152
rect 6196 10084 7512 10112
rect 6196 10053 6224 10084
rect 6043 10016 6132 10044
rect 6181 10047 6239 10053
rect 6043 10013 6055 10016
rect 5997 10007 6055 10013
rect 6181 10013 6193 10047
rect 6227 10013 6239 10047
rect 7098 10044 7104 10056
rect 7059 10016 7104 10044
rect 6181 10007 6239 10013
rect 7098 10004 7104 10016
rect 7156 10004 7162 10056
rect 7282 10044 7288 10056
rect 7243 10016 7288 10044
rect 7282 10004 7288 10016
rect 7340 10004 7346 10056
rect 7484 10053 7512 10084
rect 8202 10072 8208 10124
rect 8260 10112 8266 10124
rect 8260 10084 9536 10112
rect 8260 10072 8266 10084
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10044 7527 10047
rect 7558 10044 7564 10056
rect 7515 10016 7564 10044
rect 7515 10013 7527 10016
rect 7469 10007 7527 10013
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 8297 10047 8355 10053
rect 8297 10013 8309 10047
rect 8343 10044 8355 10047
rect 8846 10044 8852 10056
rect 8343 10016 8852 10044
rect 8343 10013 8355 10016
rect 8297 10007 8355 10013
rect 8846 10004 8852 10016
rect 8904 10004 8910 10056
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 6089 9979 6147 9985
rect 6089 9976 6101 9979
rect 5920 9948 6101 9976
rect 6089 9945 6101 9948
rect 6135 9945 6147 9979
rect 6089 9939 6147 9945
rect 6914 9936 6920 9988
rect 6972 9976 6978 9988
rect 7377 9979 7435 9985
rect 7377 9976 7389 9979
rect 6972 9948 7389 9976
rect 6972 9936 6978 9948
rect 7377 9945 7389 9948
rect 7423 9945 7435 9979
rect 7377 9939 7435 9945
rect 5353 9911 5411 9917
rect 5353 9877 5365 9911
rect 5399 9877 5411 9911
rect 8956 9908 8984 10007
rect 9508 9976 9536 10084
rect 12434 10072 12440 10124
rect 12492 10112 12498 10124
rect 13630 10112 13636 10124
rect 12492 10084 13636 10112
rect 12492 10072 12498 10084
rect 13630 10072 13636 10084
rect 13688 10072 13694 10124
rect 15194 10112 15200 10124
rect 14292 10084 15200 10112
rect 10597 10047 10655 10053
rect 10597 10013 10609 10047
rect 10643 10044 10655 10047
rect 12618 10044 12624 10056
rect 10643 10016 11008 10044
rect 12579 10016 12624 10044
rect 10643 10013 10655 10016
rect 10597 10007 10655 10013
rect 10980 9988 11008 10016
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 13357 10047 13415 10053
rect 13357 10013 13369 10047
rect 13403 10044 13415 10047
rect 14292 10044 14320 10084
rect 15194 10072 15200 10084
rect 15252 10072 15258 10124
rect 17126 10072 17132 10124
rect 17184 10112 17190 10124
rect 18156 10121 18184 10152
rect 20257 10149 20269 10183
rect 20303 10180 20315 10183
rect 21192 10180 21220 10220
rect 23290 10208 23296 10220
rect 23348 10208 23354 10260
rect 23474 10248 23480 10260
rect 23435 10220 23480 10248
rect 23474 10208 23480 10220
rect 23532 10208 23538 10260
rect 26694 10248 26700 10260
rect 24688 10220 26700 10248
rect 20303 10152 21220 10180
rect 22005 10183 22063 10189
rect 20303 10149 20315 10152
rect 20257 10143 20315 10149
rect 22005 10149 22017 10183
rect 22051 10180 22063 10183
rect 22646 10180 22652 10192
rect 22051 10152 22652 10180
rect 22051 10149 22063 10152
rect 22005 10143 22063 10149
rect 22646 10140 22652 10152
rect 22704 10140 22710 10192
rect 17865 10115 17923 10121
rect 17865 10112 17877 10115
rect 17184 10084 17877 10112
rect 17184 10072 17190 10084
rect 17865 10081 17877 10084
rect 17911 10081 17923 10115
rect 17865 10075 17923 10081
rect 18141 10115 18199 10121
rect 18141 10081 18153 10115
rect 18187 10081 18199 10115
rect 20346 10112 20352 10124
rect 18141 10075 18199 10081
rect 19352 10084 20352 10112
rect 14458 10044 14464 10056
rect 13403 10016 14320 10044
rect 14419 10016 14464 10044
rect 13403 10013 13415 10016
rect 13357 10007 13415 10013
rect 10842 9979 10900 9985
rect 10842 9976 10854 9979
rect 9508 9948 10854 9976
rect 10842 9945 10854 9948
rect 10888 9945 10900 9979
rect 10842 9939 10900 9945
rect 10962 9936 10968 9988
rect 11020 9936 11026 9988
rect 13372 9976 13400 10007
rect 14458 10004 14464 10016
rect 14516 10004 14522 10056
rect 14826 10044 14832 10056
rect 14787 10016 14832 10044
rect 14826 10004 14832 10016
rect 14884 10004 14890 10056
rect 15841 10047 15899 10053
rect 15841 10013 15853 10047
rect 15887 10044 15899 10047
rect 17770 10044 17776 10056
rect 15887 10016 17776 10044
rect 15887 10013 15899 10016
rect 15841 10007 15899 10013
rect 17770 10004 17776 10016
rect 17828 10004 17834 10056
rect 19251 10047 19309 10053
rect 19251 10013 19263 10047
rect 19297 10044 19309 10047
rect 19352 10044 19380 10084
rect 20346 10072 20352 10084
rect 20404 10112 20410 10124
rect 23750 10112 23756 10124
rect 20404 10084 23756 10112
rect 20404 10072 20410 10084
rect 23750 10072 23756 10084
rect 23808 10072 23814 10124
rect 19297 10016 19380 10044
rect 19297 10013 19309 10016
rect 19251 10007 19309 10013
rect 19426 10004 19432 10056
rect 19484 10044 19490 10056
rect 22189 10047 22247 10053
rect 19484 10016 19529 10044
rect 19484 10004 19490 10016
rect 22189 10013 22201 10047
rect 22235 10044 22247 10047
rect 22370 10044 22376 10056
rect 22235 10016 22376 10044
rect 22235 10013 22247 10016
rect 22189 10007 22247 10013
rect 22370 10004 22376 10016
rect 22428 10004 22434 10056
rect 22833 10047 22891 10053
rect 22833 10013 22845 10047
rect 22879 10013 22891 10047
rect 22833 10007 22891 10013
rect 23385 10047 23443 10053
rect 23385 10013 23397 10047
rect 23431 10044 23443 10047
rect 24688 10044 24716 10220
rect 26694 10208 26700 10220
rect 26752 10208 26758 10260
rect 26970 10208 26976 10260
rect 27028 10248 27034 10260
rect 27157 10251 27215 10257
rect 27157 10248 27169 10251
rect 27028 10220 27169 10248
rect 27028 10208 27034 10220
rect 27157 10217 27169 10220
rect 27203 10248 27215 10251
rect 27246 10248 27252 10260
rect 27203 10220 27252 10248
rect 27203 10217 27215 10220
rect 27157 10211 27215 10217
rect 27246 10208 27252 10220
rect 27304 10208 27310 10260
rect 27982 10208 27988 10260
rect 28040 10248 28046 10260
rect 28902 10248 28908 10260
rect 28040 10220 28908 10248
rect 28040 10208 28046 10220
rect 28902 10208 28908 10220
rect 28960 10208 28966 10260
rect 29178 10140 29184 10192
rect 29236 10180 29242 10192
rect 29549 10183 29607 10189
rect 29549 10180 29561 10183
rect 29236 10152 29561 10180
rect 29236 10140 29242 10152
rect 29549 10149 29561 10152
rect 29595 10149 29607 10183
rect 29549 10143 29607 10149
rect 26878 10072 26884 10124
rect 26936 10112 26942 10124
rect 27617 10115 27675 10121
rect 27617 10112 27629 10115
rect 26936 10084 27629 10112
rect 26936 10072 26942 10084
rect 27617 10081 27629 10084
rect 27663 10081 27675 10115
rect 27617 10075 27675 10081
rect 28718 10072 28724 10124
rect 28776 10112 28782 10124
rect 28776 10084 30420 10112
rect 28776 10072 28782 10084
rect 24946 10044 24952 10056
rect 23431 10016 24716 10044
rect 24907 10016 24952 10044
rect 23431 10013 23443 10016
rect 23385 10007 23443 10013
rect 11072 9948 13400 9976
rect 11072 9908 11100 9948
rect 13538 9936 13544 9988
rect 13596 9976 13602 9988
rect 14642 9976 14648 9988
rect 13596 9948 14648 9976
rect 13596 9936 13602 9948
rect 14642 9936 14648 9948
rect 14700 9936 14706 9988
rect 14737 9979 14795 9985
rect 14737 9945 14749 9979
rect 14783 9976 14795 9979
rect 16108 9979 16166 9985
rect 14783 9948 16068 9976
rect 14783 9945 14795 9948
rect 14737 9939 14795 9945
rect 8956 9880 11100 9908
rect 5353 9871 5411 9877
rect 11238 9868 11244 9920
rect 11296 9908 11302 9920
rect 11977 9911 12035 9917
rect 11977 9908 11989 9911
rect 11296 9880 11989 9908
rect 11296 9868 11302 9880
rect 11977 9877 11989 9880
rect 12023 9877 12035 9911
rect 11977 9871 12035 9877
rect 12342 9868 12348 9920
rect 12400 9908 12406 9920
rect 13722 9908 13728 9920
rect 12400 9880 13728 9908
rect 12400 9868 12406 9880
rect 13722 9868 13728 9880
rect 13780 9868 13786 9920
rect 14090 9868 14096 9920
rect 14148 9908 14154 9920
rect 15013 9911 15071 9917
rect 15013 9908 15025 9911
rect 14148 9880 15025 9908
rect 14148 9868 14154 9880
rect 15013 9877 15025 9880
rect 15059 9877 15071 9911
rect 16040 9908 16068 9948
rect 16108 9945 16120 9979
rect 16154 9976 16166 9979
rect 16390 9976 16396 9988
rect 16154 9948 16396 9976
rect 16154 9945 16166 9948
rect 16108 9939 16166 9945
rect 16390 9936 16396 9948
rect 16448 9936 16454 9988
rect 18598 9976 18604 9988
rect 17052 9948 18604 9976
rect 17052 9908 17080 9948
rect 18598 9936 18604 9948
rect 18656 9936 18662 9988
rect 19889 9979 19947 9985
rect 19889 9945 19901 9979
rect 19935 9976 19947 9979
rect 19978 9976 19984 9988
rect 19935 9948 19984 9976
rect 19935 9945 19947 9948
rect 19889 9939 19947 9945
rect 19978 9936 19984 9948
rect 20036 9976 20042 9988
rect 20438 9976 20444 9988
rect 20036 9948 20444 9976
rect 20036 9936 20042 9948
rect 20438 9936 20444 9948
rect 20496 9976 20502 9988
rect 20809 9979 20867 9985
rect 20809 9976 20821 9979
rect 20496 9948 20821 9976
rect 20496 9936 20502 9948
rect 20809 9945 20821 9948
rect 20855 9945 20867 9979
rect 20809 9939 20867 9945
rect 21025 9979 21083 9985
rect 21025 9945 21037 9979
rect 21071 9976 21083 9979
rect 21542 9976 21548 9988
rect 21071 9948 21548 9976
rect 21071 9945 21083 9948
rect 21025 9939 21083 9945
rect 21542 9936 21548 9948
rect 21600 9936 21606 9988
rect 22848 9976 22876 10007
rect 24946 10004 24952 10016
rect 25004 10004 25010 10056
rect 25133 10047 25191 10053
rect 25133 10013 25145 10047
rect 25179 10044 25191 10047
rect 25406 10044 25412 10056
rect 25179 10016 25412 10044
rect 25179 10013 25191 10016
rect 25133 10007 25191 10013
rect 25406 10004 25412 10016
rect 25464 10004 25470 10056
rect 25777 10047 25835 10053
rect 25777 10013 25789 10047
rect 25823 10044 25835 10047
rect 26896 10044 26924 10072
rect 25823 10016 26924 10044
rect 27884 10047 27942 10053
rect 25823 10013 25835 10016
rect 25777 10007 25835 10013
rect 27884 10013 27896 10047
rect 27930 10044 27942 10047
rect 29362 10044 29368 10056
rect 27930 10016 29368 10044
rect 27930 10013 27942 10016
rect 27884 10007 27942 10013
rect 23842 9976 23848 9988
rect 22848 9948 23848 9976
rect 23842 9936 23848 9948
rect 23900 9936 23906 9988
rect 25038 9936 25044 9988
rect 25096 9976 25102 9988
rect 25792 9976 25820 10007
rect 29362 10004 29368 10016
rect 29420 10004 29426 10056
rect 29730 10044 29736 10056
rect 29691 10016 29736 10044
rect 29730 10004 29736 10016
rect 29788 10004 29794 10056
rect 30392 10053 30420 10084
rect 30377 10047 30435 10053
rect 30377 10013 30389 10047
rect 30423 10013 30435 10047
rect 30377 10007 30435 10013
rect 31205 10047 31263 10053
rect 31205 10013 31217 10047
rect 31251 10013 31263 10047
rect 31205 10007 31263 10013
rect 25096 9948 25820 9976
rect 26044 9979 26102 9985
rect 25096 9936 25102 9948
rect 26044 9945 26056 9979
rect 26090 9976 26102 9979
rect 26878 9976 26884 9988
rect 26090 9948 26884 9976
rect 26090 9945 26102 9948
rect 26044 9939 26102 9945
rect 26878 9936 26884 9948
rect 26936 9936 26942 9988
rect 27430 9936 27436 9988
rect 27488 9976 27494 9988
rect 31220 9976 31248 10007
rect 27488 9948 31248 9976
rect 27488 9936 27494 9948
rect 19334 9908 19340 9920
rect 16040 9880 17080 9908
rect 19295 9880 19340 9908
rect 15013 9871 15071 9877
rect 19334 9868 19340 9880
rect 19392 9868 19398 9920
rect 20099 9911 20157 9917
rect 20099 9877 20111 9911
rect 20145 9908 20157 9911
rect 20898 9908 20904 9920
rect 20145 9880 20904 9908
rect 20145 9877 20157 9880
rect 20099 9871 20157 9877
rect 20898 9868 20904 9880
rect 20956 9868 20962 9920
rect 21174 9908 21180 9920
rect 21135 9880 21180 9908
rect 21174 9868 21180 9880
rect 21232 9868 21238 9920
rect 22649 9911 22707 9917
rect 22649 9877 22661 9911
rect 22695 9908 22707 9911
rect 23566 9908 23572 9920
rect 22695 9880 23572 9908
rect 22695 9877 22707 9880
rect 22649 9871 22707 9877
rect 23566 9868 23572 9880
rect 23624 9868 23630 9920
rect 25317 9911 25375 9917
rect 25317 9877 25329 9911
rect 25363 9908 25375 9911
rect 26970 9908 26976 9920
rect 25363 9880 26976 9908
rect 25363 9877 25375 9880
rect 25317 9871 25375 9877
rect 26970 9868 26976 9880
rect 27028 9868 27034 9920
rect 28994 9908 29000 9920
rect 28955 9880 29000 9908
rect 28994 9868 29000 9880
rect 29052 9868 29058 9920
rect 30098 9868 30104 9920
rect 30156 9908 30162 9920
rect 30193 9911 30251 9917
rect 30193 9908 30205 9911
rect 30156 9880 30205 9908
rect 30156 9868 30162 9880
rect 30193 9877 30205 9880
rect 30239 9877 30251 9911
rect 31018 9908 31024 9920
rect 30979 9880 31024 9908
rect 30193 9871 30251 9877
rect 31018 9868 31024 9880
rect 31076 9868 31082 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 7098 9664 7104 9716
rect 7156 9704 7162 9716
rect 7374 9704 7380 9716
rect 7156 9676 7380 9704
rect 7156 9664 7162 9676
rect 7374 9664 7380 9676
rect 7432 9704 7438 9716
rect 7745 9707 7803 9713
rect 7745 9704 7757 9707
rect 7432 9676 7757 9704
rect 7432 9664 7438 9676
rect 7745 9673 7757 9676
rect 7791 9673 7803 9707
rect 7745 9667 7803 9673
rect 9122 9664 9128 9716
rect 9180 9704 9186 9716
rect 12066 9704 12072 9716
rect 9180 9676 12072 9704
rect 9180 9664 9186 9676
rect 12066 9664 12072 9676
rect 12124 9664 12130 9716
rect 13648 9676 14872 9704
rect 3970 9636 3976 9648
rect 3896 9608 3976 9636
rect 3896 9577 3924 9608
rect 3970 9596 3976 9608
rect 4028 9636 4034 9648
rect 9674 9636 9680 9648
rect 4028 9608 9680 9636
rect 4028 9596 4034 9608
rect 6380 9580 6408 9608
rect 9674 9596 9680 9608
rect 9732 9596 9738 9648
rect 10226 9596 10232 9648
rect 10284 9636 10290 9648
rect 10965 9639 11023 9645
rect 10965 9636 10977 9639
rect 10284 9608 10977 9636
rect 10284 9596 10290 9608
rect 10965 9605 10977 9608
rect 11011 9605 11023 9639
rect 10965 9599 11023 9605
rect 11790 9596 11796 9648
rect 11848 9636 11854 9648
rect 12897 9639 12955 9645
rect 12897 9636 12909 9639
rect 11848 9608 11893 9636
rect 11992 9608 12909 9636
rect 11848 9596 11854 9608
rect 3881 9571 3939 9577
rect 3881 9537 3893 9571
rect 3927 9537 3939 9571
rect 3881 9531 3939 9537
rect 4148 9571 4206 9577
rect 4148 9537 4160 9571
rect 4194 9568 4206 9571
rect 4614 9568 4620 9580
rect 4194 9540 4620 9568
rect 4194 9537 4206 9540
rect 4148 9531 4206 9537
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 6362 9568 6368 9580
rect 6275 9540 6368 9568
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 6632 9571 6690 9577
rect 6632 9537 6644 9571
rect 6678 9568 6690 9571
rect 8110 9568 8116 9580
rect 6678 9540 8116 9568
rect 6678 9537 6690 9540
rect 6632 9531 6690 9537
rect 8110 9528 8116 9540
rect 8168 9528 8174 9580
rect 9013 9571 9071 9577
rect 9013 9568 9025 9571
rect 8220 9540 9025 9568
rect 5258 9364 5264 9376
rect 5219 9336 5264 9364
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 5626 9324 5632 9376
rect 5684 9364 5690 9376
rect 8220 9364 8248 9540
rect 9013 9537 9025 9540
rect 9059 9537 9071 9571
rect 9013 9531 9071 9537
rect 9490 9528 9496 9580
rect 9548 9568 9554 9580
rect 10594 9568 10600 9580
rect 9548 9540 9812 9568
rect 10555 9540 10600 9568
rect 9548 9528 9554 9540
rect 8754 9500 8760 9512
rect 8715 9472 8760 9500
rect 8754 9460 8760 9472
rect 8812 9460 8818 9512
rect 9784 9432 9812 9540
rect 10594 9528 10600 9540
rect 10652 9528 10658 9580
rect 10778 9568 10784 9580
rect 10739 9540 10784 9568
rect 10778 9528 10784 9540
rect 10836 9528 10842 9580
rect 11238 9568 11244 9580
rect 11072 9540 11244 9568
rect 9858 9460 9864 9512
rect 9916 9500 9922 9512
rect 11072 9500 11100 9540
rect 11238 9528 11244 9540
rect 11296 9568 11302 9580
rect 11992 9577 12020 9608
rect 12897 9605 12909 9608
rect 12943 9636 12955 9639
rect 13648 9636 13676 9676
rect 14844 9648 14872 9676
rect 24302 9664 24308 9716
rect 24360 9704 24366 9716
rect 25314 9704 25320 9716
rect 24360 9676 25320 9704
rect 24360 9664 24366 9676
rect 25314 9664 25320 9676
rect 25372 9664 25378 9716
rect 25406 9664 25412 9716
rect 25464 9704 25470 9716
rect 25501 9707 25559 9713
rect 25501 9704 25513 9707
rect 25464 9676 25513 9704
rect 25464 9664 25470 9676
rect 25501 9673 25513 9676
rect 25547 9673 25559 9707
rect 25501 9667 25559 9673
rect 26878 9664 26884 9716
rect 26936 9704 26942 9716
rect 26973 9707 27031 9713
rect 26973 9704 26985 9707
rect 26936 9676 26985 9704
rect 26936 9664 26942 9676
rect 26973 9673 26985 9676
rect 27019 9673 27031 9707
rect 26973 9667 27031 9673
rect 27154 9664 27160 9716
rect 27212 9704 27218 9716
rect 32490 9704 32496 9716
rect 27212 9676 32496 9704
rect 27212 9664 27218 9676
rect 32490 9664 32496 9676
rect 32548 9664 32554 9716
rect 12943 9608 13676 9636
rect 12943 9605 12955 9608
rect 12897 9599 12955 9605
rect 13722 9596 13728 9648
rect 13780 9636 13786 9648
rect 14277 9639 14335 9645
rect 14277 9636 14289 9639
rect 13780 9608 14289 9636
rect 13780 9596 13786 9608
rect 14277 9605 14289 9608
rect 14323 9605 14335 9639
rect 14826 9636 14832 9648
rect 14739 9608 14832 9636
rect 14277 9599 14335 9605
rect 14826 9596 14832 9608
rect 14884 9636 14890 9648
rect 17678 9636 17684 9648
rect 14884 9608 17684 9636
rect 14884 9596 14890 9608
rect 17678 9596 17684 9608
rect 17736 9596 17742 9648
rect 18049 9639 18107 9645
rect 18049 9605 18061 9639
rect 18095 9636 18107 9639
rect 19334 9636 19340 9648
rect 18095 9608 19340 9636
rect 18095 9605 18107 9608
rect 18049 9599 18107 9605
rect 19334 9596 19340 9608
rect 19392 9596 19398 9648
rect 19426 9596 19432 9648
rect 19484 9636 19490 9648
rect 20162 9636 20168 9648
rect 19484 9608 20168 9636
rect 19484 9596 19490 9608
rect 20162 9596 20168 9608
rect 20220 9596 20226 9648
rect 20530 9636 20536 9648
rect 20272 9608 20536 9636
rect 11609 9571 11667 9577
rect 11609 9568 11621 9571
rect 11296 9540 11621 9568
rect 11296 9528 11302 9540
rect 11609 9537 11621 9540
rect 11655 9537 11667 9571
rect 11885 9571 11943 9577
rect 11885 9568 11897 9571
rect 11609 9531 11667 9537
rect 11716 9540 11897 9568
rect 9916 9472 11100 9500
rect 9916 9460 9922 9472
rect 11146 9460 11152 9512
rect 11204 9500 11210 9512
rect 11716 9500 11744 9540
rect 11885 9537 11897 9540
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 11977 9571 12035 9577
rect 11977 9537 11989 9571
rect 12023 9537 12035 9571
rect 12710 9568 12716 9580
rect 12671 9540 12716 9568
rect 11977 9531 12035 9537
rect 12710 9528 12716 9540
rect 12768 9528 12774 9580
rect 14090 9568 14096 9580
rect 14051 9540 14096 9568
rect 14090 9528 14096 9540
rect 14148 9528 14154 9580
rect 15286 9568 15292 9580
rect 15247 9540 15292 9568
rect 15286 9528 15292 9540
rect 15344 9528 15350 9580
rect 16390 9528 16396 9580
rect 16448 9568 16454 9580
rect 17865 9571 17923 9577
rect 17865 9568 17877 9571
rect 16448 9540 17877 9568
rect 16448 9528 16454 9540
rect 17865 9537 17877 9540
rect 17911 9568 17923 9571
rect 17954 9568 17960 9580
rect 17911 9540 17960 9568
rect 17911 9537 17923 9540
rect 17865 9531 17923 9537
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 18141 9571 18199 9577
rect 18141 9537 18153 9571
rect 18187 9568 18199 9571
rect 18230 9568 18236 9580
rect 18187 9540 18236 9568
rect 18187 9537 18199 9540
rect 18141 9531 18199 9537
rect 18230 9528 18236 9540
rect 18288 9528 18294 9580
rect 18598 9528 18604 9580
rect 18656 9568 18662 9580
rect 18693 9571 18751 9577
rect 18693 9568 18705 9571
rect 18656 9540 18705 9568
rect 18656 9528 18662 9540
rect 18693 9537 18705 9540
rect 18739 9537 18751 9571
rect 18693 9531 18751 9537
rect 18782 9528 18788 9580
rect 18840 9568 18846 9580
rect 19794 9568 19800 9580
rect 18840 9540 19800 9568
rect 18840 9528 18846 9540
rect 19794 9528 19800 9540
rect 19852 9528 19858 9580
rect 20272 9577 20300 9608
rect 20530 9596 20536 9608
rect 20588 9596 20594 9648
rect 20714 9596 20720 9648
rect 20772 9636 20778 9648
rect 23385 9639 23443 9645
rect 20772 9608 22600 9636
rect 20772 9596 20778 9608
rect 20257 9571 20315 9577
rect 20257 9537 20269 9571
rect 20303 9537 20315 9571
rect 20257 9531 20315 9537
rect 20346 9528 20352 9580
rect 20404 9568 20410 9580
rect 20625 9571 20683 9577
rect 20404 9540 20449 9568
rect 20404 9528 20410 9540
rect 20625 9537 20637 9571
rect 20671 9568 20683 9571
rect 21174 9568 21180 9580
rect 20671 9540 21180 9568
rect 20671 9537 20683 9540
rect 20625 9531 20683 9537
rect 21174 9528 21180 9540
rect 21232 9528 21238 9580
rect 21266 9528 21272 9580
rect 21324 9568 21330 9580
rect 22462 9568 22468 9580
rect 21324 9540 21369 9568
rect 22423 9540 22468 9568
rect 21324 9528 21330 9540
rect 22462 9528 22468 9540
rect 22520 9528 22526 9580
rect 22572 9577 22600 9608
rect 23385 9605 23397 9639
rect 23431 9636 23443 9639
rect 23474 9636 23480 9648
rect 23431 9608 23480 9636
rect 23431 9605 23443 9608
rect 23385 9599 23443 9605
rect 23474 9596 23480 9608
rect 23532 9596 23538 9648
rect 23569 9639 23627 9645
rect 23569 9605 23581 9639
rect 23615 9636 23627 9639
rect 24394 9636 24400 9648
rect 23615 9608 24400 9636
rect 23615 9605 23627 9608
rect 23569 9599 23627 9605
rect 24394 9596 24400 9608
rect 24452 9596 24458 9648
rect 24854 9596 24860 9648
rect 24912 9636 24918 9648
rect 25133 9639 25191 9645
rect 25133 9636 25145 9639
rect 24912 9608 25145 9636
rect 24912 9596 24918 9608
rect 25133 9605 25145 9608
rect 25179 9605 25191 9639
rect 25133 9599 25191 9605
rect 25225 9639 25283 9645
rect 25225 9605 25237 9639
rect 25271 9636 25283 9639
rect 25271 9608 27614 9636
rect 25271 9605 25283 9608
rect 25225 9599 25283 9605
rect 22557 9571 22615 9577
rect 22557 9537 22569 9571
rect 22603 9537 22615 9571
rect 22830 9568 22836 9580
rect 22791 9540 22836 9568
rect 22557 9531 22615 9537
rect 22830 9528 22836 9540
rect 22888 9528 22894 9580
rect 24213 9571 24271 9577
rect 24213 9537 24225 9571
rect 24259 9568 24271 9571
rect 24486 9568 24492 9580
rect 24259 9540 24492 9568
rect 24259 9537 24271 9540
rect 24213 9531 24271 9537
rect 24486 9528 24492 9540
rect 24544 9528 24550 9580
rect 24762 9528 24768 9580
rect 24820 9568 24826 9580
rect 24949 9571 25007 9577
rect 24949 9568 24961 9571
rect 24820 9540 24961 9568
rect 24820 9528 24826 9540
rect 24949 9537 24961 9540
rect 24995 9537 25007 9571
rect 25314 9568 25320 9580
rect 25275 9540 25320 9568
rect 24949 9531 25007 9537
rect 25286 9528 25320 9540
rect 25372 9528 25378 9580
rect 26050 9528 26056 9580
rect 26108 9568 26114 9580
rect 26145 9571 26203 9577
rect 26145 9568 26157 9571
rect 26108 9540 26157 9568
rect 26108 9528 26114 9540
rect 26145 9537 26157 9540
rect 26191 9537 26203 9571
rect 26145 9531 26203 9537
rect 26970 9528 26976 9580
rect 27028 9568 27034 9580
rect 27157 9571 27215 9577
rect 27157 9568 27169 9571
rect 27028 9540 27169 9568
rect 27028 9528 27034 9540
rect 27157 9537 27169 9540
rect 27203 9537 27215 9571
rect 27157 9531 27215 9537
rect 11204 9472 11744 9500
rect 11204 9460 11210 9472
rect 13722 9460 13728 9512
rect 13780 9500 13786 9512
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 13780 9472 13921 9500
rect 13780 9460 13786 9472
rect 13909 9469 13921 9472
rect 13955 9469 13967 9503
rect 15565 9503 15623 9509
rect 15565 9500 15577 9503
rect 13909 9463 13967 9469
rect 15089 9472 15577 9500
rect 11790 9432 11796 9444
rect 9784 9404 11796 9432
rect 11790 9392 11796 9404
rect 11848 9392 11854 9444
rect 12161 9435 12219 9441
rect 12161 9401 12173 9435
rect 12207 9432 12219 9435
rect 12618 9432 12624 9444
rect 12207 9404 12624 9432
rect 12207 9401 12219 9404
rect 12161 9395 12219 9401
rect 12618 9392 12624 9404
rect 12676 9392 12682 9444
rect 5684 9336 8248 9364
rect 10137 9367 10195 9373
rect 5684 9324 5690 9336
rect 10137 9333 10149 9367
rect 10183 9364 10195 9367
rect 10226 9364 10232 9376
rect 10183 9336 10232 9364
rect 10183 9333 10195 9336
rect 10137 9327 10195 9333
rect 10226 9324 10232 9336
rect 10284 9324 10290 9376
rect 11238 9324 11244 9376
rect 11296 9364 11302 9376
rect 15089 9364 15117 9472
rect 15565 9469 15577 9472
rect 15611 9469 15623 9503
rect 16666 9500 16672 9512
rect 16579 9472 16672 9500
rect 15565 9463 15623 9469
rect 15580 9432 15608 9463
rect 16666 9460 16672 9472
rect 16724 9500 16730 9512
rect 18969 9503 19027 9509
rect 18969 9500 18981 9503
rect 16724 9472 18981 9500
rect 16724 9460 16730 9472
rect 18969 9469 18981 9472
rect 19015 9500 19027 9503
rect 19015 9472 21220 9500
rect 19015 9469 19027 9472
rect 18969 9463 19027 9469
rect 16942 9432 16948 9444
rect 15580 9404 16948 9432
rect 16942 9392 16948 9404
rect 17000 9392 17006 9444
rect 17037 9435 17095 9441
rect 17037 9401 17049 9435
rect 17083 9432 17095 9435
rect 17954 9432 17960 9444
rect 17083 9404 17960 9432
rect 17083 9401 17095 9404
rect 17037 9395 17095 9401
rect 17954 9392 17960 9404
rect 18012 9432 18018 9444
rect 18690 9432 18696 9444
rect 18012 9404 18696 9432
rect 18012 9392 18018 9404
rect 18690 9392 18696 9404
rect 18748 9392 18754 9444
rect 18984 9404 20300 9432
rect 18984 9376 19012 9404
rect 11296 9336 15117 9364
rect 11296 9324 11302 9336
rect 15654 9324 15660 9376
rect 15712 9364 15718 9376
rect 17129 9367 17187 9373
rect 17129 9364 17141 9367
rect 15712 9336 17141 9364
rect 15712 9324 15718 9336
rect 17129 9333 17141 9336
rect 17175 9333 17187 9367
rect 17129 9327 17187 9333
rect 17586 9324 17592 9376
rect 17644 9364 17650 9376
rect 17865 9367 17923 9373
rect 17865 9364 17877 9367
rect 17644 9336 17877 9364
rect 17644 9324 17650 9336
rect 17865 9333 17877 9336
rect 17911 9333 17923 9367
rect 18966 9364 18972 9376
rect 18927 9336 18972 9364
rect 17865 9327 17923 9333
rect 18966 9324 18972 9336
rect 19024 9324 19030 9376
rect 19242 9364 19248 9376
rect 19203 9336 19248 9364
rect 19242 9324 19248 9336
rect 19300 9324 19306 9376
rect 20070 9364 20076 9376
rect 20031 9336 20076 9364
rect 20070 9324 20076 9336
rect 20128 9324 20134 9376
rect 20272 9364 20300 9404
rect 20714 9392 20720 9444
rect 20772 9432 20778 9444
rect 21085 9435 21143 9441
rect 21085 9432 21097 9435
rect 20772 9404 21097 9432
rect 20772 9392 20778 9404
rect 21085 9401 21097 9404
rect 21131 9401 21143 9435
rect 21192 9432 21220 9472
rect 22094 9460 22100 9512
rect 22152 9500 22158 9512
rect 24029 9503 24087 9509
rect 24029 9500 24041 9503
rect 22152 9472 24041 9500
rect 22152 9460 22158 9472
rect 24029 9469 24041 9472
rect 24075 9469 24087 9503
rect 24029 9463 24087 9469
rect 24397 9503 24455 9509
rect 24397 9469 24409 9503
rect 24443 9500 24455 9503
rect 24670 9500 24676 9512
rect 24443 9472 24676 9500
rect 24443 9469 24455 9472
rect 24397 9463 24455 9469
rect 22186 9432 22192 9444
rect 21192 9404 22192 9432
rect 21085 9395 21143 9401
rect 22186 9392 22192 9404
rect 22244 9392 22250 9444
rect 22281 9435 22339 9441
rect 22281 9401 22293 9435
rect 22327 9432 22339 9435
rect 22922 9432 22928 9444
rect 22327 9404 22928 9432
rect 22327 9401 22339 9404
rect 22281 9395 22339 9401
rect 22922 9392 22928 9404
rect 22980 9392 22986 9444
rect 24044 9432 24072 9463
rect 24670 9460 24676 9472
rect 24728 9460 24734 9512
rect 25286 9500 25314 9528
rect 26694 9500 26700 9512
rect 25286 9472 26700 9500
rect 26694 9460 26700 9472
rect 26752 9460 26758 9512
rect 27586 9500 27614 9608
rect 27982 9596 27988 9648
rect 28040 9636 28046 9648
rect 28169 9639 28227 9645
rect 28169 9636 28181 9639
rect 28040 9608 28181 9636
rect 28040 9596 28046 9608
rect 28169 9605 28181 9608
rect 28215 9605 28227 9639
rect 28994 9636 29000 9648
rect 28169 9599 28227 9605
rect 28368 9608 29000 9636
rect 27890 9568 27896 9580
rect 27851 9540 27896 9568
rect 27890 9528 27896 9540
rect 27948 9528 27954 9580
rect 28074 9568 28080 9580
rect 28035 9540 28080 9568
rect 28074 9528 28080 9540
rect 28132 9528 28138 9580
rect 28368 9577 28396 9608
rect 28994 9596 29000 9608
rect 29052 9596 29058 9648
rect 28353 9571 28411 9577
rect 28353 9537 28365 9571
rect 28399 9537 28411 9571
rect 28626 9568 28632 9580
rect 28587 9540 28632 9568
rect 28353 9531 28411 9537
rect 28626 9528 28632 9540
rect 28684 9528 28690 9580
rect 29270 9568 29276 9580
rect 29231 9540 29276 9568
rect 29270 9528 29276 9540
rect 29328 9528 29334 9580
rect 29362 9528 29368 9580
rect 29420 9568 29426 9580
rect 29917 9571 29975 9577
rect 29917 9568 29929 9571
rect 29420 9540 29929 9568
rect 29420 9528 29426 9540
rect 29917 9537 29929 9540
rect 29963 9537 29975 9571
rect 29917 9531 29975 9537
rect 30561 9571 30619 9577
rect 30561 9537 30573 9571
rect 30607 9568 30619 9571
rect 30926 9568 30932 9580
rect 30607 9540 30932 9568
rect 30607 9537 30619 9540
rect 30561 9531 30619 9537
rect 30926 9528 30932 9540
rect 30984 9528 30990 9580
rect 31202 9568 31208 9580
rect 31163 9540 31208 9568
rect 31202 9528 31208 9540
rect 31260 9528 31266 9580
rect 27586 9472 30420 9500
rect 24946 9432 24952 9444
rect 24044 9404 24952 9432
rect 24946 9392 24952 9404
rect 25004 9432 25010 9444
rect 25130 9432 25136 9444
rect 25004 9404 25136 9432
rect 25004 9392 25010 9404
rect 25130 9392 25136 9404
rect 25188 9392 25194 9444
rect 25590 9392 25596 9444
rect 25648 9432 25654 9444
rect 30392 9441 30420 9472
rect 29089 9435 29147 9441
rect 29089 9432 29101 9435
rect 25648 9404 29101 9432
rect 25648 9392 25654 9404
rect 29089 9401 29101 9404
rect 29135 9401 29147 9435
rect 29089 9395 29147 9401
rect 30377 9435 30435 9441
rect 30377 9401 30389 9435
rect 30423 9401 30435 9435
rect 30377 9395 30435 9401
rect 20533 9367 20591 9373
rect 20533 9364 20545 9367
rect 20272 9336 20545 9364
rect 20533 9333 20545 9336
rect 20579 9364 20591 9367
rect 21358 9364 21364 9376
rect 20579 9336 21364 9364
rect 20579 9333 20591 9336
rect 20533 9327 20591 9333
rect 21358 9324 21364 9336
rect 21416 9324 21422 9376
rect 22738 9364 22744 9376
rect 22699 9336 22744 9364
rect 22738 9324 22744 9336
rect 22796 9324 22802 9376
rect 23934 9324 23940 9376
rect 23992 9364 23998 9376
rect 25498 9364 25504 9376
rect 23992 9336 25504 9364
rect 23992 9324 23998 9336
rect 25498 9324 25504 9336
rect 25556 9324 25562 9376
rect 25958 9364 25964 9376
rect 25919 9336 25964 9364
rect 25958 9324 25964 9336
rect 26016 9324 26022 9376
rect 26050 9324 26056 9376
rect 26108 9364 26114 9376
rect 29733 9367 29791 9373
rect 29733 9364 29745 9367
rect 26108 9336 29745 9364
rect 26108 9324 26114 9336
rect 29733 9333 29745 9336
rect 29779 9333 29791 9367
rect 29733 9327 29791 9333
rect 30742 9324 30748 9376
rect 30800 9364 30806 9376
rect 31021 9367 31079 9373
rect 31021 9364 31033 9367
rect 30800 9336 31033 9364
rect 30800 9324 30806 9336
rect 31021 9333 31033 9336
rect 31067 9333 31079 9367
rect 31021 9327 31079 9333
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 6917 9163 6975 9169
rect 6917 9129 6929 9163
rect 6963 9160 6975 9163
rect 7190 9160 7196 9172
rect 6963 9132 7196 9160
rect 6963 9129 6975 9132
rect 6917 9123 6975 9129
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 8018 9160 8024 9172
rect 7979 9132 8024 9160
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 8128 9132 13676 9160
rect 8128 9092 8156 9132
rect 3252 9064 8156 9092
rect 13648 9092 13676 9132
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 18690 9160 18696 9172
rect 13780 9132 18276 9160
rect 18651 9132 18696 9160
rect 13780 9120 13786 9132
rect 16206 9092 16212 9104
rect 13648 9064 16212 9092
rect 3252 8965 3280 9064
rect 16206 9052 16212 9064
rect 16264 9052 16270 9104
rect 17310 9092 17316 9104
rect 16500 9064 17316 9092
rect 6270 9024 6276 9036
rect 4540 8996 6276 9024
rect 4540 8965 4568 8996
rect 6270 8984 6276 8996
rect 6328 8984 6334 9036
rect 7558 9024 7564 9036
rect 6748 8996 7564 9024
rect 3237 8959 3295 8965
rect 3237 8925 3249 8959
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 4525 8959 4583 8965
rect 4525 8925 4537 8959
rect 4571 8925 4583 8959
rect 4525 8919 4583 8925
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8956 5227 8959
rect 5258 8956 5264 8968
rect 5215 8928 5264 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 2130 8848 2136 8900
rect 2188 8888 2194 8900
rect 5184 8888 5212 8919
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 5350 8916 5356 8968
rect 5408 8956 5414 8968
rect 5534 8956 5540 8968
rect 5408 8928 5453 8956
rect 5495 8928 5540 8956
rect 5408 8916 5414 8928
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 5810 8956 5816 8968
rect 5771 8928 5816 8956
rect 5810 8916 5816 8928
rect 5868 8916 5874 8968
rect 5902 8916 5908 8968
rect 5960 8956 5966 8968
rect 6748 8965 6776 8996
rect 7558 8984 7564 8996
rect 7616 9024 7622 9036
rect 9217 9027 9275 9033
rect 9217 9024 9229 9027
rect 7616 8996 9229 9024
rect 7616 8984 7622 8996
rect 6365 8959 6423 8965
rect 5960 8928 6005 8956
rect 5960 8916 5966 8928
rect 6365 8925 6377 8959
rect 6411 8925 6423 8959
rect 6641 8959 6699 8965
rect 6641 8956 6653 8959
rect 6365 8919 6423 8925
rect 6472 8928 6653 8956
rect 6380 8888 6408 8919
rect 2188 8860 5120 8888
rect 5184 8860 6408 8888
rect 2188 8848 2194 8860
rect 3053 8823 3111 8829
rect 3053 8789 3065 8823
rect 3099 8820 3111 8823
rect 3142 8820 3148 8832
rect 3099 8792 3148 8820
rect 3099 8789 3111 8792
rect 3053 8783 3111 8789
rect 3142 8780 3148 8792
rect 3200 8780 3206 8832
rect 4341 8823 4399 8829
rect 4341 8789 4353 8823
rect 4387 8820 4399 8823
rect 4982 8820 4988 8832
rect 4387 8792 4988 8820
rect 4387 8789 4399 8792
rect 4341 8783 4399 8789
rect 4982 8780 4988 8792
rect 5040 8780 5046 8832
rect 5092 8820 5120 8860
rect 6472 8820 6500 8928
rect 6641 8925 6653 8928
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 6733 8959 6791 8965
rect 6733 8925 6745 8959
rect 6779 8925 6791 8959
rect 7466 8956 7472 8968
rect 7427 8928 7472 8956
rect 6733 8919 6791 8925
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 7852 8965 7880 8996
rect 9217 8993 9229 8996
rect 9263 8993 9275 9027
rect 14274 9024 14280 9036
rect 9217 8987 9275 8993
rect 13648 8996 14280 9024
rect 7837 8959 7895 8965
rect 7837 8925 7849 8959
rect 7883 8925 7895 8959
rect 7837 8919 7895 8925
rect 8570 8916 8576 8968
rect 8628 8956 8634 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8628 8928 8953 8956
rect 8628 8916 8634 8928
rect 8941 8925 8953 8928
rect 8987 8956 8999 8959
rect 10042 8956 10048 8968
rect 8987 8928 10048 8956
rect 8987 8925 8999 8928
rect 8941 8919 8999 8925
rect 10042 8916 10048 8928
rect 10100 8916 10106 8968
rect 10321 8959 10379 8965
rect 10321 8925 10333 8959
rect 10367 8956 10379 8959
rect 10962 8956 10968 8968
rect 10367 8928 10968 8956
rect 10367 8925 10379 8928
rect 10321 8919 10379 8925
rect 10962 8916 10968 8928
rect 11020 8956 11026 8968
rect 12161 8959 12219 8965
rect 12161 8956 12173 8959
rect 11020 8928 12173 8956
rect 11020 8916 11026 8928
rect 12161 8925 12173 8928
rect 12207 8925 12219 8959
rect 13648 8956 13676 8996
rect 14274 8984 14280 8996
rect 14332 8984 14338 9036
rect 12161 8919 12219 8925
rect 12268 8928 13676 8956
rect 6549 8891 6607 8897
rect 6549 8857 6561 8891
rect 6595 8857 6607 8891
rect 6549 8851 6607 8857
rect 5092 8792 6500 8820
rect 6564 8820 6592 8851
rect 7282 8848 7288 8900
rect 7340 8888 7346 8900
rect 7653 8891 7711 8897
rect 7653 8888 7665 8891
rect 7340 8860 7665 8888
rect 7340 8848 7346 8860
rect 7653 8857 7665 8860
rect 7699 8857 7711 8891
rect 7653 8851 7711 8857
rect 7745 8891 7803 8897
rect 7745 8857 7757 8891
rect 7791 8888 7803 8891
rect 7791 8860 7880 8888
rect 7791 8857 7803 8860
rect 7745 8851 7803 8857
rect 7300 8820 7328 8848
rect 7852 8832 7880 8860
rect 9030 8848 9036 8900
rect 9088 8888 9094 8900
rect 9398 8888 9404 8900
rect 9088 8860 9404 8888
rect 9088 8848 9094 8860
rect 9398 8848 9404 8860
rect 9456 8848 9462 8900
rect 10134 8848 10140 8900
rect 10192 8888 10198 8900
rect 10566 8891 10624 8897
rect 10566 8888 10578 8891
rect 10192 8860 10578 8888
rect 10192 8848 10198 8860
rect 10566 8857 10578 8860
rect 10612 8857 10624 8891
rect 12268 8888 12296 8928
rect 13722 8916 13728 8968
rect 13780 8956 13786 8968
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 13780 8928 14105 8956
rect 13780 8916 13786 8928
rect 14093 8925 14105 8928
rect 14139 8925 14151 8959
rect 15102 8956 15108 8968
rect 15063 8928 15108 8956
rect 14093 8919 14151 8925
rect 15102 8916 15108 8928
rect 15160 8916 15166 8968
rect 15286 8916 15292 8968
rect 15344 8956 15350 8968
rect 16500 8965 16528 9064
rect 17310 9052 17316 9064
rect 17368 9052 17374 9104
rect 18248 9092 18276 9132
rect 18690 9120 18696 9132
rect 18748 9120 18754 9172
rect 21174 9160 21180 9172
rect 18800 9132 20760 9160
rect 21135 9132 21180 9160
rect 18800 9092 18828 9132
rect 18248 9064 18828 9092
rect 20732 9092 20760 9132
rect 21174 9120 21180 9132
rect 21232 9120 21238 9172
rect 21358 9120 21364 9172
rect 21416 9160 21422 9172
rect 22278 9160 22284 9172
rect 21416 9132 22284 9160
rect 21416 9120 21422 9132
rect 22278 9120 22284 9132
rect 22336 9160 22342 9172
rect 22738 9160 22744 9172
rect 22336 9132 22744 9160
rect 22336 9120 22342 9132
rect 22738 9120 22744 9132
rect 22796 9120 22802 9172
rect 22830 9120 22836 9172
rect 22888 9160 22894 9172
rect 23477 9163 23535 9169
rect 23477 9160 23489 9163
rect 22888 9132 23489 9160
rect 22888 9120 22894 9132
rect 23477 9129 23489 9132
rect 23523 9129 23535 9163
rect 23477 9123 23535 9129
rect 23750 9120 23756 9172
rect 23808 9160 23814 9172
rect 29825 9163 29883 9169
rect 29825 9160 29837 9163
rect 23808 9132 29837 9160
rect 23808 9120 23814 9132
rect 29825 9129 29837 9132
rect 29871 9160 29883 9163
rect 32766 9160 32772 9172
rect 29871 9132 32772 9160
rect 29871 9129 29883 9132
rect 29825 9123 29883 9129
rect 32766 9120 32772 9132
rect 32824 9120 32830 9172
rect 21910 9092 21916 9104
rect 20732 9064 21916 9092
rect 21910 9052 21916 9064
rect 21968 9052 21974 9104
rect 25498 9052 25504 9104
rect 25556 9092 25562 9104
rect 25777 9095 25835 9101
rect 25777 9092 25789 9095
rect 25556 9064 25789 9092
rect 25556 9052 25562 9064
rect 25777 9061 25789 9064
rect 25823 9061 25835 9095
rect 25777 9055 25835 9061
rect 26234 9052 26240 9104
rect 26292 9092 26298 9104
rect 31021 9095 31079 9101
rect 31021 9092 31033 9095
rect 26292 9064 31033 9092
rect 26292 9052 26298 9064
rect 31021 9061 31033 9064
rect 31067 9061 31079 9095
rect 31021 9055 31079 9061
rect 16666 9024 16672 9036
rect 16627 8996 16672 9024
rect 16666 8984 16672 8996
rect 16724 8984 16730 9036
rect 24394 9024 24400 9036
rect 24355 8996 24400 9024
rect 24394 8984 24400 8996
rect 24452 8984 24458 9036
rect 29178 9024 29184 9036
rect 26160 8996 29184 9024
rect 15381 8959 15439 8965
rect 15381 8956 15393 8959
rect 15344 8928 15393 8956
rect 15344 8916 15350 8928
rect 15381 8925 15393 8928
rect 15427 8925 15439 8959
rect 15381 8919 15439 8925
rect 16485 8959 16543 8965
rect 16485 8925 16497 8959
rect 16531 8956 16543 8959
rect 16574 8956 16580 8968
rect 16531 8928 16580 8956
rect 16531 8925 16543 8928
rect 16485 8919 16543 8925
rect 16574 8916 16580 8928
rect 16632 8916 16638 8968
rect 16761 8959 16819 8965
rect 16761 8925 16773 8959
rect 16807 8956 16819 8959
rect 17126 8956 17132 8968
rect 16807 8928 17132 8956
rect 16807 8925 16819 8928
rect 16761 8919 16819 8925
rect 17126 8916 17132 8928
rect 17184 8916 17190 8968
rect 17313 8959 17371 8965
rect 17313 8925 17325 8959
rect 17359 8956 17371 8959
rect 17862 8956 17868 8968
rect 17359 8928 17868 8956
rect 17359 8925 17371 8928
rect 17313 8919 17371 8925
rect 17862 8916 17868 8928
rect 17920 8916 17926 8968
rect 19797 8959 19855 8965
rect 19797 8925 19809 8959
rect 19843 8956 19855 8959
rect 20622 8956 20628 8968
rect 19843 8928 20628 8956
rect 19843 8925 19855 8928
rect 19797 8919 19855 8925
rect 20622 8916 20628 8928
rect 20680 8956 20686 8968
rect 22097 8959 22155 8965
rect 22097 8956 22109 8959
rect 20680 8928 22109 8956
rect 20680 8916 20686 8928
rect 22097 8925 22109 8928
rect 22143 8956 22155 8959
rect 24412 8956 24440 8984
rect 22143 8928 24440 8956
rect 24664 8959 24722 8965
rect 22143 8925 22155 8928
rect 22097 8919 22155 8925
rect 24664 8925 24676 8959
rect 24710 8956 24722 8959
rect 25958 8956 25964 8968
rect 24710 8928 25964 8956
rect 24710 8925 24722 8928
rect 24664 8919 24722 8925
rect 25958 8916 25964 8928
rect 26016 8916 26022 8968
rect 10566 8851 10624 8857
rect 11256 8860 12296 8888
rect 12428 8891 12486 8897
rect 6564 8792 7328 8820
rect 7834 8780 7840 8832
rect 7892 8780 7898 8832
rect 8478 8780 8484 8832
rect 8536 8820 8542 8832
rect 11256 8820 11284 8860
rect 12428 8857 12440 8891
rect 12474 8888 12486 8891
rect 12526 8888 12532 8900
rect 12474 8860 12532 8888
rect 12474 8857 12486 8860
rect 12428 8851 12486 8857
rect 12526 8848 12532 8860
rect 12584 8848 12590 8900
rect 16390 8888 16396 8900
rect 13280 8860 16396 8888
rect 8536 8792 11284 8820
rect 8536 8780 8542 8792
rect 11330 8780 11336 8832
rect 11388 8820 11394 8832
rect 11701 8823 11759 8829
rect 11701 8820 11713 8823
rect 11388 8792 11713 8820
rect 11388 8780 11394 8792
rect 11701 8789 11713 8792
rect 11747 8789 11759 8823
rect 11701 8783 11759 8789
rect 11790 8780 11796 8832
rect 11848 8820 11854 8832
rect 13280 8820 13308 8860
rect 11848 8792 13308 8820
rect 11848 8780 11854 8792
rect 13354 8780 13360 8832
rect 13412 8820 13418 8832
rect 14292 8829 14320 8860
rect 16390 8848 16396 8860
rect 16448 8848 16454 8900
rect 16666 8848 16672 8900
rect 16724 8888 16730 8900
rect 17586 8897 17592 8900
rect 16853 8891 16911 8897
rect 16853 8888 16865 8891
rect 16724 8860 16865 8888
rect 16724 8848 16730 8860
rect 16853 8857 16865 8860
rect 16899 8857 16911 8891
rect 17580 8888 17592 8897
rect 17547 8860 17592 8888
rect 16853 8851 16911 8857
rect 17580 8851 17592 8860
rect 17586 8848 17592 8851
rect 17644 8848 17650 8900
rect 17678 8848 17684 8900
rect 17736 8888 17742 8900
rect 20064 8891 20122 8897
rect 17736 8860 20024 8888
rect 17736 8848 17742 8860
rect 13541 8823 13599 8829
rect 13541 8820 13553 8823
rect 13412 8792 13553 8820
rect 13412 8780 13418 8792
rect 13541 8789 13553 8792
rect 13587 8789 13599 8823
rect 13541 8783 13599 8789
rect 14277 8823 14335 8829
rect 14277 8789 14289 8823
rect 14323 8789 14335 8823
rect 14918 8820 14924 8832
rect 14879 8792 14924 8820
rect 14277 8783 14335 8789
rect 14918 8780 14924 8792
rect 14976 8780 14982 8832
rect 15289 8823 15347 8829
rect 15289 8789 15301 8823
rect 15335 8820 15347 8823
rect 17954 8820 17960 8832
rect 15335 8792 17960 8820
rect 15335 8789 15347 8792
rect 15289 8783 15347 8789
rect 17954 8780 17960 8792
rect 18012 8780 18018 8832
rect 19996 8820 20024 8860
rect 20064 8857 20076 8891
rect 20110 8888 20122 8891
rect 21818 8888 21824 8900
rect 20110 8860 21824 8888
rect 20110 8857 20122 8860
rect 20064 8851 20122 8857
rect 21818 8848 21824 8860
rect 21876 8848 21882 8900
rect 22364 8891 22422 8897
rect 22364 8857 22376 8891
rect 22410 8888 22422 8891
rect 26160 8888 26188 8996
rect 29178 8984 29184 8996
rect 29236 8984 29242 9036
rect 26237 8959 26295 8965
rect 26237 8925 26249 8959
rect 26283 8956 26295 8959
rect 26326 8956 26332 8968
rect 26283 8928 26332 8956
rect 26283 8925 26295 8928
rect 26237 8919 26295 8925
rect 26326 8916 26332 8928
rect 26384 8916 26390 8968
rect 26602 8956 26608 8968
rect 26563 8928 26608 8956
rect 26602 8916 26608 8928
rect 26660 8916 26666 8968
rect 26694 8916 26700 8968
rect 26752 8956 26758 8968
rect 27338 8956 27344 8968
rect 26752 8928 27344 8956
rect 26752 8916 26758 8928
rect 27338 8916 27344 8928
rect 27396 8916 27402 8968
rect 27798 8956 27804 8968
rect 27759 8928 27804 8956
rect 27798 8916 27804 8928
rect 27856 8916 27862 8968
rect 28074 8956 28080 8968
rect 28035 8928 28080 8956
rect 28074 8916 28080 8928
rect 28132 8916 28138 8968
rect 28350 8956 28356 8968
rect 28311 8928 28356 8956
rect 28350 8916 28356 8928
rect 28408 8916 28414 8968
rect 28626 8956 28632 8968
rect 28539 8928 28632 8956
rect 28626 8916 28632 8928
rect 28684 8956 28690 8968
rect 29641 8959 29699 8965
rect 29641 8956 29653 8959
rect 28684 8928 29653 8956
rect 28684 8916 28690 8928
rect 29641 8925 29653 8928
rect 29687 8956 29699 8959
rect 30190 8956 30196 8968
rect 29687 8928 30196 8956
rect 29687 8925 29699 8928
rect 29641 8919 29699 8925
rect 30190 8916 30196 8928
rect 30248 8916 30254 8968
rect 30561 8959 30619 8965
rect 30561 8925 30573 8959
rect 30607 8956 30619 8959
rect 30650 8956 30656 8968
rect 30607 8928 30656 8956
rect 30607 8925 30619 8928
rect 30561 8919 30619 8925
rect 30650 8916 30656 8928
rect 30708 8916 30714 8968
rect 31202 8956 31208 8968
rect 31163 8928 31208 8956
rect 31202 8916 31208 8928
rect 31260 8916 31266 8968
rect 31846 8956 31852 8968
rect 31807 8928 31852 8956
rect 31846 8916 31852 8928
rect 31904 8916 31910 8968
rect 22410 8860 26188 8888
rect 26421 8891 26479 8897
rect 22410 8857 22422 8860
rect 22364 8851 22422 8857
rect 26421 8857 26433 8891
rect 26467 8857 26479 8891
rect 26421 8851 26479 8857
rect 26513 8891 26571 8897
rect 26513 8857 26525 8891
rect 26559 8888 26571 8891
rect 26559 8860 28120 8888
rect 26559 8857 26571 8860
rect 26513 8851 26571 8857
rect 24302 8820 24308 8832
rect 19996 8792 24308 8820
rect 24302 8780 24308 8792
rect 24360 8780 24366 8832
rect 24854 8780 24860 8832
rect 24912 8820 24918 8832
rect 26436 8820 26464 8851
rect 24912 8792 26464 8820
rect 24912 8780 24918 8792
rect 26602 8780 26608 8832
rect 26660 8820 26666 8832
rect 26789 8823 26847 8829
rect 26789 8820 26801 8823
rect 26660 8792 26801 8820
rect 26660 8780 26666 8792
rect 26789 8789 26801 8792
rect 26835 8789 26847 8823
rect 26789 8783 26847 8789
rect 26878 8780 26884 8832
rect 26936 8820 26942 8832
rect 27430 8820 27436 8832
rect 26936 8792 27436 8820
rect 26936 8780 26942 8792
rect 27430 8780 27436 8792
rect 27488 8780 27494 8832
rect 28092 8820 28120 8860
rect 28166 8848 28172 8900
rect 28224 8888 28230 8900
rect 28224 8860 28269 8888
rect 28224 8848 28230 8860
rect 29914 8848 29920 8900
rect 29972 8888 29978 8900
rect 29972 8860 31708 8888
rect 29972 8848 29978 8860
rect 29730 8820 29736 8832
rect 28092 8792 29736 8820
rect 29730 8780 29736 8792
rect 29788 8780 29794 8832
rect 30377 8823 30435 8829
rect 30377 8789 30389 8823
rect 30423 8820 30435 8823
rect 30558 8820 30564 8832
rect 30423 8792 30564 8820
rect 30423 8789 30435 8792
rect 30377 8783 30435 8789
rect 30558 8780 30564 8792
rect 30616 8780 30622 8832
rect 31680 8829 31708 8860
rect 31665 8823 31723 8829
rect 31665 8789 31677 8823
rect 31711 8789 31723 8823
rect 31665 8783 31723 8789
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 3697 8619 3755 8625
rect 3697 8585 3709 8619
rect 3743 8585 3755 8619
rect 3697 8579 3755 8585
rect 4341 8619 4399 8625
rect 4341 8585 4353 8619
rect 4387 8616 4399 8619
rect 5166 8616 5172 8628
rect 4387 8588 5172 8616
rect 4387 8585 4399 8588
rect 4341 8579 4399 8585
rect 3712 8548 3740 8579
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 5626 8616 5632 8628
rect 5587 8588 5632 8616
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 9493 8619 9551 8625
rect 9493 8616 9505 8619
rect 5828 8588 9505 8616
rect 5718 8548 5724 8560
rect 3712 8520 5724 8548
rect 5718 8508 5724 8520
rect 5776 8508 5782 8560
rect 1302 8440 1308 8492
rect 1360 8480 1366 8492
rect 1581 8483 1639 8489
rect 1581 8480 1593 8483
rect 1360 8452 1593 8480
rect 1360 8440 1366 8452
rect 1581 8449 1593 8452
rect 1627 8449 1639 8483
rect 1581 8443 1639 8449
rect 3881 8483 3939 8489
rect 3881 8449 3893 8483
rect 3927 8480 3939 8483
rect 3970 8480 3976 8492
rect 3927 8452 3976 8480
rect 3927 8449 3939 8452
rect 3881 8443 3939 8449
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8449 4583 8483
rect 4525 8443 4583 8449
rect 4540 8412 4568 8443
rect 4890 8440 4896 8492
rect 4948 8480 4954 8492
rect 4985 8483 5043 8489
rect 4985 8480 4997 8483
rect 4948 8452 4997 8480
rect 4948 8440 4954 8452
rect 4985 8449 4997 8452
rect 5031 8449 5043 8483
rect 4985 8443 5043 8449
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8480 5227 8483
rect 5626 8480 5632 8492
rect 5215 8452 5632 8480
rect 5215 8449 5227 8452
rect 5169 8443 5227 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 5828 8489 5856 8588
rect 9493 8585 9505 8588
rect 9539 8585 9551 8619
rect 10318 8616 10324 8628
rect 10279 8588 10324 8616
rect 9493 8579 9551 8585
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 11885 8619 11943 8625
rect 11885 8616 11897 8619
rect 10980 8588 11897 8616
rect 8478 8548 8484 8560
rect 7208 8520 8484 8548
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8480 6699 8483
rect 7006 8480 7012 8492
rect 6687 8452 7012 8480
rect 6687 8449 6699 8452
rect 6641 8443 6699 8449
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8449 7159 8483
rect 7101 8443 7159 8449
rect 5074 8412 5080 8424
rect 4540 8384 4936 8412
rect 5035 8384 5080 8412
rect 1397 8279 1455 8285
rect 1397 8245 1409 8279
rect 1443 8276 1455 8279
rect 1946 8276 1952 8288
rect 1443 8248 1952 8276
rect 1443 8245 1455 8248
rect 1397 8239 1455 8245
rect 1946 8236 1952 8248
rect 2004 8236 2010 8288
rect 4908 8276 4936 8384
rect 5074 8372 5080 8384
rect 5132 8372 5138 8424
rect 5258 8372 5264 8424
rect 5316 8412 5322 8424
rect 7116 8412 7144 8443
rect 5316 8384 7144 8412
rect 5316 8372 5322 8384
rect 7208 8344 7236 8520
rect 8478 8508 8484 8520
rect 8536 8508 8542 8560
rect 9125 8551 9183 8557
rect 9125 8517 9137 8551
rect 9171 8548 9183 8551
rect 9858 8548 9864 8560
rect 9171 8520 9864 8548
rect 9171 8517 9183 8520
rect 9125 8511 9183 8517
rect 9858 8508 9864 8520
rect 9916 8508 9922 8560
rect 10870 8508 10876 8560
rect 10928 8548 10934 8560
rect 10980 8548 11008 8588
rect 11885 8585 11897 8588
rect 11931 8585 11943 8619
rect 13906 8616 13912 8628
rect 13867 8588 13912 8616
rect 11885 8579 11943 8585
rect 13906 8576 13912 8588
rect 13964 8576 13970 8628
rect 16574 8576 16580 8628
rect 16632 8576 16638 8628
rect 16666 8576 16672 8628
rect 16724 8616 16730 8628
rect 18598 8616 18604 8628
rect 16724 8588 18604 8616
rect 16724 8576 16730 8588
rect 18598 8576 18604 8588
rect 18656 8616 18662 8628
rect 19245 8619 19303 8625
rect 19245 8616 19257 8619
rect 18656 8588 19257 8616
rect 18656 8576 18662 8588
rect 19245 8585 19257 8588
rect 19291 8585 19303 8619
rect 24486 8616 24492 8628
rect 19245 8579 19303 8585
rect 19352 8588 24164 8616
rect 24447 8588 24492 8616
rect 10928 8520 11008 8548
rect 10928 8508 10934 8520
rect 11698 8508 11704 8560
rect 11756 8548 11762 8560
rect 14458 8548 14464 8560
rect 11756 8520 11801 8548
rect 12820 8520 14464 8548
rect 11756 8508 11762 8520
rect 7374 8480 7380 8492
rect 7335 8452 7380 8480
rect 7374 8440 7380 8452
rect 7432 8440 7438 8492
rect 8294 8480 8300 8492
rect 8255 8452 8300 8480
rect 8294 8440 8300 8452
rect 8352 8440 8358 8492
rect 8386 8440 8392 8492
rect 8444 8480 8450 8492
rect 9306 8480 9312 8492
rect 8444 8452 9312 8480
rect 8444 8440 8450 8452
rect 9306 8440 9312 8452
rect 9364 8440 9370 8492
rect 9490 8440 9496 8492
rect 9548 8480 9554 8492
rect 9953 8483 10011 8489
rect 9953 8480 9965 8483
rect 9548 8452 9965 8480
rect 9548 8440 9554 8452
rect 9953 8449 9965 8452
rect 9999 8449 10011 8483
rect 10134 8480 10140 8492
rect 10095 8452 10140 8480
rect 9953 8443 10011 8449
rect 10134 8440 10140 8452
rect 10192 8440 10198 8492
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8449 10839 8483
rect 10781 8443 10839 8449
rect 10965 8483 11023 8489
rect 10965 8449 10977 8483
rect 11011 8480 11023 8483
rect 11238 8480 11244 8492
rect 11011 8452 11244 8480
rect 11011 8449 11023 8452
rect 10965 8443 11023 8449
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8412 7343 8415
rect 9766 8412 9772 8424
rect 7331 8384 9772 8412
rect 7331 8381 7343 8384
rect 7285 8375 7343 8381
rect 9766 8372 9772 8384
rect 9824 8372 9830 8424
rect 10796 8412 10824 8443
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 11514 8480 11520 8492
rect 11475 8452 11520 8480
rect 11514 8440 11520 8452
rect 11572 8440 11578 8492
rect 12710 8480 12716 8492
rect 12671 8452 12716 8480
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 12820 8412 12848 8520
rect 14458 8508 14464 8520
rect 14516 8548 14522 8560
rect 14829 8551 14887 8557
rect 14829 8548 14841 8551
rect 14516 8520 14841 8548
rect 14516 8508 14522 8520
rect 14829 8517 14841 8520
rect 14875 8548 14887 8551
rect 14918 8548 14924 8560
rect 14875 8520 14924 8548
rect 14875 8517 14887 8520
rect 14829 8511 14887 8517
rect 14918 8508 14924 8520
rect 14976 8508 14982 8560
rect 16592 8548 16620 8576
rect 19352 8548 19380 8588
rect 15672 8520 16620 8548
rect 16684 8520 19380 8548
rect 12897 8483 12955 8489
rect 12897 8449 12909 8483
rect 12943 8449 12955 8483
rect 13538 8480 13544 8492
rect 13499 8452 13544 8480
rect 12897 8443 12955 8449
rect 10796 8384 12848 8412
rect 12912 8412 12940 8443
rect 13538 8440 13544 8452
rect 13596 8440 13602 8492
rect 13722 8480 13728 8492
rect 13683 8452 13728 8480
rect 13722 8440 13728 8452
rect 13780 8440 13786 8492
rect 15672 8489 15700 8520
rect 15657 8483 15715 8489
rect 15657 8449 15669 8483
rect 15703 8449 15715 8483
rect 15657 8443 15715 8449
rect 15841 8483 15899 8489
rect 15841 8449 15853 8483
rect 15887 8480 15899 8483
rect 16574 8480 16580 8492
rect 15887 8452 16580 8480
rect 15887 8449 15899 8452
rect 15841 8443 15899 8449
rect 16574 8440 16580 8452
rect 16632 8440 16638 8492
rect 13740 8412 13768 8440
rect 12912 8384 13768 8412
rect 14642 8372 14648 8424
rect 14700 8412 14706 8424
rect 16684 8412 16712 8520
rect 19426 8508 19432 8560
rect 19484 8548 19490 8560
rect 19889 8551 19947 8557
rect 19889 8548 19901 8551
rect 19484 8520 19901 8548
rect 19484 8508 19490 8520
rect 19889 8517 19901 8520
rect 19935 8517 19947 8551
rect 20254 8548 20260 8560
rect 20215 8520 20260 8548
rect 19889 8511 19947 8517
rect 20254 8508 20260 8520
rect 20312 8508 20318 8560
rect 24136 8557 24164 8588
rect 24486 8576 24492 8588
rect 24544 8576 24550 8628
rect 26050 8616 26056 8628
rect 24964 8588 26056 8616
rect 24121 8551 24179 8557
rect 24121 8517 24133 8551
rect 24167 8517 24179 8551
rect 24121 8511 24179 8517
rect 24213 8551 24271 8557
rect 24213 8517 24225 8551
rect 24259 8548 24271 8551
rect 24964 8548 24992 8588
rect 26050 8576 26056 8588
rect 26108 8576 26114 8628
rect 26326 8616 26332 8628
rect 26287 8588 26332 8616
rect 26326 8576 26332 8588
rect 26384 8576 26390 8628
rect 28166 8616 28172 8628
rect 27264 8588 28172 8616
rect 25958 8548 25964 8560
rect 24259 8520 24992 8548
rect 25056 8520 25964 8548
rect 24259 8517 24271 8520
rect 24213 8511 24271 8517
rect 17126 8480 17132 8492
rect 17087 8452 17132 8480
rect 17126 8440 17132 8452
rect 17184 8440 17190 8492
rect 17218 8440 17224 8492
rect 17276 8480 17282 8492
rect 17862 8480 17868 8492
rect 17276 8452 17321 8480
rect 17823 8452 17868 8480
rect 17276 8440 17282 8452
rect 17862 8440 17868 8452
rect 17920 8440 17926 8492
rect 18138 8489 18144 8492
rect 18132 8480 18144 8489
rect 18099 8452 18144 8480
rect 18132 8443 18144 8452
rect 18138 8440 18144 8443
rect 18196 8440 18202 8492
rect 20070 8480 20076 8492
rect 20031 8452 20076 8480
rect 20070 8440 20076 8452
rect 20128 8440 20134 8492
rect 22094 8489 22100 8492
rect 20901 8483 20959 8489
rect 20901 8480 20913 8483
rect 20171 8452 20913 8480
rect 14700 8384 16712 8412
rect 17405 8415 17463 8421
rect 14700 8372 14706 8384
rect 17405 8381 17417 8415
rect 17451 8412 17463 8415
rect 17770 8412 17776 8424
rect 17451 8384 17776 8412
rect 17451 8381 17463 8384
rect 17405 8375 17463 8381
rect 17770 8372 17776 8384
rect 17828 8372 17834 8424
rect 18966 8372 18972 8424
rect 19024 8412 19030 8424
rect 20171 8412 20199 8452
rect 20901 8449 20913 8452
rect 20947 8449 20959 8483
rect 20901 8443 20959 8449
rect 22088 8443 22100 8489
rect 22152 8480 22158 8492
rect 22152 8452 22188 8480
rect 22094 8440 22100 8443
rect 22152 8440 22158 8452
rect 23934 8440 23940 8492
rect 23992 8480 23998 8492
rect 23992 8452 24037 8480
rect 23992 8440 23998 8452
rect 19024 8384 20199 8412
rect 19024 8372 19030 8384
rect 20622 8372 20628 8424
rect 20680 8412 20686 8424
rect 21821 8415 21879 8421
rect 21821 8412 21833 8415
rect 20680 8384 21833 8412
rect 20680 8372 20686 8384
rect 21821 8381 21833 8384
rect 21867 8381 21879 8415
rect 24136 8412 24164 8511
rect 25056 8492 25084 8520
rect 25958 8508 25964 8520
rect 26016 8508 26022 8560
rect 24302 8480 24308 8492
rect 24263 8452 24308 8480
rect 24302 8440 24308 8452
rect 24360 8440 24366 8492
rect 24949 8483 25007 8489
rect 24949 8449 24961 8483
rect 24995 8480 25007 8483
rect 25038 8480 25044 8492
rect 24995 8452 25044 8480
rect 24995 8449 25007 8452
rect 24949 8443 25007 8449
rect 25038 8440 25044 8452
rect 25096 8440 25102 8492
rect 25216 8483 25274 8489
rect 25216 8449 25228 8483
rect 25262 8480 25274 8483
rect 25590 8480 25596 8492
rect 25262 8452 25596 8480
rect 25262 8449 25274 8452
rect 25216 8443 25274 8449
rect 25590 8440 25596 8452
rect 25648 8440 25654 8492
rect 25774 8440 25780 8492
rect 25832 8480 25838 8492
rect 27264 8480 27292 8588
rect 28166 8576 28172 8588
rect 28224 8576 28230 8628
rect 28350 8576 28356 8628
rect 28408 8616 28414 8628
rect 28721 8619 28779 8625
rect 28721 8616 28733 8619
rect 28408 8588 28733 8616
rect 28408 8576 28414 8588
rect 28721 8585 28733 8588
rect 28767 8585 28779 8619
rect 29178 8616 29184 8628
rect 29139 8588 29184 8616
rect 28721 8579 28779 8585
rect 29178 8576 29184 8588
rect 29236 8576 29242 8628
rect 29730 8576 29736 8628
rect 29788 8616 29794 8628
rect 31113 8619 31171 8625
rect 31113 8616 31125 8619
rect 29788 8588 31125 8616
rect 29788 8576 29794 8588
rect 31113 8585 31125 8588
rect 31159 8585 31171 8619
rect 31113 8579 31171 8585
rect 32674 8576 32680 8628
rect 32732 8616 32738 8628
rect 32953 8619 33011 8625
rect 32953 8616 32965 8619
rect 32732 8588 32965 8616
rect 32732 8576 32738 8588
rect 32953 8585 32965 8588
rect 32999 8585 33011 8619
rect 32953 8579 33011 8585
rect 27608 8551 27666 8557
rect 27608 8517 27620 8551
rect 27654 8548 27666 8551
rect 29917 8551 29975 8557
rect 29917 8548 29929 8551
rect 27654 8520 29929 8548
rect 27654 8517 27666 8520
rect 27608 8511 27666 8517
rect 29917 8517 29929 8520
rect 29963 8517 29975 8551
rect 29917 8511 29975 8517
rect 25832 8452 27292 8480
rect 27341 8483 27399 8489
rect 25832 8440 25838 8452
rect 27341 8449 27353 8483
rect 27387 8449 27399 8483
rect 27341 8443 27399 8449
rect 24854 8412 24860 8424
rect 24136 8384 24860 8412
rect 21821 8375 21879 8381
rect 24854 8372 24860 8384
rect 24912 8372 24918 8424
rect 25958 8372 25964 8424
rect 26016 8412 26022 8424
rect 27356 8412 27384 8443
rect 27430 8440 27436 8492
rect 27488 8480 27494 8492
rect 29365 8483 29423 8489
rect 29365 8480 29377 8483
rect 27488 8452 29377 8480
rect 27488 8440 27494 8452
rect 29365 8449 29377 8452
rect 29411 8449 29423 8483
rect 29822 8480 29828 8492
rect 29783 8452 29828 8480
rect 29365 8443 29423 8449
rect 29822 8440 29828 8452
rect 29880 8440 29886 8492
rect 30009 8483 30067 8489
rect 30009 8449 30021 8483
rect 30055 8449 30067 8483
rect 30009 8443 30067 8449
rect 30653 8483 30711 8489
rect 30653 8449 30665 8483
rect 30699 8480 30711 8483
rect 30834 8480 30840 8492
rect 30699 8452 30840 8480
rect 30699 8449 30711 8452
rect 30653 8443 30711 8449
rect 26016 8384 27384 8412
rect 26016 8372 26022 8384
rect 28350 8372 28356 8424
rect 28408 8412 28414 8424
rect 30024 8412 30052 8443
rect 30834 8440 30840 8452
rect 30892 8440 30898 8492
rect 31297 8483 31355 8489
rect 31297 8449 31309 8483
rect 31343 8449 31355 8483
rect 31297 8443 31355 8449
rect 32493 8483 32551 8489
rect 32493 8449 32505 8483
rect 32539 8449 32551 8483
rect 33134 8480 33140 8492
rect 33095 8452 33140 8480
rect 32493 8443 32551 8449
rect 28408 8384 30052 8412
rect 28408 8372 28414 8384
rect 7558 8344 7564 8356
rect 5276 8316 7236 8344
rect 7519 8316 7564 8344
rect 5276 8276 5304 8316
rect 7558 8304 7564 8316
rect 7616 8304 7622 8356
rect 8110 8344 8116 8356
rect 8071 8316 8116 8344
rect 8110 8304 8116 8316
rect 8168 8304 8174 8356
rect 9306 8304 9312 8356
rect 9364 8344 9370 8356
rect 10134 8344 10140 8356
rect 9364 8316 10140 8344
rect 9364 8304 9370 8316
rect 10134 8304 10140 8316
rect 10192 8304 10198 8356
rect 10686 8304 10692 8356
rect 10744 8344 10750 8356
rect 10873 8347 10931 8353
rect 10873 8344 10885 8347
rect 10744 8316 10885 8344
rect 10744 8304 10750 8316
rect 10873 8313 10885 8316
rect 10919 8313 10931 8347
rect 14918 8344 14924 8356
rect 10873 8307 10931 8313
rect 11992 8316 14924 8344
rect 6454 8276 6460 8288
rect 4908 8248 5304 8276
rect 6415 8248 6460 8276
rect 6454 8236 6460 8248
rect 6512 8236 6518 8288
rect 6638 8236 6644 8288
rect 6696 8276 6702 8288
rect 7101 8279 7159 8285
rect 7101 8276 7113 8279
rect 6696 8248 7113 8276
rect 6696 8236 6702 8248
rect 7101 8245 7113 8248
rect 7147 8245 7159 8279
rect 7101 8239 7159 8245
rect 7650 8236 7656 8288
rect 7708 8276 7714 8288
rect 11992 8276 12020 8316
rect 14918 8304 14924 8316
rect 14976 8344 14982 8356
rect 15013 8347 15071 8353
rect 15013 8344 15025 8347
rect 14976 8316 15025 8344
rect 14976 8304 14982 8316
rect 15013 8313 15025 8316
rect 15059 8313 15071 8347
rect 15013 8307 15071 8313
rect 15194 8304 15200 8356
rect 15252 8344 15258 8356
rect 15841 8347 15899 8353
rect 15841 8344 15853 8347
rect 15252 8316 15853 8344
rect 15252 8304 15258 8316
rect 15841 8313 15853 8316
rect 15887 8344 15899 8347
rect 16390 8344 16396 8356
rect 15887 8316 16396 8344
rect 15887 8313 15899 8316
rect 15841 8307 15899 8313
rect 16390 8304 16396 8316
rect 16448 8304 16454 8356
rect 18874 8304 18880 8356
rect 18932 8344 18938 8356
rect 20717 8347 20775 8353
rect 20717 8344 20729 8347
rect 18932 8316 20729 8344
rect 18932 8304 18938 8316
rect 20717 8313 20729 8316
rect 20763 8313 20775 8347
rect 20717 8307 20775 8313
rect 28276 8316 29960 8344
rect 28276 8288 28304 8316
rect 13078 8276 13084 8288
rect 7708 8248 12020 8276
rect 13039 8248 13084 8276
rect 7708 8236 7714 8248
rect 13078 8236 13084 8248
rect 13136 8236 13142 8288
rect 13446 8236 13452 8288
rect 13504 8276 13510 8288
rect 16022 8276 16028 8288
rect 13504 8248 16028 8276
rect 13504 8236 13510 8248
rect 16022 8236 16028 8248
rect 16080 8236 16086 8288
rect 16114 8236 16120 8288
rect 16172 8276 16178 8288
rect 21450 8276 21456 8288
rect 16172 8248 21456 8276
rect 16172 8236 16178 8248
rect 21450 8236 21456 8248
rect 21508 8236 21514 8288
rect 22186 8236 22192 8288
rect 22244 8276 22250 8288
rect 23201 8279 23259 8285
rect 23201 8276 23213 8279
rect 22244 8248 23213 8276
rect 22244 8236 22250 8248
rect 23201 8245 23213 8248
rect 23247 8245 23259 8279
rect 23201 8239 23259 8245
rect 28258 8236 28264 8288
rect 28316 8236 28322 8288
rect 29932 8276 29960 8316
rect 30006 8304 30012 8356
rect 30064 8344 30070 8356
rect 30469 8347 30527 8353
rect 30469 8344 30481 8347
rect 30064 8316 30481 8344
rect 30064 8304 30070 8316
rect 30469 8313 30481 8316
rect 30515 8313 30527 8347
rect 31312 8344 31340 8443
rect 30469 8307 30527 8313
rect 30576 8316 31340 8344
rect 32309 8347 32367 8353
rect 30576 8276 30604 8316
rect 32309 8313 32321 8347
rect 32355 8344 32367 8347
rect 32398 8344 32404 8356
rect 32355 8316 32404 8344
rect 32355 8313 32367 8316
rect 32309 8307 32367 8313
rect 32398 8304 32404 8316
rect 32456 8304 32462 8356
rect 32508 8344 32536 8443
rect 33134 8440 33140 8452
rect 33192 8440 33198 8492
rect 33956 8483 34014 8489
rect 33956 8449 33968 8483
rect 34002 8480 34014 8483
rect 34698 8480 34704 8492
rect 34002 8452 34704 8480
rect 34002 8449 34014 8452
rect 33956 8443 34014 8449
rect 34698 8440 34704 8452
rect 34756 8440 34762 8492
rect 32950 8372 32956 8424
rect 33008 8412 33014 8424
rect 33689 8415 33747 8421
rect 33689 8412 33701 8415
rect 33008 8384 33701 8412
rect 33008 8372 33014 8384
rect 33689 8381 33701 8384
rect 33735 8381 33747 8415
rect 33689 8375 33747 8381
rect 33594 8344 33600 8356
rect 32508 8316 33600 8344
rect 33594 8304 33600 8316
rect 33652 8304 33658 8356
rect 29932 8248 30604 8276
rect 35069 8279 35127 8285
rect 35069 8245 35081 8279
rect 35115 8276 35127 8279
rect 35434 8276 35440 8288
rect 35115 8248 35440 8276
rect 35115 8245 35127 8248
rect 35069 8239 35127 8245
rect 35434 8236 35440 8248
rect 35492 8236 35498 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 2038 8032 2044 8084
rect 2096 8072 2102 8084
rect 2096 8044 5028 8072
rect 2096 8032 2102 8044
rect 2685 8007 2743 8013
rect 2685 8004 2697 8007
rect 1688 7976 2697 8004
rect 1688 7877 1716 7976
rect 2685 7973 2697 7976
rect 2731 8004 2743 8007
rect 4614 8004 4620 8016
rect 2731 7976 4620 8004
rect 2731 7973 2743 7976
rect 2685 7967 2743 7973
rect 4614 7964 4620 7976
rect 4672 7964 4678 8016
rect 5000 8004 5028 8044
rect 9490 8032 9496 8084
rect 9548 8072 9554 8084
rect 9766 8072 9772 8084
rect 9548 8044 9772 8072
rect 9548 8032 9554 8044
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 9858 8032 9864 8084
rect 9916 8072 9922 8084
rect 9953 8075 10011 8081
rect 9953 8072 9965 8075
rect 9916 8044 9965 8072
rect 9916 8032 9922 8044
rect 9953 8041 9965 8044
rect 9999 8041 10011 8075
rect 10410 8072 10416 8084
rect 10371 8044 10416 8072
rect 9953 8035 10011 8041
rect 10410 8032 10416 8044
rect 10468 8032 10474 8084
rect 10594 8032 10600 8084
rect 10652 8072 10658 8084
rect 10965 8075 11023 8081
rect 10965 8072 10977 8075
rect 10652 8044 10977 8072
rect 10652 8032 10658 8044
rect 10965 8041 10977 8044
rect 11011 8041 11023 8075
rect 10965 8035 11023 8041
rect 11425 8075 11483 8081
rect 11425 8041 11437 8075
rect 11471 8072 11483 8075
rect 12434 8072 12440 8084
rect 11471 8044 12440 8072
rect 11471 8041 11483 8044
rect 11425 8035 11483 8041
rect 12434 8032 12440 8044
rect 12492 8032 12498 8084
rect 12989 8075 13047 8081
rect 12989 8041 13001 8075
rect 13035 8072 13047 8075
rect 13538 8072 13544 8084
rect 13035 8044 13544 8072
rect 13035 8041 13047 8044
rect 12989 8035 13047 8041
rect 13538 8032 13544 8044
rect 13596 8032 13602 8084
rect 16114 8072 16120 8084
rect 16075 8044 16120 8072
rect 16114 8032 16120 8044
rect 16172 8032 16178 8084
rect 16574 8072 16580 8084
rect 16535 8044 16580 8072
rect 16574 8032 16580 8044
rect 16632 8032 16638 8084
rect 17494 8072 17500 8084
rect 17455 8044 17500 8072
rect 17494 8032 17500 8044
rect 17552 8032 17558 8084
rect 18049 8075 18107 8081
rect 18049 8041 18061 8075
rect 18095 8072 18107 8075
rect 18138 8072 18144 8084
rect 18095 8044 18144 8072
rect 18095 8041 18107 8044
rect 18049 8035 18107 8041
rect 18138 8032 18144 8044
rect 18196 8032 18202 8084
rect 19797 8075 19855 8081
rect 19797 8041 19809 8075
rect 19843 8072 19855 8075
rect 21266 8072 21272 8084
rect 19843 8044 21272 8072
rect 19843 8041 19855 8044
rect 19797 8035 19855 8041
rect 21266 8032 21272 8044
rect 21324 8032 21330 8084
rect 21913 8075 21971 8081
rect 21913 8041 21925 8075
rect 21959 8072 21971 8075
rect 22094 8072 22100 8084
rect 21959 8044 22100 8072
rect 21959 8041 21971 8044
rect 21913 8035 21971 8041
rect 22094 8032 22100 8044
rect 22152 8032 22158 8084
rect 22278 8072 22284 8084
rect 22239 8044 22284 8072
rect 22278 8032 22284 8044
rect 22336 8032 22342 8084
rect 23201 8075 23259 8081
rect 23201 8041 23213 8075
rect 23247 8072 23259 8075
rect 27430 8072 27436 8084
rect 23247 8044 27436 8072
rect 23247 8041 23259 8044
rect 23201 8035 23259 8041
rect 27430 8032 27436 8044
rect 27488 8032 27494 8084
rect 29086 8032 29092 8084
rect 29144 8072 29150 8084
rect 31481 8075 31539 8081
rect 31481 8072 31493 8075
rect 29144 8044 31493 8072
rect 29144 8032 29150 8044
rect 31481 8041 31493 8044
rect 31527 8041 31539 8075
rect 34698 8072 34704 8084
rect 34659 8044 34704 8072
rect 31481 8035 31539 8041
rect 34698 8032 34704 8044
rect 34756 8032 34762 8084
rect 9306 8004 9312 8016
rect 5000 7976 9312 8004
rect 9306 7964 9312 7976
rect 9364 7964 9370 8016
rect 9398 7964 9404 8016
rect 9456 8004 9462 8016
rect 9456 7976 9501 8004
rect 9456 7964 9462 7976
rect 12250 7964 12256 8016
rect 12308 8004 12314 8016
rect 16482 8004 16488 8016
rect 12308 7976 16488 8004
rect 12308 7964 12314 7976
rect 16482 7964 16488 7976
rect 16540 7964 16546 8016
rect 2317 7939 2375 7945
rect 2317 7905 2329 7939
rect 2363 7936 2375 7939
rect 4706 7936 4712 7948
rect 2363 7908 4712 7936
rect 2363 7905 2375 7908
rect 2317 7899 2375 7905
rect 4706 7896 4712 7908
rect 4764 7896 4770 7948
rect 8941 7939 8999 7945
rect 8941 7905 8953 7939
rect 8987 7936 8999 7939
rect 8987 7908 9076 7936
rect 8987 7905 8999 7908
rect 8941 7899 8999 7905
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7837 1731 7871
rect 1673 7831 1731 7837
rect 1762 7828 1768 7880
rect 1820 7868 1826 7880
rect 1946 7868 1952 7880
rect 1820 7840 1865 7868
rect 1907 7840 1952 7868
rect 1820 7828 1826 7840
rect 1946 7828 1952 7840
rect 2004 7828 2010 7880
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7868 3295 7871
rect 3510 7868 3516 7880
rect 3283 7840 3516 7868
rect 3283 7837 3295 7840
rect 3237 7831 3295 7837
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 5442 7868 5448 7880
rect 4295 7840 5304 7868
rect 5403 7840 5448 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 2314 7760 2320 7812
rect 2372 7800 2378 7812
rect 4433 7803 4491 7809
rect 2372 7772 2728 7800
rect 2372 7760 2378 7772
rect 2700 7732 2728 7772
rect 4433 7769 4445 7803
rect 4479 7800 4491 7803
rect 5074 7800 5080 7812
rect 4479 7772 5080 7800
rect 4479 7769 4491 7772
rect 4433 7763 4491 7769
rect 5074 7760 5080 7772
rect 5132 7760 5138 7812
rect 5276 7800 5304 7840
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 6086 7868 6092 7880
rect 6047 7840 6092 7868
rect 6086 7828 6092 7840
rect 6144 7828 6150 7880
rect 6178 7828 6184 7880
rect 6236 7868 6242 7880
rect 6730 7868 6736 7880
rect 6236 7840 6736 7868
rect 6236 7828 6242 7840
rect 6730 7828 6736 7840
rect 6788 7828 6794 7880
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 7469 7871 7527 7877
rect 7469 7837 7481 7871
rect 7515 7868 7527 7871
rect 7650 7868 7656 7880
rect 7515 7840 7656 7868
rect 7515 7837 7527 7840
rect 7469 7831 7527 7837
rect 5626 7800 5632 7812
rect 5276 7772 5632 7800
rect 5626 7760 5632 7772
rect 5684 7760 5690 7812
rect 7024 7800 7052 7831
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 7745 7871 7803 7877
rect 7745 7837 7757 7871
rect 7791 7868 7803 7871
rect 8110 7868 8116 7880
rect 7791 7840 8116 7868
rect 7791 7837 7803 7840
rect 7745 7831 7803 7837
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 8846 7800 8852 7812
rect 7024 7772 8852 7800
rect 8846 7760 8852 7772
rect 8904 7760 8910 7812
rect 8938 7804 8944 7856
rect 8996 7844 9002 7856
rect 9048 7844 9076 7908
rect 9140 7908 9628 7936
rect 9140 7877 9168 7908
rect 8996 7816 9076 7844
rect 9125 7871 9183 7877
rect 9125 7837 9137 7871
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7868 9275 7871
rect 9306 7868 9312 7880
rect 9263 7840 9312 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 9306 7828 9312 7840
rect 9364 7828 9370 7880
rect 9398 7828 9404 7880
rect 9456 7864 9462 7880
rect 9493 7871 9551 7877
rect 9493 7868 9505 7871
rect 9490 7864 9505 7868
rect 9456 7837 9505 7864
rect 9539 7837 9551 7871
rect 9600 7868 9628 7908
rect 9858 7896 9864 7948
rect 9916 7936 9922 7948
rect 9916 7908 11560 7936
rect 9916 7896 9922 7908
rect 10134 7868 10140 7880
rect 9600 7840 10140 7868
rect 9456 7836 9551 7837
rect 9456 7828 9462 7836
rect 9493 7831 9551 7836
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 10226 7828 10232 7880
rect 10284 7868 10290 7880
rect 10502 7868 10508 7880
rect 10284 7840 10329 7868
rect 10463 7840 10508 7868
rect 10284 7828 10290 7840
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 11149 7871 11207 7877
rect 11149 7837 11161 7871
rect 11195 7837 11207 7871
rect 11149 7831 11207 7837
rect 11241 7871 11299 7877
rect 11241 7837 11253 7871
rect 11287 7868 11299 7871
rect 11330 7868 11336 7880
rect 11287 7840 11336 7868
rect 11287 7837 11299 7840
rect 11241 7831 11299 7837
rect 8996 7804 9002 7816
rect 9766 7760 9772 7812
rect 9824 7800 9830 7812
rect 10686 7800 10692 7812
rect 9824 7772 10692 7800
rect 9824 7760 9830 7772
rect 10686 7760 10692 7772
rect 10744 7760 10750 7812
rect 11164 7800 11192 7831
rect 11330 7828 11336 7840
rect 11388 7828 11394 7880
rect 11532 7877 11560 7908
rect 11606 7896 11612 7948
rect 11664 7936 11670 7948
rect 11977 7939 12035 7945
rect 11977 7936 11989 7939
rect 11664 7908 11989 7936
rect 11664 7896 11670 7908
rect 11977 7905 11989 7908
rect 12023 7905 12035 7939
rect 12434 7936 12440 7948
rect 12347 7908 12440 7936
rect 11977 7899 12035 7905
rect 12434 7896 12440 7908
rect 12492 7936 12498 7948
rect 13449 7939 13507 7945
rect 13449 7936 13461 7939
rect 12492 7908 13461 7936
rect 12492 7896 12498 7908
rect 13449 7905 13461 7908
rect 13495 7936 13507 7939
rect 14458 7936 14464 7948
rect 13495 7908 13676 7936
rect 14419 7908 14464 7936
rect 13495 7905 13507 7908
rect 13449 7899 13507 7905
rect 11517 7871 11575 7877
rect 11517 7837 11529 7871
rect 11563 7837 11575 7871
rect 11517 7831 11575 7837
rect 12161 7871 12219 7877
rect 12161 7837 12173 7871
rect 12207 7837 12219 7871
rect 12161 7831 12219 7837
rect 12176 7800 12204 7831
rect 12250 7828 12256 7880
rect 12308 7868 12314 7880
rect 12526 7868 12532 7880
rect 12308 7840 12353 7868
rect 12487 7840 12532 7868
rect 12308 7828 12314 7840
rect 12526 7828 12532 7840
rect 12584 7828 12590 7880
rect 12986 7828 12992 7880
rect 13044 7868 13050 7880
rect 13173 7871 13231 7877
rect 13173 7868 13185 7871
rect 13044 7840 13185 7868
rect 13044 7828 13050 7840
rect 13173 7837 13185 7840
rect 13219 7837 13231 7871
rect 13173 7831 13231 7837
rect 13265 7871 13323 7877
rect 13265 7837 13277 7871
rect 13311 7868 13323 7871
rect 13354 7868 13360 7880
rect 13311 7840 13360 7868
rect 13311 7837 13323 7840
rect 13265 7831 13323 7837
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 13538 7868 13544 7880
rect 13499 7840 13544 7868
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 13648 7868 13676 7908
rect 14458 7896 14464 7908
rect 14516 7896 14522 7948
rect 14737 7939 14795 7945
rect 14737 7905 14749 7939
rect 14783 7936 14795 7939
rect 16298 7936 16304 7948
rect 14783 7908 16304 7936
rect 14783 7905 14795 7908
rect 14737 7899 14795 7905
rect 13906 7868 13912 7880
rect 13648 7840 13912 7868
rect 13906 7828 13912 7840
rect 13964 7868 13970 7880
rect 14752 7868 14780 7899
rect 16298 7896 16304 7908
rect 16356 7896 16362 7948
rect 16592 7936 16620 8032
rect 20162 7964 20168 8016
rect 20220 8004 20226 8016
rect 20714 8004 20720 8016
rect 20220 7976 20720 8004
rect 20220 7964 20226 7976
rect 20714 7964 20720 7976
rect 20772 7964 20778 8016
rect 21542 7964 21548 8016
rect 21600 8004 21606 8016
rect 25409 8007 25467 8013
rect 21600 7976 23888 8004
rect 21600 7964 21606 7976
rect 16592 7908 17448 7936
rect 13964 7840 14780 7868
rect 13964 7828 13970 7840
rect 15102 7828 15108 7880
rect 15160 7868 15166 7880
rect 16577 7871 16635 7877
rect 16577 7868 16589 7871
rect 15160 7840 16589 7868
rect 15160 7828 15166 7840
rect 16577 7837 16589 7840
rect 16623 7837 16635 7871
rect 16577 7831 16635 7837
rect 16853 7871 16911 7877
rect 16853 7837 16865 7871
rect 16899 7868 16911 7871
rect 16942 7868 16948 7880
rect 16899 7840 16948 7868
rect 16899 7837 16911 7840
rect 16853 7831 16911 7837
rect 16942 7828 16948 7840
rect 17000 7828 17006 7880
rect 17420 7877 17448 7908
rect 17494 7896 17500 7948
rect 17552 7936 17558 7948
rect 17552 7908 21128 7936
rect 17552 7896 17558 7908
rect 17405 7871 17463 7877
rect 17405 7837 17417 7871
rect 17451 7837 17463 7871
rect 18046 7868 18052 7880
rect 18007 7840 18052 7868
rect 17405 7831 17463 7837
rect 18046 7828 18052 7840
rect 18104 7828 18110 7880
rect 18230 7868 18236 7880
rect 18191 7840 18236 7868
rect 18230 7828 18236 7840
rect 18288 7828 18294 7880
rect 18325 7871 18383 7877
rect 18325 7837 18337 7871
rect 18371 7868 18383 7871
rect 19242 7868 19248 7880
rect 18371 7840 19248 7868
rect 18371 7837 18383 7840
rect 18325 7831 18383 7837
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 20438 7868 20444 7880
rect 20399 7840 20444 7868
rect 20438 7828 20444 7840
rect 20496 7828 20502 7880
rect 21100 7877 21128 7908
rect 22186 7896 22192 7948
rect 22244 7936 22250 7948
rect 22373 7939 22431 7945
rect 22373 7936 22385 7939
rect 22244 7908 22385 7936
rect 22244 7896 22250 7908
rect 22373 7905 22385 7908
rect 22419 7905 22431 7939
rect 22373 7899 22431 7905
rect 22756 7908 23060 7936
rect 21085 7871 21143 7877
rect 21085 7837 21097 7871
rect 21131 7837 21143 7871
rect 21085 7831 21143 7837
rect 22097 7871 22155 7877
rect 22097 7837 22109 7871
rect 22143 7868 22155 7871
rect 22756 7868 22784 7908
rect 22922 7868 22928 7880
rect 22143 7840 22784 7868
rect 22883 7840 22928 7868
rect 22143 7837 22155 7840
rect 22097 7831 22155 7837
rect 22922 7828 22928 7840
rect 22980 7828 22986 7880
rect 23032 7877 23060 7908
rect 23474 7896 23480 7948
rect 23532 7936 23538 7948
rect 23658 7936 23664 7948
rect 23532 7908 23664 7936
rect 23532 7896 23538 7908
rect 23658 7896 23664 7908
rect 23716 7896 23722 7948
rect 23860 7877 23888 7976
rect 25409 7973 25421 8007
rect 25455 8004 25467 8007
rect 25455 7976 27476 8004
rect 25455 7973 25467 7976
rect 25409 7967 25467 7973
rect 26602 7936 26608 7948
rect 25240 7908 26608 7936
rect 23017 7871 23075 7877
rect 23017 7837 23029 7871
rect 23063 7868 23075 7871
rect 23845 7871 23903 7877
rect 23063 7840 23796 7868
rect 23063 7837 23075 7840
rect 23017 7831 23075 7837
rect 11164 7772 12204 7800
rect 4338 7732 4344 7744
rect 2700 7704 4344 7732
rect 4338 7692 4344 7704
rect 4396 7692 4402 7744
rect 4617 7735 4675 7741
rect 4617 7701 4629 7735
rect 4663 7732 4675 7735
rect 4798 7732 4804 7744
rect 4663 7704 4804 7732
rect 4663 7701 4675 7704
rect 4617 7695 4675 7701
rect 4798 7692 4804 7704
rect 4856 7692 4862 7744
rect 5261 7735 5319 7741
rect 5261 7701 5273 7735
rect 5307 7732 5319 7735
rect 5810 7732 5816 7744
rect 5307 7704 5816 7732
rect 5307 7701 5319 7704
rect 5261 7695 5319 7701
rect 5810 7692 5816 7704
rect 5868 7692 5874 7744
rect 5905 7735 5963 7741
rect 5905 7701 5917 7735
rect 5951 7732 5963 7735
rect 6454 7732 6460 7744
rect 5951 7704 6460 7732
rect 5951 7701 5963 7704
rect 5905 7695 5963 7701
rect 6454 7692 6460 7704
rect 6512 7692 6518 7744
rect 6825 7735 6883 7741
rect 6825 7701 6837 7735
rect 6871 7732 6883 7735
rect 8478 7732 8484 7744
rect 6871 7704 8484 7732
rect 6871 7701 6883 7704
rect 6825 7695 6883 7701
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 9582 7692 9588 7744
rect 9640 7732 9646 7744
rect 10042 7732 10048 7744
rect 9640 7704 10048 7732
rect 9640 7692 9646 7704
rect 10042 7692 10048 7704
rect 10100 7692 10106 7744
rect 10134 7692 10140 7744
rect 10192 7732 10198 7744
rect 11164 7732 11192 7772
rect 15470 7760 15476 7812
rect 15528 7800 15534 7812
rect 15749 7803 15807 7809
rect 15749 7800 15761 7803
rect 15528 7772 15761 7800
rect 15528 7760 15534 7772
rect 15749 7769 15761 7772
rect 15795 7769 15807 7803
rect 15749 7763 15807 7769
rect 15933 7803 15991 7809
rect 15933 7769 15945 7803
rect 15979 7769 15991 7803
rect 15933 7763 15991 7769
rect 16761 7803 16819 7809
rect 16761 7769 16773 7803
rect 16807 7800 16819 7803
rect 17954 7800 17960 7812
rect 16807 7772 17960 7800
rect 16807 7769 16819 7772
rect 16761 7763 16819 7769
rect 10192 7704 11192 7732
rect 10192 7692 10198 7704
rect 13722 7692 13728 7744
rect 13780 7732 13786 7744
rect 15948 7732 15976 7763
rect 17954 7760 17960 7772
rect 18012 7760 18018 7812
rect 19426 7800 19432 7812
rect 19387 7772 19432 7800
rect 19426 7760 19432 7772
rect 19484 7760 19490 7812
rect 19613 7803 19671 7809
rect 19613 7769 19625 7803
rect 19659 7800 19671 7803
rect 20346 7800 20352 7812
rect 19659 7772 20352 7800
rect 19659 7769 19671 7772
rect 19613 7763 19671 7769
rect 13780 7704 15976 7732
rect 13780 7692 13786 7704
rect 16022 7692 16028 7744
rect 16080 7732 16086 7744
rect 16574 7732 16580 7744
rect 16080 7704 16580 7732
rect 16080 7692 16086 7704
rect 16574 7692 16580 7704
rect 16632 7692 16638 7744
rect 17402 7692 17408 7744
rect 17460 7732 17466 7744
rect 19628 7732 19656 7763
rect 20346 7760 20352 7772
rect 20404 7760 20410 7812
rect 22462 7760 22468 7812
rect 22520 7800 22526 7812
rect 23768 7800 23796 7840
rect 23845 7837 23857 7871
rect 23891 7837 23903 7871
rect 23845 7831 23903 7837
rect 23934 7828 23940 7880
rect 23992 7868 23998 7880
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 23992 7840 24593 7868
rect 23992 7828 23998 7840
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 25130 7868 25136 7880
rect 25091 7840 25136 7868
rect 24581 7831 24639 7837
rect 25130 7828 25136 7840
rect 25188 7828 25194 7880
rect 25240 7877 25268 7908
rect 26602 7896 26608 7908
rect 26660 7896 26666 7948
rect 26973 7939 27031 7945
rect 26973 7905 26985 7939
rect 27019 7905 27031 7939
rect 27338 7936 27344 7948
rect 26973 7899 27031 7905
rect 27264 7908 27344 7936
rect 25225 7871 25283 7877
rect 25225 7837 25237 7871
rect 25271 7837 25283 7871
rect 25225 7831 25283 7837
rect 25406 7828 25412 7880
rect 25464 7868 25470 7880
rect 26053 7871 26111 7877
rect 26053 7868 26065 7871
rect 25464 7840 26065 7868
rect 25464 7828 25470 7840
rect 26053 7837 26065 7840
rect 26099 7837 26111 7871
rect 26053 7831 26111 7837
rect 26694 7828 26700 7880
rect 26752 7868 26758 7880
rect 26789 7871 26847 7877
rect 26789 7868 26801 7871
rect 26752 7840 26801 7868
rect 26752 7828 26758 7840
rect 26789 7837 26801 7840
rect 26835 7837 26847 7871
rect 26789 7831 26847 7837
rect 24486 7800 24492 7812
rect 22520 7772 23704 7800
rect 23768 7772 24492 7800
rect 22520 7760 22526 7772
rect 17460 7704 19656 7732
rect 20257 7735 20315 7741
rect 17460 7692 17466 7704
rect 20257 7701 20269 7735
rect 20303 7732 20315 7735
rect 20530 7732 20536 7744
rect 20303 7704 20536 7732
rect 20303 7701 20315 7704
rect 20257 7695 20315 7701
rect 20530 7692 20536 7704
rect 20588 7692 20594 7744
rect 20714 7692 20720 7744
rect 20772 7732 20778 7744
rect 23676 7741 23704 7772
rect 24486 7760 24492 7772
rect 24544 7760 24550 7812
rect 25038 7760 25044 7812
rect 25096 7800 25102 7812
rect 26988 7800 27016 7899
rect 27264 7877 27292 7908
rect 27338 7896 27344 7908
rect 27396 7896 27402 7948
rect 27448 7936 27476 7976
rect 27614 7964 27620 8016
rect 27672 8004 27678 8016
rect 28626 8004 28632 8016
rect 27672 7976 28632 8004
rect 27672 7964 27678 7976
rect 28626 7964 28632 7976
rect 28684 7964 28690 8016
rect 28994 7964 29000 8016
rect 29052 8004 29058 8016
rect 30193 8007 30251 8013
rect 30193 8004 30205 8007
rect 29052 7976 30205 8004
rect 29052 7964 29058 7976
rect 30193 7973 30205 7976
rect 30239 7973 30251 8007
rect 30193 7967 30251 7973
rect 29270 7936 29276 7948
rect 27448 7908 29276 7936
rect 29270 7896 29276 7908
rect 29328 7896 29334 7948
rect 29454 7896 29460 7948
rect 29512 7936 29518 7948
rect 29512 7908 29776 7936
rect 29512 7896 29518 7908
rect 27065 7871 27123 7877
rect 27065 7837 27077 7871
rect 27111 7868 27123 7871
rect 27249 7871 27307 7877
rect 27111 7840 27200 7868
rect 27111 7837 27123 7840
rect 27065 7831 27123 7837
rect 25096 7772 27016 7800
rect 27172 7800 27200 7840
rect 27249 7837 27261 7871
rect 27295 7837 27307 7871
rect 27522 7868 27528 7880
rect 27483 7840 27528 7868
rect 27249 7831 27307 7837
rect 27522 7828 27528 7840
rect 27580 7828 27586 7880
rect 27614 7828 27620 7880
rect 27672 7868 27678 7880
rect 29748 7877 29776 7908
rect 35176 7908 36124 7936
rect 35176 7880 35204 7908
rect 28997 7871 29055 7877
rect 28997 7868 29009 7871
rect 27672 7840 29009 7868
rect 27672 7828 27678 7840
rect 28997 7837 29009 7840
rect 29043 7837 29055 7871
rect 28997 7831 29055 7837
rect 29549 7871 29607 7877
rect 29549 7837 29561 7871
rect 29595 7837 29607 7871
rect 29549 7831 29607 7837
rect 29733 7871 29791 7877
rect 29733 7837 29745 7871
rect 29779 7837 29791 7871
rect 29733 7831 29791 7837
rect 30377 7871 30435 7877
rect 30377 7837 30389 7871
rect 30423 7868 30435 7871
rect 30466 7868 30472 7880
rect 30423 7840 30472 7868
rect 30423 7837 30435 7840
rect 30377 7831 30435 7837
rect 28074 7800 28080 7812
rect 27172 7772 28080 7800
rect 25096 7760 25102 7772
rect 28074 7760 28080 7772
rect 28132 7760 28138 7812
rect 28169 7803 28227 7809
rect 28169 7769 28181 7803
rect 28215 7800 28227 7803
rect 28258 7800 28264 7812
rect 28215 7772 28264 7800
rect 28215 7769 28227 7772
rect 28169 7763 28227 7769
rect 28258 7760 28264 7772
rect 28316 7760 28322 7812
rect 28353 7803 28411 7809
rect 28353 7769 28365 7803
rect 28399 7800 28411 7803
rect 29564 7800 29592 7831
rect 30466 7828 30472 7840
rect 30524 7828 30530 7880
rect 31018 7868 31024 7880
rect 30979 7840 31024 7868
rect 31018 7828 31024 7840
rect 31076 7828 31082 7880
rect 31662 7868 31668 7880
rect 31623 7840 31668 7868
rect 31662 7828 31668 7840
rect 31720 7828 31726 7880
rect 32309 7871 32367 7877
rect 32309 7837 32321 7871
rect 32355 7868 32367 7871
rect 32950 7868 32956 7880
rect 32355 7840 32956 7868
rect 32355 7837 32367 7840
rect 32309 7831 32367 7837
rect 32950 7828 32956 7840
rect 33008 7828 33014 7880
rect 34885 7871 34943 7877
rect 34885 7868 34897 7871
rect 33060 7840 34897 7868
rect 29822 7800 29828 7812
rect 28399 7772 29828 7800
rect 28399 7769 28411 7772
rect 28353 7763 28411 7769
rect 29822 7760 29828 7772
rect 29880 7800 29886 7812
rect 32576 7803 32634 7809
rect 29880 7772 31754 7800
rect 29880 7760 29886 7772
rect 20901 7735 20959 7741
rect 20901 7732 20913 7735
rect 20772 7704 20913 7732
rect 20772 7692 20778 7704
rect 20901 7701 20913 7704
rect 20947 7701 20959 7735
rect 20901 7695 20959 7701
rect 23661 7735 23719 7741
rect 23661 7701 23673 7735
rect 23707 7701 23719 7735
rect 23661 7695 23719 7701
rect 23750 7692 23756 7744
rect 23808 7732 23814 7744
rect 24397 7735 24455 7741
rect 24397 7732 24409 7735
rect 23808 7704 24409 7732
rect 23808 7692 23814 7704
rect 24397 7701 24409 7704
rect 24443 7701 24455 7735
rect 24397 7695 24455 7701
rect 25498 7692 25504 7744
rect 25556 7732 25562 7744
rect 25869 7735 25927 7741
rect 25869 7732 25881 7735
rect 25556 7704 25881 7732
rect 25556 7692 25562 7704
rect 25869 7701 25881 7704
rect 25915 7701 25927 7735
rect 25869 7695 25927 7701
rect 26694 7692 26700 7744
rect 26752 7732 26758 7744
rect 28813 7735 28871 7741
rect 28813 7732 28825 7735
rect 26752 7704 28825 7732
rect 26752 7692 26758 7704
rect 28813 7701 28825 7704
rect 28859 7701 28871 7735
rect 28813 7695 28871 7701
rect 28902 7692 28908 7744
rect 28960 7732 28966 7744
rect 29641 7735 29699 7741
rect 29641 7732 29653 7735
rect 28960 7704 29653 7732
rect 28960 7692 28966 7704
rect 29641 7701 29653 7704
rect 29687 7701 29699 7735
rect 29641 7695 29699 7701
rect 30374 7692 30380 7744
rect 30432 7732 30438 7744
rect 30837 7735 30895 7741
rect 30837 7732 30849 7735
rect 30432 7704 30849 7732
rect 30432 7692 30438 7704
rect 30837 7701 30849 7704
rect 30883 7701 30895 7735
rect 31726 7732 31754 7772
rect 32576 7769 32588 7803
rect 32622 7800 32634 7803
rect 32858 7800 32864 7812
rect 32622 7772 32864 7800
rect 32622 7769 32634 7772
rect 32576 7763 32634 7769
rect 32858 7760 32864 7772
rect 32916 7760 32922 7812
rect 33060 7744 33088 7840
rect 34885 7837 34897 7840
rect 34931 7837 34943 7871
rect 35158 7868 35164 7880
rect 35119 7840 35164 7868
rect 34885 7831 34943 7837
rect 34900 7800 34928 7831
rect 35158 7828 35164 7840
rect 35216 7828 35222 7880
rect 36096 7877 36124 7908
rect 35805 7871 35863 7877
rect 35805 7837 35817 7871
rect 35851 7837 35863 7871
rect 35805 7831 35863 7837
rect 36081 7871 36139 7877
rect 36081 7837 36093 7871
rect 36127 7837 36139 7871
rect 36081 7831 36139 7837
rect 35820 7800 35848 7831
rect 34900 7772 35848 7800
rect 33042 7732 33048 7744
rect 31726 7704 33048 7732
rect 30837 7695 30895 7701
rect 33042 7692 33048 7704
rect 33100 7692 33106 7744
rect 33689 7735 33747 7741
rect 33689 7701 33701 7735
rect 33735 7732 33747 7735
rect 34698 7732 34704 7744
rect 33735 7704 34704 7732
rect 33735 7701 33747 7704
rect 33689 7695 33747 7701
rect 34698 7692 34704 7704
rect 34756 7692 34762 7744
rect 35069 7735 35127 7741
rect 35069 7701 35081 7735
rect 35115 7732 35127 7735
rect 35434 7732 35440 7744
rect 35115 7704 35440 7732
rect 35115 7701 35127 7704
rect 35069 7695 35127 7701
rect 35434 7692 35440 7704
rect 35492 7692 35498 7744
rect 35618 7732 35624 7744
rect 35579 7704 35624 7732
rect 35618 7692 35624 7704
rect 35676 7692 35682 7744
rect 35989 7735 36047 7741
rect 35989 7701 36001 7735
rect 36035 7732 36047 7735
rect 36078 7732 36084 7744
rect 36035 7704 36084 7732
rect 36035 7701 36047 7704
rect 35989 7695 36047 7701
rect 36078 7692 36084 7704
rect 36136 7692 36142 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 1397 7531 1455 7537
rect 1397 7497 1409 7531
rect 1443 7528 1455 7531
rect 1762 7528 1768 7540
rect 1443 7500 1768 7528
rect 1443 7497 1455 7500
rect 1397 7491 1455 7497
rect 1762 7488 1768 7500
rect 1820 7488 1826 7540
rect 2314 7528 2320 7540
rect 2275 7500 2320 7528
rect 2314 7488 2320 7500
rect 2372 7488 2378 7540
rect 2958 7528 2964 7540
rect 2516 7500 2774 7528
rect 2919 7500 2964 7528
rect 934 7352 940 7404
rect 992 7392 998 7404
rect 2516 7401 2544 7500
rect 2746 7460 2774 7500
rect 2958 7488 2964 7500
rect 3016 7488 3022 7540
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 5445 7531 5503 7537
rect 5445 7528 5457 7531
rect 4120 7500 5457 7528
rect 4120 7488 4126 7500
rect 5445 7497 5457 7500
rect 5491 7497 5503 7531
rect 5445 7491 5503 7497
rect 5810 7488 5816 7540
rect 5868 7528 5874 7540
rect 5868 7500 8708 7528
rect 5868 7488 5874 7500
rect 2746 7432 4108 7460
rect 3878 7401 3884 7404
rect 1581 7395 1639 7401
rect 1581 7392 1593 7395
rect 992 7364 1593 7392
rect 992 7352 998 7364
rect 1581 7361 1593 7364
rect 1627 7361 1639 7395
rect 1581 7355 1639 7361
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7361 2559 7395
rect 2501 7355 2559 7361
rect 3145 7395 3203 7401
rect 3145 7361 3157 7395
rect 3191 7361 3203 7395
rect 3145 7355 3203 7361
rect 3872 7355 3884 7401
rect 3936 7392 3942 7404
rect 4080 7392 4108 7432
rect 4338 7420 4344 7472
rect 4396 7460 4402 7472
rect 6178 7460 6184 7472
rect 4396 7432 6184 7460
rect 4396 7420 4402 7432
rect 6178 7420 6184 7432
rect 6236 7420 6242 7472
rect 8478 7469 8484 7472
rect 8472 7460 8484 7469
rect 6380 7432 8248 7460
rect 8439 7432 8484 7460
rect 6380 7404 6408 7432
rect 3936 7364 3972 7392
rect 4080 7364 4660 7392
rect 3160 7188 3188 7355
rect 3878 7352 3884 7355
rect 3936 7352 3942 7364
rect 3602 7324 3608 7336
rect 3563 7296 3608 7324
rect 3602 7284 3608 7296
rect 3660 7284 3666 7336
rect 4632 7324 4660 7364
rect 4798 7352 4804 7404
rect 4856 7392 4862 7404
rect 5629 7395 5687 7401
rect 5629 7392 5641 7395
rect 4856 7364 5641 7392
rect 4856 7352 4862 7364
rect 5629 7361 5641 7364
rect 5675 7361 5687 7395
rect 6362 7392 6368 7404
rect 6323 7364 6368 7392
rect 5629 7355 5687 7361
rect 6362 7352 6368 7364
rect 6420 7352 6426 7404
rect 6454 7352 6460 7404
rect 6512 7392 6518 7404
rect 8220 7401 8248 7432
rect 8472 7423 8484 7432
rect 8478 7420 8484 7423
rect 8536 7420 8542 7472
rect 8680 7460 8708 7500
rect 9490 7488 9496 7540
rect 9548 7528 9554 7540
rect 10042 7528 10048 7540
rect 9548 7500 10048 7528
rect 9548 7488 9554 7500
rect 10042 7488 10048 7500
rect 10100 7528 10106 7540
rect 10410 7528 10416 7540
rect 10100 7500 10416 7528
rect 10100 7488 10106 7500
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 15102 7528 15108 7540
rect 12268 7500 15108 7528
rect 12130 7463 12188 7469
rect 12130 7460 12142 7463
rect 8680 7432 12142 7460
rect 12130 7429 12142 7432
rect 12176 7429 12188 7463
rect 12130 7423 12188 7429
rect 6621 7395 6679 7401
rect 6621 7392 6633 7395
rect 6512 7364 6633 7392
rect 6512 7352 6518 7364
rect 6621 7361 6633 7364
rect 6667 7361 6679 7395
rect 6621 7355 6679 7361
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7361 8263 7395
rect 9490 7392 9496 7404
rect 8205 7355 8263 7361
rect 8312 7364 9496 7392
rect 4632 7296 5580 7324
rect 4614 7216 4620 7268
rect 4672 7256 4678 7268
rect 4985 7259 5043 7265
rect 4985 7256 4997 7259
rect 4672 7228 4997 7256
rect 4672 7216 4678 7228
rect 4985 7225 4997 7228
rect 5031 7256 5043 7259
rect 5258 7256 5264 7268
rect 5031 7228 5264 7256
rect 5031 7225 5043 7228
rect 4985 7219 5043 7225
rect 5258 7216 5264 7228
rect 5316 7216 5322 7268
rect 5442 7188 5448 7200
rect 3160 7160 5448 7188
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 5552 7188 5580 7296
rect 8110 7284 8116 7336
rect 8168 7324 8174 7336
rect 8312 7324 8340 7364
rect 9490 7352 9496 7364
rect 9548 7352 9554 7404
rect 10134 7352 10140 7404
rect 10192 7392 10198 7404
rect 10321 7395 10379 7401
rect 10321 7392 10333 7395
rect 10192 7364 10333 7392
rect 10192 7352 10198 7364
rect 10321 7361 10333 7364
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 10962 7352 10968 7404
rect 11020 7392 11026 7404
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 11020 7364 11897 7392
rect 11020 7352 11026 7364
rect 11885 7361 11897 7364
rect 11931 7361 11943 7395
rect 12268 7392 12296 7500
rect 15102 7488 15108 7500
rect 15160 7488 15166 7540
rect 15470 7528 15476 7540
rect 15431 7500 15476 7528
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 18230 7488 18236 7540
rect 18288 7528 18294 7540
rect 18598 7528 18604 7540
rect 18288 7500 18604 7528
rect 18288 7488 18294 7500
rect 18598 7488 18604 7500
rect 18656 7528 18662 7540
rect 18656 7500 19334 7528
rect 18656 7488 18662 7500
rect 12342 7420 12348 7472
rect 12400 7460 12406 7472
rect 18325 7463 18383 7469
rect 18325 7460 18337 7463
rect 12400 7432 18337 7460
rect 12400 7420 12406 7432
rect 18325 7429 18337 7432
rect 18371 7429 18383 7463
rect 18325 7423 18383 7429
rect 11885 7355 11943 7361
rect 11992 7364 12296 7392
rect 8168 7296 8340 7324
rect 8168 7284 8174 7296
rect 9766 7284 9772 7336
rect 9824 7324 9830 7336
rect 10045 7327 10103 7333
rect 10045 7324 10057 7327
rect 9824 7296 10057 7324
rect 9824 7284 9830 7296
rect 10045 7293 10057 7296
rect 10091 7293 10103 7327
rect 11992 7324 12020 7364
rect 12434 7352 12440 7404
rect 12492 7392 12498 7404
rect 12492 7364 12940 7392
rect 12492 7352 12498 7364
rect 10045 7287 10103 7293
rect 10152 7296 12020 7324
rect 12912 7324 12940 7364
rect 13078 7352 13084 7404
rect 13136 7392 13142 7404
rect 15657 7395 15715 7401
rect 13136 7364 14504 7392
rect 13136 7352 13142 7364
rect 13446 7324 13452 7336
rect 12912 7296 13452 7324
rect 9398 7216 9404 7268
rect 9456 7256 9462 7268
rect 10152 7256 10180 7296
rect 13446 7284 13452 7296
rect 13504 7284 13510 7336
rect 14476 7333 14504 7364
rect 15657 7361 15669 7395
rect 15703 7361 15715 7395
rect 15657 7355 15715 7361
rect 14185 7327 14243 7333
rect 14185 7293 14197 7327
rect 14231 7293 14243 7327
rect 14185 7287 14243 7293
rect 14461 7327 14519 7333
rect 14461 7293 14473 7327
rect 14507 7324 14519 7327
rect 15672 7324 15700 7355
rect 15746 7352 15752 7404
rect 15804 7392 15810 7404
rect 16022 7392 16028 7404
rect 15804 7364 15849 7392
rect 15983 7364 16028 7392
rect 15804 7352 15810 7364
rect 16022 7352 16028 7364
rect 16080 7352 16086 7404
rect 16574 7352 16580 7404
rect 16632 7392 16638 7404
rect 16945 7395 17003 7401
rect 16945 7392 16957 7395
rect 16632 7364 16957 7392
rect 16632 7352 16638 7364
rect 16945 7361 16957 7364
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 17126 7352 17132 7404
rect 17184 7392 17190 7404
rect 18233 7395 18291 7401
rect 18233 7392 18245 7395
rect 17184 7364 18245 7392
rect 17184 7352 17190 7364
rect 18233 7361 18245 7364
rect 18279 7361 18291 7395
rect 19306 7392 19334 7500
rect 20346 7488 20352 7540
rect 20404 7528 20410 7540
rect 22370 7528 22376 7540
rect 20404 7500 21128 7528
rect 22331 7500 22376 7528
rect 20404 7488 20410 7500
rect 21100 7469 21128 7500
rect 22370 7488 22376 7500
rect 22428 7488 22434 7540
rect 22738 7488 22744 7540
rect 22796 7528 22802 7540
rect 25777 7531 25835 7537
rect 25777 7528 25789 7531
rect 22796 7500 25789 7528
rect 22796 7488 22802 7500
rect 25777 7497 25789 7500
rect 25823 7497 25835 7531
rect 25777 7491 25835 7497
rect 27338 7488 27344 7540
rect 27396 7528 27402 7540
rect 28353 7531 28411 7537
rect 28353 7528 28365 7531
rect 27396 7500 28365 7528
rect 27396 7488 27402 7500
rect 28353 7497 28365 7500
rect 28399 7497 28411 7531
rect 29270 7528 29276 7540
rect 28353 7491 28411 7497
rect 28966 7500 29276 7528
rect 21085 7463 21143 7469
rect 21085 7429 21097 7463
rect 21131 7460 21143 7463
rect 22189 7463 22247 7469
rect 22189 7460 22201 7463
rect 21131 7432 22201 7460
rect 21131 7429 21143 7432
rect 21085 7423 21143 7429
rect 22189 7429 22201 7432
rect 22235 7429 22247 7463
rect 22189 7423 22247 7429
rect 24026 7420 24032 7472
rect 24084 7460 24090 7472
rect 24210 7460 24216 7472
rect 24084 7432 24216 7460
rect 24084 7420 24090 7432
rect 24210 7420 24216 7432
rect 24268 7460 24274 7472
rect 24268 7432 24440 7460
rect 24268 7420 24274 7432
rect 19521 7395 19579 7401
rect 19521 7392 19533 7395
rect 19306 7364 19533 7392
rect 18233 7355 18291 7361
rect 19521 7361 19533 7364
rect 19567 7361 19579 7395
rect 20898 7392 20904 7404
rect 20859 7364 20904 7392
rect 19521 7355 19579 7361
rect 20898 7352 20904 7364
rect 20956 7352 20962 7404
rect 22005 7395 22063 7401
rect 22005 7361 22017 7395
rect 22051 7392 22063 7395
rect 22094 7392 22100 7404
rect 22051 7364 22100 7392
rect 22051 7361 22063 7364
rect 22005 7355 22063 7361
rect 22094 7352 22100 7364
rect 22152 7352 22158 7404
rect 23014 7392 23020 7404
rect 22975 7364 23020 7392
rect 23014 7352 23020 7364
rect 23072 7352 23078 7404
rect 23658 7392 23664 7404
rect 23619 7364 23664 7392
rect 23658 7352 23664 7364
rect 23716 7352 23722 7404
rect 24302 7392 24308 7404
rect 24263 7364 24308 7392
rect 24302 7352 24308 7364
rect 24360 7352 24366 7404
rect 24412 7401 24440 7432
rect 24486 7420 24492 7472
rect 24544 7460 24550 7472
rect 27240 7463 27298 7469
rect 24544 7432 27200 7460
rect 24544 7420 24550 7432
rect 24397 7395 24455 7401
rect 24397 7361 24409 7395
rect 24443 7361 24455 7395
rect 24397 7355 24455 7361
rect 24673 7395 24731 7401
rect 24673 7361 24685 7395
rect 24719 7392 24731 7395
rect 24762 7392 24768 7404
rect 24719 7364 24768 7392
rect 24719 7361 24731 7364
rect 24673 7355 24731 7361
rect 24762 7352 24768 7364
rect 24820 7352 24826 7404
rect 25314 7392 25320 7404
rect 25275 7364 25320 7392
rect 25314 7352 25320 7364
rect 25372 7352 25378 7404
rect 25958 7392 25964 7404
rect 25919 7364 25964 7392
rect 25958 7352 25964 7364
rect 26016 7352 26022 7404
rect 26973 7395 27031 7401
rect 26973 7361 26985 7395
rect 27019 7392 27031 7395
rect 27062 7392 27068 7404
rect 27019 7364 27068 7392
rect 27019 7361 27031 7364
rect 26973 7355 27031 7361
rect 27062 7352 27068 7364
rect 27120 7352 27126 7404
rect 27172 7392 27200 7432
rect 27240 7429 27252 7463
rect 27286 7460 27298 7463
rect 28074 7460 28080 7472
rect 27286 7432 28080 7460
rect 27286 7429 27298 7432
rect 27240 7423 27298 7429
rect 28074 7420 28080 7432
rect 28132 7420 28138 7472
rect 28966 7392 28994 7500
rect 29270 7488 29276 7500
rect 29328 7528 29334 7540
rect 29411 7531 29469 7537
rect 29411 7528 29423 7531
rect 29328 7500 29423 7528
rect 29328 7488 29334 7500
rect 29411 7497 29423 7500
rect 29457 7528 29469 7531
rect 30669 7531 30727 7537
rect 30669 7528 30681 7531
rect 29457 7500 30681 7528
rect 29457 7497 29469 7500
rect 29411 7491 29469 7497
rect 30669 7497 30681 7500
rect 30715 7497 30727 7531
rect 30834 7528 30840 7540
rect 30795 7500 30840 7528
rect 30669 7491 30727 7497
rect 30834 7488 30840 7500
rect 30892 7488 30898 7540
rect 32858 7528 32864 7540
rect 32819 7500 32864 7528
rect 32858 7488 32864 7500
rect 32916 7488 32922 7540
rect 33229 7531 33287 7537
rect 33229 7497 33241 7531
rect 33275 7528 33287 7531
rect 34698 7528 34704 7540
rect 33275 7500 34704 7528
rect 33275 7497 33287 7500
rect 33229 7491 33287 7497
rect 34698 7488 34704 7500
rect 34756 7488 34762 7540
rect 35161 7531 35219 7537
rect 35161 7497 35173 7531
rect 35207 7528 35219 7531
rect 36078 7528 36084 7540
rect 35207 7500 36084 7528
rect 35207 7497 35219 7500
rect 35161 7491 35219 7497
rect 36078 7488 36084 7500
rect 36136 7488 36142 7540
rect 30469 7463 30527 7469
rect 30469 7429 30481 7463
rect 30515 7429 30527 7463
rect 30469 7423 30527 7429
rect 29178 7392 29184 7404
rect 27172 7364 28994 7392
rect 29139 7364 29184 7392
rect 29178 7352 29184 7364
rect 29236 7392 29242 7404
rect 30484 7392 30512 7423
rect 32766 7420 32772 7472
rect 32824 7460 32830 7472
rect 34048 7463 34106 7469
rect 32824 7432 33364 7460
rect 32824 7420 32830 7432
rect 31202 7392 31208 7404
rect 29236 7364 29316 7392
rect 30484 7364 31208 7392
rect 29236 7352 29242 7364
rect 16114 7324 16120 7336
rect 14507 7296 16120 7324
rect 14507 7293 14519 7296
rect 14461 7287 14519 7293
rect 14200 7256 14228 7287
rect 16114 7284 16120 7296
rect 16172 7284 16178 7336
rect 17221 7327 17279 7333
rect 17221 7293 17233 7327
rect 17267 7324 17279 7327
rect 17402 7324 17408 7336
rect 17267 7296 17408 7324
rect 17267 7293 17279 7296
rect 17221 7287 17279 7293
rect 17402 7284 17408 7296
rect 17460 7284 17466 7336
rect 19245 7327 19303 7333
rect 19245 7293 19257 7327
rect 19291 7324 19303 7327
rect 20438 7324 20444 7336
rect 19291 7296 20444 7324
rect 19291 7293 19303 7296
rect 19245 7287 19303 7293
rect 9456 7228 10180 7256
rect 13188 7228 14228 7256
rect 9456 7216 9462 7228
rect 6546 7188 6552 7200
rect 5552 7160 6552 7188
rect 6546 7148 6552 7160
rect 6604 7148 6610 7200
rect 6638 7148 6644 7200
rect 6696 7188 6702 7200
rect 7745 7191 7803 7197
rect 7745 7188 7757 7191
rect 6696 7160 7757 7188
rect 6696 7148 6702 7160
rect 7745 7157 7757 7160
rect 7791 7157 7803 7191
rect 7745 7151 7803 7157
rect 9214 7148 9220 7200
rect 9272 7188 9278 7200
rect 9585 7191 9643 7197
rect 9585 7188 9597 7191
rect 9272 7160 9597 7188
rect 9272 7148 9278 7160
rect 9585 7157 9597 7160
rect 9631 7157 9643 7191
rect 9585 7151 9643 7157
rect 10686 7148 10692 7200
rect 10744 7188 10750 7200
rect 13188 7188 13216 7228
rect 14918 7216 14924 7268
rect 14976 7256 14982 7268
rect 15933 7259 15991 7265
rect 15933 7256 15945 7259
rect 14976 7228 15945 7256
rect 14976 7216 14982 7228
rect 15933 7225 15945 7228
rect 15979 7256 15991 7259
rect 19260 7256 19288 7287
rect 20438 7284 20444 7296
rect 20496 7284 20502 7336
rect 21269 7327 21327 7333
rect 21269 7293 21281 7327
rect 21315 7324 21327 7327
rect 23934 7324 23940 7336
rect 21315 7296 23940 7324
rect 21315 7293 21327 7296
rect 21269 7287 21327 7293
rect 23934 7284 23940 7296
rect 23992 7284 23998 7336
rect 28074 7284 28080 7336
rect 28132 7324 28138 7336
rect 28902 7324 28908 7336
rect 28132 7296 28908 7324
rect 28132 7284 28138 7296
rect 28902 7284 28908 7296
rect 28960 7284 28966 7336
rect 15979 7228 19288 7256
rect 15979 7225 15991 7228
rect 15933 7219 15991 7225
rect 20254 7216 20260 7268
rect 20312 7256 20318 7268
rect 23477 7259 23535 7265
rect 23477 7256 23489 7259
rect 20312 7228 23489 7256
rect 20312 7216 20318 7228
rect 23477 7225 23489 7228
rect 23523 7225 23535 7259
rect 23477 7219 23535 7225
rect 24394 7216 24400 7268
rect 24452 7256 24458 7268
rect 25133 7259 25191 7265
rect 25133 7256 25145 7259
rect 24452 7228 25145 7256
rect 24452 7216 24458 7228
rect 25133 7225 25145 7228
rect 25179 7225 25191 7259
rect 29288 7256 29316 7364
rect 31202 7352 31208 7364
rect 31260 7352 31266 7404
rect 31481 7395 31539 7401
rect 31481 7361 31493 7395
rect 31527 7361 31539 7395
rect 31481 7355 31539 7361
rect 32401 7395 32459 7401
rect 32401 7361 32413 7395
rect 32447 7392 32459 7395
rect 32490 7392 32496 7404
rect 32447 7364 32496 7392
rect 32447 7361 32459 7364
rect 32401 7355 32459 7361
rect 30190 7284 30196 7336
rect 30248 7324 30254 7336
rect 31496 7324 31524 7355
rect 32490 7352 32496 7364
rect 32548 7352 32554 7404
rect 33042 7392 33048 7404
rect 33003 7364 33048 7392
rect 33042 7352 33048 7364
rect 33100 7352 33106 7404
rect 33336 7401 33364 7432
rect 34048 7429 34060 7463
rect 34094 7460 34106 7463
rect 35618 7460 35624 7472
rect 34094 7432 35624 7460
rect 34094 7429 34106 7432
rect 34048 7423 34106 7429
rect 35618 7420 35624 7432
rect 35676 7420 35682 7472
rect 33321 7395 33379 7401
rect 33321 7361 33333 7395
rect 33367 7392 33379 7395
rect 35158 7392 35164 7404
rect 33367 7364 35164 7392
rect 33367 7361 33379 7364
rect 33321 7355 33379 7361
rect 35158 7352 35164 7364
rect 35216 7352 35222 7404
rect 35710 7352 35716 7404
rect 35768 7392 35774 7404
rect 35805 7395 35863 7401
rect 35805 7392 35817 7395
rect 35768 7364 35817 7392
rect 35768 7352 35774 7364
rect 35805 7361 35817 7364
rect 35851 7361 35863 7395
rect 36446 7392 36452 7404
rect 36407 7364 36452 7392
rect 35805 7355 35863 7361
rect 36446 7352 36452 7364
rect 36504 7352 36510 7404
rect 30248 7296 31524 7324
rect 30248 7284 30254 7296
rect 32950 7284 32956 7336
rect 33008 7324 33014 7336
rect 33781 7327 33839 7333
rect 33781 7324 33793 7327
rect 33008 7296 33793 7324
rect 33008 7284 33014 7296
rect 33781 7293 33793 7296
rect 33827 7293 33839 7327
rect 33781 7287 33839 7293
rect 31938 7256 31944 7268
rect 29288 7228 31944 7256
rect 25133 7219 25191 7225
rect 31938 7216 31944 7228
rect 31996 7216 32002 7268
rect 34790 7216 34796 7268
rect 34848 7256 34854 7268
rect 36265 7259 36323 7265
rect 36265 7256 36277 7259
rect 34848 7228 36277 7256
rect 34848 7216 34854 7228
rect 36265 7225 36277 7228
rect 36311 7225 36323 7259
rect 36265 7219 36323 7225
rect 10744 7160 13216 7188
rect 10744 7148 10750 7160
rect 13262 7148 13268 7200
rect 13320 7188 13326 7200
rect 13320 7160 13365 7188
rect 13320 7148 13326 7160
rect 13446 7148 13452 7200
rect 13504 7188 13510 7200
rect 15654 7188 15660 7200
rect 13504 7160 15660 7188
rect 13504 7148 13510 7160
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 22833 7191 22891 7197
rect 22833 7157 22845 7191
rect 22879 7188 22891 7191
rect 23198 7188 23204 7200
rect 22879 7160 23204 7188
rect 22879 7157 22891 7160
rect 22833 7151 22891 7157
rect 23198 7148 23204 7160
rect 23256 7148 23262 7200
rect 24118 7188 24124 7200
rect 24079 7160 24124 7188
rect 24118 7148 24124 7160
rect 24176 7148 24182 7200
rect 24581 7191 24639 7197
rect 24581 7157 24593 7191
rect 24627 7188 24639 7191
rect 24946 7188 24952 7200
rect 24627 7160 24952 7188
rect 24627 7157 24639 7160
rect 24581 7151 24639 7157
rect 24946 7148 24952 7160
rect 25004 7148 25010 7200
rect 29178 7148 29184 7200
rect 29236 7188 29242 7200
rect 30653 7191 30711 7197
rect 30653 7188 30665 7191
rect 29236 7160 30665 7188
rect 29236 7148 29242 7160
rect 30653 7157 30665 7160
rect 30699 7157 30711 7191
rect 30653 7151 30711 7157
rect 31297 7191 31355 7197
rect 31297 7157 31309 7191
rect 31343 7188 31355 7191
rect 32122 7188 32128 7200
rect 31343 7160 32128 7188
rect 31343 7157 31355 7160
rect 31297 7151 31355 7157
rect 32122 7148 32128 7160
rect 32180 7148 32186 7200
rect 32217 7191 32275 7197
rect 32217 7157 32229 7191
rect 32263 7188 32275 7191
rect 33410 7188 33416 7200
rect 32263 7160 33416 7188
rect 32263 7157 32275 7160
rect 32217 7151 32275 7157
rect 33410 7148 33416 7160
rect 33468 7148 33474 7200
rect 35434 7148 35440 7200
rect 35492 7188 35498 7200
rect 35621 7191 35679 7197
rect 35621 7188 35633 7191
rect 35492 7160 35633 7188
rect 35492 7148 35498 7160
rect 35621 7157 35633 7160
rect 35667 7157 35679 7191
rect 35621 7151 35679 7157
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1765 6987 1823 6993
rect 1765 6953 1777 6987
rect 1811 6984 1823 6987
rect 2130 6984 2136 6996
rect 1811 6956 2136 6984
rect 1811 6953 1823 6956
rect 1765 6947 1823 6953
rect 2130 6944 2136 6956
rect 2188 6944 2194 6996
rect 2958 6944 2964 6996
rect 3016 6984 3022 6996
rect 3053 6987 3111 6993
rect 3053 6984 3065 6987
rect 3016 6956 3065 6984
rect 3016 6944 3022 6956
rect 3053 6953 3065 6956
rect 3099 6953 3111 6987
rect 3053 6947 3111 6953
rect 3252 6956 9168 6984
rect 3050 6848 3056 6860
rect 1964 6820 3056 6848
rect 1964 6789 1992 6820
rect 3050 6808 3056 6820
rect 3108 6808 3114 6860
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6749 2007 6783
rect 1949 6743 2007 6749
rect 2593 6783 2651 6789
rect 2593 6749 2605 6783
rect 2639 6780 2651 6783
rect 2958 6780 2964 6792
rect 2639 6752 2964 6780
rect 2639 6749 2651 6752
rect 2593 6743 2651 6749
rect 2958 6740 2964 6752
rect 3016 6740 3022 6792
rect 3252 6789 3280 6956
rect 5169 6919 5227 6925
rect 5169 6885 5181 6919
rect 5215 6916 5227 6919
rect 7650 6916 7656 6928
rect 5215 6888 5948 6916
rect 5215 6885 5227 6888
rect 5169 6879 5227 6885
rect 3602 6808 3608 6860
rect 3660 6848 3666 6860
rect 3789 6851 3847 6857
rect 3789 6848 3801 6851
rect 3660 6820 3801 6848
rect 3660 6808 3666 6820
rect 3789 6817 3801 6820
rect 3835 6817 3847 6851
rect 5626 6848 5632 6860
rect 5587 6820 5632 6848
rect 3789 6811 3847 6817
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 5920 6848 5948 6888
rect 6932 6888 7656 6916
rect 5994 6848 6000 6860
rect 5920 6820 6000 6848
rect 4062 6789 4068 6792
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6749 3295 6783
rect 4056 6780 4068 6789
rect 4023 6752 4068 6780
rect 3237 6743 3295 6749
rect 4056 6743 4068 6752
rect 4062 6740 4068 6743
rect 4120 6740 4126 6792
rect 5920 6789 5948 6820
rect 5994 6808 6000 6820
rect 6052 6808 6058 6860
rect 6932 6857 6960 6888
rect 7650 6876 7656 6888
rect 7708 6876 7714 6928
rect 9140 6916 9168 6956
rect 9214 6944 9220 6996
rect 9272 6984 9278 6996
rect 9272 6956 9317 6984
rect 9272 6944 9278 6956
rect 9398 6944 9404 6996
rect 9456 6984 9462 6996
rect 11701 6987 11759 6993
rect 9456 6956 9501 6984
rect 10336 6956 11652 6984
rect 9456 6944 9462 6956
rect 10336 6916 10364 6956
rect 9140 6888 10364 6916
rect 11624 6916 11652 6956
rect 11701 6953 11713 6987
rect 11747 6984 11759 6987
rect 12250 6984 12256 6996
rect 11747 6956 12256 6984
rect 11747 6953 11759 6956
rect 11701 6947 11759 6953
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 12989 6987 13047 6993
rect 12989 6953 13001 6987
rect 13035 6984 13047 6987
rect 13998 6984 14004 6996
rect 13035 6956 14004 6984
rect 13035 6953 13047 6956
rect 12989 6947 13047 6953
rect 13998 6944 14004 6956
rect 14056 6944 14062 6996
rect 16022 6984 16028 6996
rect 14108 6956 16028 6984
rect 12342 6916 12348 6928
rect 11624 6888 12348 6916
rect 12342 6876 12348 6888
rect 12400 6876 12406 6928
rect 12802 6876 12808 6928
rect 12860 6916 12866 6928
rect 13173 6919 13231 6925
rect 13173 6916 13185 6919
rect 12860 6888 13185 6916
rect 12860 6876 12866 6888
rect 13173 6885 13185 6888
rect 13219 6885 13231 6919
rect 13173 6879 13231 6885
rect 6089 6851 6147 6857
rect 6089 6817 6101 6851
rect 6135 6848 6147 6851
rect 6917 6851 6975 6857
rect 6135 6820 6868 6848
rect 6135 6817 6147 6820
rect 6089 6811 6147 6817
rect 6840 6792 6868 6820
rect 6917 6817 6929 6851
rect 6963 6817 6975 6851
rect 6917 6811 6975 6817
rect 7558 6808 7564 6860
rect 7616 6848 7622 6860
rect 9033 6851 9091 6857
rect 9033 6848 9045 6851
rect 7616 6820 9045 6848
rect 7616 6808 7622 6820
rect 9033 6817 9045 6820
rect 9079 6817 9091 6851
rect 10321 6851 10379 6857
rect 10321 6848 10333 6851
rect 9033 6811 9091 6817
rect 9140 6820 10333 6848
rect 5813 6783 5871 6789
rect 5813 6749 5825 6783
rect 5859 6749 5871 6783
rect 5813 6743 5871 6749
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6749 5963 6783
rect 6178 6780 6184 6792
rect 6139 6752 6184 6780
rect 5905 6743 5963 6749
rect 4522 6672 4528 6724
rect 4580 6712 4586 6724
rect 5829 6712 5857 6743
rect 6178 6740 6184 6752
rect 6236 6740 6242 6792
rect 6822 6740 6828 6792
rect 6880 6780 6886 6792
rect 7193 6783 7251 6789
rect 7193 6780 7205 6783
rect 6880 6752 7205 6780
rect 6880 6740 6886 6752
rect 7193 6749 7205 6752
rect 7239 6749 7251 6783
rect 8202 6780 8208 6792
rect 7193 6743 7251 6749
rect 7300 6752 8208 6780
rect 7300 6712 7328 6752
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6780 8447 6783
rect 8662 6780 8668 6792
rect 8435 6752 8668 6780
rect 8435 6749 8447 6752
rect 8389 6743 8447 6749
rect 8662 6740 8668 6752
rect 8720 6740 8726 6792
rect 8754 6740 8760 6792
rect 8812 6780 8818 6792
rect 9140 6780 9168 6820
rect 10321 6817 10333 6820
rect 10367 6817 10379 6851
rect 14108 6848 14136 6956
rect 16022 6944 16028 6956
rect 16080 6944 16086 6996
rect 16298 6944 16304 6996
rect 16356 6984 16362 6996
rect 16393 6987 16451 6993
rect 16393 6984 16405 6987
rect 16356 6956 16405 6984
rect 16356 6944 16362 6956
rect 16393 6953 16405 6956
rect 16439 6953 16451 6987
rect 16393 6947 16451 6953
rect 16666 6944 16672 6996
rect 16724 6984 16730 6996
rect 16724 6956 19334 6984
rect 16724 6944 16730 6956
rect 18046 6876 18052 6928
rect 18104 6916 18110 6928
rect 18417 6919 18475 6925
rect 18417 6916 18429 6919
rect 18104 6888 18429 6916
rect 18104 6876 18110 6888
rect 18417 6885 18429 6888
rect 18463 6916 18475 6919
rect 18782 6916 18788 6928
rect 18463 6888 18788 6916
rect 18463 6885 18475 6888
rect 18417 6879 18475 6885
rect 18782 6876 18788 6888
rect 18840 6876 18846 6928
rect 10321 6811 10379 6817
rect 11348 6820 14136 6848
rect 8812 6752 9168 6780
rect 9217 6783 9275 6789
rect 8812 6740 8818 6752
rect 9217 6749 9229 6783
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 4580 6684 7328 6712
rect 4580 6672 4586 6684
rect 7926 6672 7932 6724
rect 7984 6712 7990 6724
rect 8941 6715 8999 6721
rect 8941 6712 8953 6715
rect 7984 6684 8953 6712
rect 7984 6672 7990 6684
rect 8941 6681 8953 6684
rect 8987 6681 8999 6715
rect 8941 6675 8999 6681
rect 9030 6672 9036 6724
rect 9088 6712 9094 6724
rect 9232 6712 9260 6743
rect 9398 6740 9404 6792
rect 9456 6780 9462 6792
rect 11348 6780 11376 6820
rect 15194 6808 15200 6860
rect 15252 6848 15258 6860
rect 19306 6848 19334 6956
rect 19904 6956 20944 6984
rect 19904 6848 19932 6956
rect 15252 6820 16252 6848
rect 19306 6820 19932 6848
rect 20916 6848 20944 6956
rect 21726 6944 21732 6996
rect 21784 6984 21790 6996
rect 25958 6984 25964 6996
rect 21784 6956 25964 6984
rect 21784 6944 21790 6956
rect 25958 6944 25964 6956
rect 26016 6944 26022 6996
rect 28721 6987 28779 6993
rect 28721 6953 28733 6987
rect 28767 6984 28779 6987
rect 29178 6984 29184 6996
rect 28767 6956 29184 6984
rect 28767 6953 28779 6956
rect 28721 6947 28779 6953
rect 29178 6944 29184 6956
rect 29236 6984 29242 6996
rect 33873 6987 33931 6993
rect 33873 6984 33885 6987
rect 29236 6956 33885 6984
rect 29236 6944 29242 6956
rect 33873 6953 33885 6956
rect 33919 6984 33931 6987
rect 34606 6984 34612 6996
rect 33919 6956 34612 6984
rect 33919 6953 33931 6956
rect 33873 6947 33931 6953
rect 34606 6944 34612 6956
rect 34664 6984 34670 6996
rect 34885 6987 34943 6993
rect 34885 6984 34897 6987
rect 34664 6956 34897 6984
rect 34664 6944 34670 6956
rect 34885 6953 34897 6956
rect 34931 6953 34943 6987
rect 34885 6947 34943 6953
rect 24026 6876 24032 6928
rect 24084 6916 24090 6928
rect 24394 6916 24400 6928
rect 24084 6888 24400 6916
rect 24084 6876 24090 6888
rect 24394 6876 24400 6888
rect 24452 6876 24458 6928
rect 24670 6876 24676 6928
rect 24728 6876 24734 6928
rect 24857 6919 24915 6925
rect 24857 6885 24869 6919
rect 24903 6916 24915 6919
rect 24946 6916 24952 6928
rect 24903 6888 24952 6916
rect 24903 6885 24915 6888
rect 24857 6879 24915 6885
rect 24946 6876 24952 6888
rect 25004 6876 25010 6928
rect 25038 6876 25044 6928
rect 25096 6916 25102 6928
rect 29454 6916 29460 6928
rect 25096 6888 29460 6916
rect 25096 6876 25102 6888
rect 29454 6876 29460 6888
rect 29512 6876 29518 6928
rect 32217 6919 32275 6925
rect 32217 6885 32229 6919
rect 32263 6885 32275 6919
rect 32217 6879 32275 6885
rect 35621 6919 35679 6925
rect 35621 6885 35633 6919
rect 35667 6885 35679 6919
rect 35621 6879 35679 6885
rect 21450 6848 21456 6860
rect 20916 6820 21456 6848
rect 15252 6808 15258 6820
rect 9456 6752 11376 6780
rect 9456 6740 9462 6752
rect 11974 6740 11980 6792
rect 12032 6780 12038 6792
rect 12897 6783 12955 6789
rect 12897 6780 12909 6783
rect 12032 6752 12909 6780
rect 12032 6740 12038 6752
rect 12897 6749 12909 6752
rect 12943 6749 12955 6783
rect 12897 6743 12955 6749
rect 12986 6740 12992 6792
rect 13044 6780 13050 6792
rect 13044 6752 13089 6780
rect 13044 6740 13050 6752
rect 13170 6740 13176 6792
rect 13228 6780 13234 6792
rect 13538 6780 13544 6792
rect 13228 6752 13544 6780
rect 13228 6740 13234 6752
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 14093 6783 14151 6789
rect 14093 6749 14105 6783
rect 14139 6780 14151 6783
rect 16114 6780 16120 6792
rect 14139 6752 14780 6780
rect 16075 6752 16120 6780
rect 14139 6749 14151 6752
rect 14093 6743 14151 6749
rect 14752 6724 14780 6752
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 16224 6789 16252 6820
rect 21450 6808 21456 6820
rect 21508 6808 21514 6860
rect 24302 6808 24308 6860
rect 24360 6848 24366 6860
rect 24688 6848 24716 6876
rect 29086 6848 29092 6860
rect 24360 6820 24716 6848
rect 24946 6820 29092 6848
rect 24360 6808 24366 6820
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6749 16267 6783
rect 16482 6780 16488 6792
rect 16443 6752 16488 6780
rect 16209 6743 16267 6749
rect 16482 6740 16488 6752
rect 16540 6740 16546 6792
rect 17037 6783 17095 6789
rect 17037 6749 17049 6783
rect 17083 6780 17095 6783
rect 17862 6780 17868 6792
rect 17083 6752 17868 6780
rect 17083 6749 17095 6752
rect 17037 6743 17095 6749
rect 10594 6721 10600 6724
rect 9088 6684 9260 6712
rect 9088 6672 9094 6684
rect 10588 6675 10600 6721
rect 10652 6712 10658 6724
rect 10652 6684 10688 6712
rect 10594 6672 10600 6675
rect 10652 6672 10658 6684
rect 10870 6672 10876 6724
rect 10928 6712 10934 6724
rect 10928 6684 12112 6712
rect 10928 6672 10934 6684
rect 2409 6647 2467 6653
rect 2409 6613 2421 6647
rect 2455 6644 2467 6647
rect 5626 6644 5632 6656
rect 2455 6616 5632 6644
rect 2455 6613 2467 6616
rect 2409 6607 2467 6613
rect 5626 6604 5632 6616
rect 5684 6604 5690 6656
rect 6454 6604 6460 6656
rect 6512 6644 6518 6656
rect 8205 6647 8263 6653
rect 8205 6644 8217 6647
rect 6512 6616 8217 6644
rect 6512 6604 6518 6616
rect 8205 6613 8217 6616
rect 8251 6613 8263 6647
rect 8205 6607 8263 6613
rect 9582 6604 9588 6656
rect 9640 6644 9646 6656
rect 10686 6644 10692 6656
rect 9640 6616 10692 6644
rect 9640 6604 9646 6616
rect 10686 6604 10692 6616
rect 10744 6604 10750 6656
rect 12084 6644 12112 6684
rect 12158 6672 12164 6724
rect 12216 6712 12222 6724
rect 12713 6715 12771 6721
rect 12713 6712 12725 6715
rect 12216 6684 12725 6712
rect 12216 6672 12222 6684
rect 12713 6681 12725 6684
rect 12759 6681 12771 6715
rect 14360 6715 14418 6721
rect 12713 6675 12771 6681
rect 13096 6684 14320 6712
rect 13096 6644 13124 6684
rect 12084 6616 13124 6644
rect 14292 6644 14320 6684
rect 14360 6681 14372 6715
rect 14406 6712 14418 6715
rect 14550 6712 14556 6724
rect 14406 6684 14556 6712
rect 14406 6681 14418 6684
rect 14360 6675 14418 6681
rect 14550 6672 14556 6684
rect 14608 6672 14614 6724
rect 14734 6672 14740 6724
rect 14792 6712 14798 6724
rect 17052 6712 17080 6743
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 19058 6740 19064 6792
rect 19116 6780 19122 6792
rect 19245 6783 19303 6789
rect 19245 6780 19257 6783
rect 19116 6752 19257 6780
rect 19116 6740 19122 6752
rect 19245 6749 19257 6752
rect 19291 6749 19303 6783
rect 19245 6743 19303 6749
rect 19334 6740 19340 6792
rect 19392 6780 19398 6792
rect 19889 6783 19947 6789
rect 19889 6780 19901 6783
rect 19392 6752 19901 6780
rect 19392 6740 19398 6752
rect 19889 6749 19901 6752
rect 19935 6780 19947 6783
rect 20622 6780 20628 6792
rect 19935 6752 20628 6780
rect 19935 6749 19947 6752
rect 19889 6743 19947 6749
rect 20622 6740 20628 6752
rect 20680 6780 20686 6792
rect 21818 6780 21824 6792
rect 20680 6752 21824 6780
rect 20680 6740 20686 6752
rect 21818 6740 21824 6752
rect 21876 6740 21882 6792
rect 22088 6783 22146 6789
rect 22088 6749 22100 6783
rect 22134 6780 22146 6783
rect 23750 6780 23756 6792
rect 22134 6752 23756 6780
rect 22134 6749 22146 6752
rect 22088 6743 22146 6749
rect 23750 6740 23756 6752
rect 23808 6740 23814 6792
rect 23845 6783 23903 6789
rect 23845 6749 23857 6783
rect 23891 6780 23903 6783
rect 24486 6780 24492 6792
rect 23891 6752 24492 6780
rect 23891 6749 23903 6752
rect 23845 6743 23903 6749
rect 24486 6740 24492 6752
rect 24544 6740 24550 6792
rect 24596 6789 24624 6820
rect 24581 6783 24639 6789
rect 24581 6749 24593 6783
rect 24627 6749 24639 6783
rect 24581 6743 24639 6749
rect 24673 6783 24731 6789
rect 24673 6749 24685 6783
rect 24719 6780 24731 6783
rect 24762 6780 24768 6792
rect 24719 6752 24768 6780
rect 24719 6749 24731 6752
rect 24673 6743 24731 6749
rect 24762 6740 24768 6752
rect 24820 6740 24826 6792
rect 24946 6789 24974 6820
rect 29086 6808 29092 6820
rect 29144 6808 29150 6860
rect 24946 6783 25007 6789
rect 24946 6749 24961 6783
rect 24995 6749 25007 6783
rect 25590 6780 25596 6792
rect 25551 6752 25596 6780
rect 24946 6748 25007 6749
rect 24949 6743 25007 6748
rect 25590 6740 25596 6752
rect 25648 6740 25654 6792
rect 26142 6740 26148 6792
rect 26200 6780 26206 6792
rect 26237 6783 26295 6789
rect 26237 6780 26249 6783
rect 26200 6752 26249 6780
rect 26200 6740 26206 6752
rect 26237 6749 26249 6752
rect 26283 6749 26295 6783
rect 26237 6743 26295 6749
rect 26326 6740 26332 6792
rect 26384 6780 26390 6792
rect 26881 6783 26939 6789
rect 26881 6780 26893 6783
rect 26384 6752 26893 6780
rect 26384 6740 26390 6752
rect 26881 6749 26893 6752
rect 26927 6749 26939 6783
rect 28074 6780 28080 6792
rect 28035 6752 28080 6780
rect 26881 6743 26939 6749
rect 28074 6740 28080 6752
rect 28132 6740 28138 6792
rect 29270 6780 29276 6792
rect 28757 6752 29276 6780
rect 20162 6721 20168 6724
rect 14792 6684 17080 6712
rect 17304 6715 17362 6721
rect 14792 6672 14798 6684
rect 17304 6681 17316 6715
rect 17350 6712 17362 6715
rect 20156 6712 20168 6721
rect 17350 6684 19472 6712
rect 20123 6684 20168 6712
rect 17350 6681 17362 6684
rect 17304 6675 17362 6681
rect 15102 6644 15108 6656
rect 14292 6616 15108 6644
rect 15102 6604 15108 6616
rect 15160 6604 15166 6656
rect 15194 6604 15200 6656
rect 15252 6644 15258 6656
rect 15473 6647 15531 6653
rect 15473 6644 15485 6647
rect 15252 6616 15485 6644
rect 15252 6604 15258 6616
rect 15473 6613 15485 6616
rect 15519 6613 15531 6647
rect 15930 6644 15936 6656
rect 15891 6616 15936 6644
rect 15473 6607 15531 6613
rect 15930 6604 15936 6616
rect 15988 6604 15994 6656
rect 16298 6604 16304 6656
rect 16356 6644 16362 6656
rect 19337 6647 19395 6653
rect 19337 6644 19349 6647
rect 16356 6616 19349 6644
rect 16356 6604 16362 6616
rect 19337 6613 19349 6616
rect 19383 6613 19395 6647
rect 19444 6644 19472 6684
rect 20156 6675 20168 6684
rect 20162 6672 20168 6675
rect 20220 6672 20226 6724
rect 23290 6712 23296 6724
rect 21284 6684 23296 6712
rect 21284 6656 21312 6684
rect 23290 6672 23296 6684
rect 23348 6672 23354 6724
rect 25130 6712 25136 6724
rect 23676 6684 25136 6712
rect 20714 6644 20720 6656
rect 19444 6616 20720 6644
rect 19337 6607 19395 6613
rect 20714 6604 20720 6616
rect 20772 6604 20778 6656
rect 21266 6644 21272 6656
rect 21179 6616 21272 6644
rect 21266 6604 21272 6616
rect 21324 6604 21330 6656
rect 21358 6604 21364 6656
rect 21416 6644 21422 6656
rect 23201 6647 23259 6653
rect 23201 6644 23213 6647
rect 21416 6616 23213 6644
rect 21416 6604 21422 6616
rect 23201 6613 23213 6616
rect 23247 6644 23259 6647
rect 23382 6644 23388 6656
rect 23247 6616 23388 6644
rect 23247 6613 23259 6616
rect 23201 6607 23259 6613
rect 23382 6604 23388 6616
rect 23440 6604 23446 6656
rect 23676 6653 23704 6684
rect 25130 6672 25136 6684
rect 25188 6672 25194 6724
rect 26510 6712 26516 6724
rect 26068 6684 26516 6712
rect 23661 6647 23719 6653
rect 23661 6613 23673 6647
rect 23707 6613 23719 6647
rect 24394 6644 24400 6656
rect 24355 6616 24400 6644
rect 23661 6607 23719 6613
rect 24394 6604 24400 6616
rect 24452 6604 24458 6656
rect 25222 6604 25228 6656
rect 25280 6644 25286 6656
rect 26068 6653 26096 6684
rect 26510 6672 26516 6684
rect 26568 6672 26574 6724
rect 28534 6712 28540 6724
rect 28495 6684 28540 6712
rect 28534 6672 28540 6684
rect 28592 6672 28598 6724
rect 28757 6721 28785 6752
rect 29270 6740 29276 6752
rect 29328 6740 29334 6792
rect 29730 6780 29736 6792
rect 29691 6752 29736 6780
rect 29730 6740 29736 6752
rect 29788 6780 29794 6792
rect 29788 6752 30144 6780
rect 29788 6740 29794 6752
rect 28742 6715 28800 6721
rect 28742 6681 28754 6715
rect 28788 6681 28800 6715
rect 29822 6712 29828 6724
rect 28742 6675 28800 6681
rect 28828 6684 29828 6712
rect 25409 6647 25467 6653
rect 25409 6644 25421 6647
rect 25280 6616 25421 6644
rect 25280 6604 25286 6616
rect 25409 6613 25421 6616
rect 25455 6613 25467 6647
rect 25409 6607 25467 6613
rect 26053 6647 26111 6653
rect 26053 6613 26065 6647
rect 26099 6613 26111 6647
rect 26053 6607 26111 6613
rect 26418 6604 26424 6656
rect 26476 6644 26482 6656
rect 26697 6647 26755 6653
rect 26697 6644 26709 6647
rect 26476 6616 26709 6644
rect 26476 6604 26482 6616
rect 26697 6613 26709 6616
rect 26743 6613 26755 6647
rect 26697 6607 26755 6613
rect 27893 6647 27951 6653
rect 27893 6613 27905 6647
rect 27939 6644 27951 6647
rect 28828 6644 28856 6684
rect 29822 6672 29828 6684
rect 29880 6672 29886 6724
rect 30006 6721 30012 6724
rect 30000 6712 30012 6721
rect 29967 6684 30012 6712
rect 30000 6675 30012 6684
rect 30006 6672 30012 6675
rect 30064 6672 30070 6724
rect 30116 6712 30144 6752
rect 31754 6740 31760 6792
rect 31812 6780 31818 6792
rect 31812 6752 31857 6780
rect 31812 6740 31818 6752
rect 32122 6712 32128 6724
rect 30116 6684 32128 6712
rect 32122 6672 32128 6684
rect 32180 6672 32186 6724
rect 32232 6712 32260 6879
rect 32490 6808 32496 6860
rect 32548 6848 32554 6860
rect 35636 6848 35664 6879
rect 37550 6848 37556 6860
rect 32548 6820 34100 6848
rect 35636 6820 37556 6848
rect 32548 6808 32554 6820
rect 34072 6792 34100 6820
rect 37550 6808 37556 6820
rect 37608 6808 37614 6860
rect 32306 6740 32312 6792
rect 32364 6780 32370 6792
rect 32401 6783 32459 6789
rect 32401 6780 32413 6783
rect 32364 6752 32413 6780
rect 32364 6740 32370 6752
rect 32401 6749 32413 6752
rect 32447 6749 32459 6783
rect 32401 6743 32459 6749
rect 32766 6740 32772 6792
rect 32824 6780 32830 6792
rect 33413 6783 33471 6789
rect 33413 6780 33425 6783
rect 32824 6752 33425 6780
rect 32824 6740 32830 6752
rect 33413 6749 33425 6752
rect 33459 6749 33471 6783
rect 34054 6780 34060 6792
rect 34015 6752 34060 6780
rect 33413 6743 33471 6749
rect 34054 6740 34060 6752
rect 34112 6740 34118 6792
rect 35802 6780 35808 6792
rect 35763 6752 35808 6780
rect 35802 6740 35808 6752
rect 35860 6740 35866 6792
rect 36449 6783 36507 6789
rect 36449 6749 36461 6783
rect 36495 6749 36507 6783
rect 36449 6743 36507 6749
rect 33502 6712 33508 6724
rect 32232 6684 33508 6712
rect 33502 6672 33508 6684
rect 33560 6672 33566 6724
rect 34698 6712 34704 6724
rect 34659 6684 34704 6712
rect 34698 6672 34704 6684
rect 34756 6672 34762 6724
rect 36464 6712 36492 6743
rect 35084 6684 36492 6712
rect 27939 6616 28856 6644
rect 28905 6647 28963 6653
rect 27939 6613 27951 6616
rect 27893 6607 27951 6613
rect 28905 6613 28917 6647
rect 28951 6644 28963 6647
rect 30466 6644 30472 6656
rect 28951 6616 30472 6644
rect 28951 6613 28963 6616
rect 28905 6607 28963 6613
rect 30466 6604 30472 6616
rect 30524 6604 30530 6656
rect 31113 6647 31171 6653
rect 31113 6613 31125 6647
rect 31159 6644 31171 6647
rect 31202 6644 31208 6656
rect 31159 6616 31208 6644
rect 31159 6613 31171 6616
rect 31113 6607 31171 6613
rect 31202 6604 31208 6616
rect 31260 6604 31266 6656
rect 31573 6647 31631 6653
rect 31573 6613 31585 6647
rect 31619 6644 31631 6647
rect 32858 6644 32864 6656
rect 31619 6616 32864 6644
rect 31619 6613 31631 6616
rect 31573 6607 31631 6613
rect 32858 6604 32864 6616
rect 32916 6604 32922 6656
rect 33229 6647 33287 6653
rect 33229 6613 33241 6647
rect 33275 6644 33287 6647
rect 33870 6644 33876 6656
rect 33275 6616 33876 6644
rect 33275 6613 33287 6616
rect 33229 6607 33287 6613
rect 33870 6604 33876 6616
rect 33928 6604 33934 6656
rect 34882 6604 34888 6656
rect 34940 6653 34946 6656
rect 35084 6653 35112 6684
rect 34940 6647 34959 6653
rect 34947 6613 34959 6647
rect 34940 6607 34959 6613
rect 35069 6647 35127 6653
rect 35069 6613 35081 6647
rect 35115 6613 35127 6647
rect 35069 6607 35127 6613
rect 36265 6647 36323 6653
rect 36265 6613 36277 6647
rect 36311 6644 36323 6647
rect 37642 6644 37648 6656
rect 36311 6616 37648 6644
rect 36311 6613 36323 6616
rect 36265 6607 36323 6613
rect 34940 6604 34946 6607
rect 37642 6604 37648 6616
rect 37700 6604 37706 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 1762 6440 1768 6452
rect 1723 6412 1768 6440
rect 1762 6400 1768 6412
rect 1820 6400 1826 6452
rect 3053 6443 3111 6449
rect 3053 6409 3065 6443
rect 3099 6409 3111 6443
rect 3053 6403 3111 6409
rect 3697 6443 3755 6449
rect 3697 6409 3709 6443
rect 3743 6440 3755 6443
rect 3878 6440 3884 6452
rect 3743 6412 3884 6440
rect 3743 6409 3755 6412
rect 3697 6403 3755 6409
rect 3068 6372 3096 6403
rect 3878 6400 3884 6412
rect 3936 6400 3942 6452
rect 3970 6400 3976 6452
rect 4028 6440 4034 6452
rect 4706 6440 4712 6452
rect 4028 6412 4712 6440
rect 4028 6400 4034 6412
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 5813 6443 5871 6449
rect 5813 6409 5825 6443
rect 5859 6440 5871 6443
rect 6086 6440 6092 6452
rect 5859 6412 6092 6440
rect 5859 6409 5871 6412
rect 5813 6403 5871 6409
rect 6086 6400 6092 6412
rect 6144 6400 6150 6452
rect 6472 6412 9076 6440
rect 4430 6372 4436 6384
rect 3068 6344 4436 6372
rect 4430 6332 4436 6344
rect 4488 6332 4494 6384
rect 5445 6375 5503 6381
rect 5445 6341 5457 6375
rect 5491 6372 5503 6375
rect 6365 6375 6423 6381
rect 6365 6372 6377 6375
rect 5491 6344 6377 6372
rect 5491 6341 5503 6344
rect 5445 6335 5503 6341
rect 6365 6341 6377 6344
rect 6411 6341 6423 6375
rect 6365 6335 6423 6341
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 2409 6307 2467 6313
rect 2409 6273 2421 6307
rect 2455 6273 2467 6307
rect 2409 6267 2467 6273
rect 2685 6307 2743 6313
rect 2685 6273 2697 6307
rect 2731 6304 2743 6307
rect 3237 6307 3295 6313
rect 3237 6304 3249 6307
rect 2731 6276 3249 6304
rect 2731 6273 2743 6276
rect 2685 6267 2743 6273
rect 3237 6273 3249 6276
rect 3283 6273 3295 6307
rect 3878 6304 3884 6316
rect 3839 6276 3884 6304
rect 3237 6267 3295 6273
rect 1964 6168 1992 6267
rect 2424 6236 2452 6267
rect 2774 6236 2780 6248
rect 2424 6208 2780 6236
rect 2774 6196 2780 6208
rect 2832 6196 2838 6248
rect 3252 6236 3280 6267
rect 3878 6264 3884 6276
rect 3936 6264 3942 6316
rect 4522 6304 4528 6316
rect 4483 6276 4528 6304
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 4614 6264 4620 6316
rect 4672 6304 4678 6316
rect 4672 6276 4717 6304
rect 4672 6264 4678 6276
rect 4798 6264 4804 6316
rect 4856 6304 4862 6316
rect 4893 6307 4951 6313
rect 4893 6304 4905 6307
rect 4856 6276 4905 6304
rect 4856 6264 4862 6276
rect 4893 6273 4905 6276
rect 4939 6273 4951 6307
rect 4893 6267 4951 6273
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 5629 6307 5687 6313
rect 5629 6304 5641 6307
rect 5592 6276 5641 6304
rect 5592 6264 5598 6276
rect 5629 6273 5641 6276
rect 5675 6273 5687 6307
rect 6472 6304 6500 6412
rect 7282 6372 7288 6384
rect 6564 6344 7288 6372
rect 6564 6313 6592 6344
rect 7282 6332 7288 6344
rect 7340 6332 7346 6384
rect 7374 6332 7380 6384
rect 7432 6372 7438 6384
rect 7653 6375 7711 6381
rect 7653 6372 7665 6375
rect 7432 6344 7665 6372
rect 7432 6332 7438 6344
rect 7653 6341 7665 6344
rect 7699 6372 7711 6375
rect 8478 6372 8484 6384
rect 7699 6344 8484 6372
rect 7699 6341 7711 6344
rect 7653 6335 7711 6341
rect 8478 6332 8484 6344
rect 8536 6332 8542 6384
rect 8573 6375 8631 6381
rect 8573 6341 8585 6375
rect 8619 6372 8631 6375
rect 8938 6372 8944 6384
rect 8619 6344 8944 6372
rect 8619 6341 8631 6344
rect 8573 6335 8631 6341
rect 8938 6332 8944 6344
rect 8996 6332 9002 6384
rect 9048 6372 9076 6412
rect 9490 6400 9496 6452
rect 9548 6440 9554 6452
rect 9585 6443 9643 6449
rect 9585 6440 9597 6443
rect 9548 6412 9597 6440
rect 9548 6400 9554 6412
rect 9585 6409 9597 6412
rect 9631 6409 9643 6443
rect 9585 6403 9643 6409
rect 10134 6400 10140 6452
rect 10192 6400 10198 6452
rect 10594 6440 10600 6452
rect 10555 6412 10600 6440
rect 10594 6400 10600 6412
rect 10652 6400 10658 6452
rect 10686 6400 10692 6452
rect 10744 6440 10750 6452
rect 10744 6412 12020 6440
rect 10744 6400 10750 6412
rect 10152 6372 10180 6400
rect 9048 6344 9674 6372
rect 5629 6267 5687 6273
rect 5736 6276 6500 6304
rect 6549 6307 6607 6313
rect 5736 6236 5764 6276
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6638 6264 6644 6316
rect 6696 6304 6702 6316
rect 6917 6307 6975 6313
rect 6696 6276 6741 6304
rect 6696 6264 6702 6276
rect 6917 6273 6929 6307
rect 6963 6273 6975 6307
rect 6917 6267 6975 6273
rect 3252 6208 5764 6236
rect 5810 6196 5816 6248
rect 5868 6236 5874 6248
rect 6932 6236 6960 6267
rect 7006 6264 7012 6316
rect 7064 6304 7070 6316
rect 7469 6307 7527 6313
rect 7469 6304 7481 6307
rect 7064 6276 7481 6304
rect 7064 6264 7070 6276
rect 7469 6273 7481 6276
rect 7515 6304 7527 6307
rect 8662 6304 8668 6316
rect 7515 6276 8668 6304
rect 7515 6273 7527 6276
rect 7469 6267 7527 6273
rect 8662 6264 8668 6276
rect 8720 6264 8726 6316
rect 8757 6307 8815 6313
rect 8757 6273 8769 6307
rect 8803 6273 8815 6307
rect 8757 6267 8815 6273
rect 5868 6208 6960 6236
rect 5868 6196 5874 6208
rect 8386 6196 8392 6248
rect 8444 6236 8450 6248
rect 8772 6236 8800 6267
rect 8444 6208 8800 6236
rect 8444 6196 8450 6208
rect 8846 6196 8852 6248
rect 8904 6236 8910 6248
rect 8941 6239 8999 6245
rect 8941 6236 8953 6239
rect 8904 6208 8953 6236
rect 8904 6196 8910 6208
rect 8941 6205 8953 6208
rect 8987 6205 8999 6239
rect 9646 6236 9674 6344
rect 9784 6344 10180 6372
rect 9784 6313 9812 6344
rect 10226 6332 10232 6384
rect 10284 6372 10290 6384
rect 11517 6375 11575 6381
rect 11517 6372 11529 6375
rect 10284 6344 11529 6372
rect 10284 6332 10290 6344
rect 11517 6341 11529 6344
rect 11563 6341 11575 6375
rect 11992 6372 12020 6412
rect 12710 6400 12716 6452
rect 12768 6440 12774 6452
rect 12805 6443 12863 6449
rect 12805 6440 12817 6443
rect 12768 6412 12817 6440
rect 12768 6400 12774 6412
rect 12805 6409 12817 6412
rect 12851 6409 12863 6443
rect 12805 6403 12863 6409
rect 12986 6400 12992 6452
rect 13044 6440 13050 6452
rect 14277 6443 14335 6449
rect 14277 6440 14289 6443
rect 13044 6412 14289 6440
rect 13044 6400 13050 6412
rect 14277 6409 14289 6412
rect 14323 6409 14335 6443
rect 14277 6403 14335 6409
rect 15102 6400 15108 6452
rect 15160 6440 15166 6452
rect 16482 6440 16488 6452
rect 15160 6412 16488 6440
rect 15160 6400 15166 6412
rect 16482 6400 16488 6412
rect 16540 6400 16546 6452
rect 24670 6440 24676 6452
rect 16592 6412 24676 6440
rect 13170 6372 13176 6384
rect 11517 6335 11575 6341
rect 11624 6344 11928 6372
rect 11992 6344 13176 6372
rect 9769 6307 9827 6313
rect 9769 6273 9781 6307
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 9861 6307 9919 6313
rect 9861 6273 9873 6307
rect 9907 6304 9919 6307
rect 9950 6304 9956 6316
rect 9907 6276 9956 6304
rect 9907 6273 9919 6276
rect 9861 6267 9919 6273
rect 9950 6264 9956 6276
rect 10008 6264 10014 6316
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6304 10195 6307
rect 10502 6304 10508 6316
rect 10183 6276 10508 6304
rect 10183 6273 10195 6276
rect 10137 6267 10195 6273
rect 10502 6264 10508 6276
rect 10560 6264 10566 6316
rect 10778 6304 10784 6316
rect 10739 6276 10784 6304
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 11624 6304 11652 6344
rect 10888 6276 11652 6304
rect 10888 6236 10916 6276
rect 11698 6264 11704 6316
rect 11756 6304 11762 6316
rect 11793 6307 11851 6313
rect 11793 6304 11805 6307
rect 11756 6276 11805 6304
rect 11756 6264 11762 6276
rect 11793 6273 11805 6276
rect 11839 6273 11851 6307
rect 11900 6304 11928 6344
rect 13170 6332 13176 6344
rect 13228 6332 13234 6384
rect 13817 6375 13875 6381
rect 13817 6372 13829 6375
rect 13280 6344 13829 6372
rect 13280 6316 13308 6344
rect 13817 6341 13829 6344
rect 13863 6341 13875 6375
rect 13817 6335 13875 6341
rect 15286 6332 15292 6384
rect 15344 6372 15350 6384
rect 16592 6372 16620 6412
rect 24670 6400 24676 6412
rect 24728 6400 24734 6452
rect 31846 6440 31852 6452
rect 24872 6412 31852 6440
rect 15344 6344 16620 6372
rect 18408 6375 18466 6381
rect 15344 6332 15350 6344
rect 18408 6341 18420 6375
rect 18454 6372 18466 6375
rect 18874 6372 18880 6384
rect 18454 6344 18880 6372
rect 18454 6341 18466 6344
rect 18408 6335 18466 6341
rect 18874 6332 18880 6344
rect 18932 6332 18938 6384
rect 19242 6332 19248 6384
rect 19300 6372 19306 6384
rect 20162 6372 20168 6384
rect 19300 6344 20168 6372
rect 19300 6332 19306 6344
rect 20162 6332 20168 6344
rect 20220 6332 20226 6384
rect 21174 6332 21180 6384
rect 21232 6372 21238 6384
rect 24872 6372 24900 6412
rect 31846 6400 31852 6412
rect 31904 6400 31910 6452
rect 36173 6443 36231 6449
rect 36173 6409 36185 6443
rect 36219 6440 36231 6443
rect 36446 6440 36452 6452
rect 36219 6412 36452 6440
rect 36219 6409 36231 6412
rect 36173 6403 36231 6409
rect 36446 6400 36452 6412
rect 36504 6400 36510 6452
rect 26234 6372 26240 6384
rect 21232 6344 24900 6372
rect 24964 6344 26240 6372
rect 21232 6332 21238 6344
rect 12342 6304 12348 6316
rect 11900 6276 12348 6304
rect 11793 6267 11851 6273
rect 12342 6264 12348 6276
rect 12400 6264 12406 6316
rect 12986 6304 12992 6316
rect 12947 6276 12992 6304
rect 12986 6264 12992 6276
rect 13044 6264 13050 6316
rect 13081 6307 13139 6313
rect 13081 6273 13093 6307
rect 13127 6304 13139 6307
rect 13262 6304 13268 6316
rect 13127 6276 13268 6304
rect 13127 6273 13139 6276
rect 13081 6267 13139 6273
rect 13262 6264 13268 6276
rect 13320 6264 13326 6316
rect 13357 6307 13415 6313
rect 13357 6273 13369 6307
rect 13403 6273 13415 6307
rect 14090 6304 14096 6316
rect 14051 6276 14096 6304
rect 13357 6267 13415 6273
rect 11606 6236 11612 6248
rect 9646 6208 10916 6236
rect 11567 6208 11612 6236
rect 8941 6199 8999 6205
rect 11606 6196 11612 6208
rect 11664 6196 11670 6248
rect 13372 6236 13400 6267
rect 14090 6264 14096 6276
rect 14148 6264 14154 6316
rect 14734 6304 14740 6316
rect 14695 6276 14740 6304
rect 14734 6264 14740 6276
rect 14792 6264 14798 6316
rect 15010 6313 15016 6316
rect 15004 6304 15016 6313
rect 14971 6276 15016 6304
rect 15004 6267 15016 6276
rect 15010 6264 15016 6267
rect 15068 6264 15074 6316
rect 17218 6264 17224 6316
rect 17276 6304 17282 6316
rect 19978 6304 19984 6316
rect 17276 6276 19984 6304
rect 17276 6264 17282 6276
rect 19978 6264 19984 6276
rect 20036 6264 20042 6316
rect 20438 6304 20444 6316
rect 20399 6276 20444 6304
rect 20438 6264 20444 6276
rect 20496 6264 20502 6316
rect 21634 6304 21640 6316
rect 20548 6276 21640 6304
rect 11808 6208 13400 6236
rect 1964 6140 2774 6168
rect 2225 6103 2283 6109
rect 2225 6069 2237 6103
rect 2271 6100 2283 6103
rect 2406 6100 2412 6112
rect 2271 6072 2412 6100
rect 2271 6069 2283 6072
rect 2225 6063 2283 6069
rect 2406 6060 2412 6072
rect 2464 6060 2470 6112
rect 2746 6100 2774 6140
rect 2866 6128 2872 6180
rect 2924 6168 2930 6180
rect 2924 6140 10180 6168
rect 2924 6128 2930 6140
rect 3326 6100 3332 6112
rect 2746 6072 3332 6100
rect 3326 6060 3332 6072
rect 3384 6060 3390 6112
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 4341 6103 4399 6109
rect 4341 6100 4353 6103
rect 4120 6072 4353 6100
rect 4120 6060 4126 6072
rect 4341 6069 4353 6072
rect 4387 6069 4399 6103
rect 4341 6063 4399 6069
rect 4801 6103 4859 6109
rect 4801 6069 4813 6103
rect 4847 6100 4859 6103
rect 5534 6100 5540 6112
rect 4847 6072 5540 6100
rect 4847 6069 4859 6072
rect 4801 6063 4859 6069
rect 5534 6060 5540 6072
rect 5592 6100 5598 6112
rect 6822 6100 6828 6112
rect 5592 6072 6828 6100
rect 5592 6060 5598 6072
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 7742 6060 7748 6112
rect 7800 6100 7806 6112
rect 9582 6100 9588 6112
rect 7800 6072 9588 6100
rect 7800 6060 7806 6072
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 10042 6100 10048 6112
rect 10003 6072 10048 6100
rect 10042 6060 10048 6072
rect 10100 6060 10106 6112
rect 10152 6100 10180 6140
rect 10226 6128 10232 6180
rect 10284 6168 10290 6180
rect 11808 6168 11836 6208
rect 13814 6196 13820 6248
rect 13872 6236 13878 6248
rect 13909 6239 13967 6245
rect 13909 6236 13921 6239
rect 13872 6208 13921 6236
rect 13872 6196 13878 6208
rect 13909 6205 13921 6208
rect 13955 6205 13967 6239
rect 13909 6199 13967 6205
rect 16114 6196 16120 6248
rect 16172 6236 16178 6248
rect 16669 6239 16727 6245
rect 16669 6236 16681 6239
rect 16172 6208 16681 6236
rect 16172 6196 16178 6208
rect 16669 6205 16681 6208
rect 16715 6205 16727 6239
rect 16669 6199 16727 6205
rect 16945 6239 17003 6245
rect 16945 6205 16957 6239
rect 16991 6236 17003 6239
rect 17678 6236 17684 6248
rect 16991 6208 17684 6236
rect 16991 6205 17003 6208
rect 16945 6199 17003 6205
rect 17678 6196 17684 6208
rect 17736 6196 17742 6248
rect 18141 6239 18199 6245
rect 18141 6205 18153 6239
rect 18187 6205 18199 6239
rect 18141 6199 18199 6205
rect 11974 6168 11980 6180
rect 10284 6140 11836 6168
rect 11935 6140 11980 6168
rect 10284 6128 10290 6140
rect 11974 6128 11980 6140
rect 12032 6128 12038 6180
rect 13265 6171 13323 6177
rect 13265 6137 13277 6171
rect 13311 6168 13323 6171
rect 13311 6140 13952 6168
rect 13311 6137 13323 6140
rect 13265 6131 13323 6137
rect 13924 6112 13952 6140
rect 11422 6100 11428 6112
rect 10152 6072 11428 6100
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 11514 6060 11520 6112
rect 11572 6100 11578 6112
rect 11572 6072 11617 6100
rect 11572 6060 11578 6072
rect 13354 6060 13360 6112
rect 13412 6100 13418 6112
rect 13817 6103 13875 6109
rect 13817 6100 13829 6103
rect 13412 6072 13829 6100
rect 13412 6060 13418 6072
rect 13817 6069 13829 6072
rect 13863 6069 13875 6103
rect 13817 6063 13875 6069
rect 13906 6060 13912 6112
rect 13964 6060 13970 6112
rect 16114 6100 16120 6112
rect 16075 6072 16120 6100
rect 16114 6060 16120 6072
rect 16172 6060 16178 6112
rect 18156 6100 18184 6199
rect 19242 6196 19248 6248
rect 19300 6236 19306 6248
rect 20548 6236 20576 6276
rect 21634 6264 21640 6276
rect 21692 6264 21698 6316
rect 21818 6264 21824 6316
rect 21876 6304 21882 6316
rect 22278 6304 22284 6316
rect 21876 6276 22284 6304
rect 21876 6264 21882 6276
rect 22278 6264 22284 6276
rect 22336 6264 22342 6316
rect 22548 6307 22606 6313
rect 22548 6273 22560 6307
rect 22594 6304 22606 6307
rect 22830 6304 22836 6316
rect 22594 6276 22836 6304
rect 22594 6273 22606 6276
rect 22548 6267 22606 6273
rect 22830 6264 22836 6276
rect 22888 6264 22894 6316
rect 24121 6307 24179 6313
rect 24121 6273 24133 6307
rect 24167 6273 24179 6307
rect 24302 6304 24308 6316
rect 24263 6276 24308 6304
rect 24121 6267 24179 6273
rect 19300 6208 20576 6236
rect 20717 6239 20775 6245
rect 19300 6196 19306 6208
rect 20717 6205 20729 6239
rect 20763 6236 20775 6239
rect 21450 6236 21456 6248
rect 20763 6208 21456 6236
rect 20763 6205 20775 6208
rect 20717 6199 20775 6205
rect 21450 6196 21456 6208
rect 21508 6196 21514 6248
rect 24136 6236 24164 6267
rect 24302 6264 24308 6276
rect 24360 6264 24366 6316
rect 24964 6313 24992 6344
rect 26234 6332 26240 6344
rect 26292 6372 26298 6384
rect 29730 6372 29736 6384
rect 26292 6344 27108 6372
rect 26292 6332 26298 6344
rect 27080 6316 27108 6344
rect 27448 6344 29736 6372
rect 24949 6307 25007 6313
rect 24949 6273 24961 6307
rect 24995 6273 25007 6307
rect 24949 6267 25007 6273
rect 25216 6307 25274 6313
rect 25216 6273 25228 6307
rect 25262 6304 25274 6307
rect 25498 6304 25504 6316
rect 25262 6276 25504 6304
rect 25262 6273 25274 6276
rect 25216 6267 25274 6273
rect 25498 6264 25504 6276
rect 25556 6264 25562 6316
rect 27062 6264 27068 6316
rect 27120 6304 27126 6316
rect 27448 6313 27476 6344
rect 27433 6307 27491 6313
rect 27433 6304 27445 6307
rect 27120 6276 27445 6304
rect 27120 6264 27126 6276
rect 27433 6273 27445 6276
rect 27479 6273 27491 6307
rect 27433 6267 27491 6273
rect 27522 6264 27528 6316
rect 27580 6264 27586 6316
rect 27700 6307 27758 6313
rect 27700 6273 27712 6307
rect 27746 6304 27758 6307
rect 28994 6304 29000 6316
rect 27746 6276 29000 6304
rect 27746 6273 27758 6276
rect 27700 6267 27758 6273
rect 28994 6264 29000 6276
rect 29052 6264 29058 6316
rect 29288 6313 29316 6344
rect 29730 6332 29736 6344
rect 29788 6332 29794 6384
rect 29822 6332 29828 6384
rect 29880 6372 29886 6384
rect 32950 6372 32956 6384
rect 29880 6344 31340 6372
rect 29880 6332 29886 6344
rect 29273 6307 29331 6313
rect 29273 6273 29285 6307
rect 29319 6273 29331 6307
rect 29273 6267 29331 6273
rect 29540 6307 29598 6313
rect 29540 6273 29552 6307
rect 29586 6304 29598 6307
rect 30374 6304 30380 6316
rect 29586 6276 30380 6304
rect 29586 6273 29598 6276
rect 29540 6267 29598 6273
rect 30374 6264 30380 6276
rect 30432 6264 30438 6316
rect 31312 6313 31340 6344
rect 32140 6344 32956 6372
rect 31297 6307 31355 6313
rect 31297 6273 31309 6307
rect 31343 6273 31355 6307
rect 31297 6267 31355 6273
rect 24854 6236 24860 6248
rect 24136 6208 24860 6236
rect 24854 6196 24860 6208
rect 24912 6196 24918 6248
rect 27540 6236 27568 6264
rect 32140 6248 32168 6344
rect 32950 6332 32956 6344
rect 33008 6372 33014 6384
rect 34232 6375 34290 6381
rect 33008 6344 34008 6372
rect 33008 6332 33014 6344
rect 32398 6313 32404 6316
rect 32392 6304 32404 6313
rect 32359 6276 32404 6304
rect 32392 6267 32404 6276
rect 32398 6264 32404 6267
rect 32456 6264 32462 6316
rect 33980 6313 34008 6344
rect 34232 6341 34244 6375
rect 34278 6372 34290 6375
rect 34790 6372 34796 6384
rect 34278 6344 34796 6372
rect 34278 6341 34290 6344
rect 34232 6335 34290 6341
rect 34790 6332 34796 6344
rect 34848 6332 34854 6384
rect 35805 6375 35863 6381
rect 35805 6372 35817 6375
rect 35360 6344 35817 6372
rect 33965 6307 34023 6313
rect 33965 6273 33977 6307
rect 34011 6273 34023 6307
rect 33965 6267 34023 6273
rect 32122 6236 32128 6248
rect 26068 6208 27568 6236
rect 32083 6208 32128 6236
rect 19150 6128 19156 6180
rect 19208 6168 19214 6180
rect 19521 6171 19579 6177
rect 19521 6168 19533 6171
rect 19208 6140 19533 6168
rect 19208 6128 19214 6140
rect 19521 6137 19533 6140
rect 19567 6137 19579 6171
rect 19521 6131 19579 6137
rect 23474 6128 23480 6180
rect 23532 6168 23538 6180
rect 23661 6171 23719 6177
rect 23661 6168 23673 6171
rect 23532 6140 23673 6168
rect 23532 6128 23538 6140
rect 23661 6137 23673 6140
rect 23707 6137 23719 6171
rect 24762 6168 24768 6180
rect 23661 6131 23719 6137
rect 24412 6140 24768 6168
rect 19334 6100 19340 6112
rect 18156 6072 19340 6100
rect 19334 6060 19340 6072
rect 19392 6060 19398 6112
rect 19610 6060 19616 6112
rect 19668 6100 19674 6112
rect 24412 6100 24440 6140
rect 24762 6128 24768 6140
rect 24820 6128 24826 6180
rect 19668 6072 24440 6100
rect 24489 6103 24547 6109
rect 19668 6060 19674 6072
rect 24489 6069 24501 6103
rect 24535 6100 24547 6103
rect 26068 6100 26096 6208
rect 32122 6196 32128 6208
rect 32180 6196 32186 6248
rect 26142 6128 26148 6180
rect 26200 6168 26206 6180
rect 26200 6140 27476 6168
rect 26200 6128 26206 6140
rect 24535 6072 26096 6100
rect 26329 6103 26387 6109
rect 24535 6069 24547 6072
rect 24489 6063 24547 6069
rect 26329 6069 26341 6103
rect 26375 6100 26387 6103
rect 27246 6100 27252 6112
rect 26375 6072 27252 6100
rect 26375 6069 26387 6072
rect 26329 6063 26387 6069
rect 27246 6060 27252 6072
rect 27304 6060 27310 6112
rect 27448 6100 27476 6140
rect 35360 6112 35388 6344
rect 35805 6341 35817 6344
rect 35851 6341 35863 6375
rect 35805 6335 35863 6341
rect 35894 6332 35900 6384
rect 35952 6372 35958 6384
rect 36005 6375 36063 6381
rect 36005 6372 36017 6375
rect 35952 6344 36017 6372
rect 35952 6332 35958 6344
rect 36005 6341 36017 6344
rect 36051 6341 36063 6375
rect 36005 6335 36063 6341
rect 37274 6264 37280 6316
rect 37332 6304 37338 6316
rect 37461 6307 37519 6313
rect 37461 6304 37473 6307
rect 37332 6276 37473 6304
rect 37332 6264 37338 6276
rect 37461 6273 37473 6276
rect 37507 6273 37519 6307
rect 37461 6267 37519 6273
rect 27798 6100 27804 6112
rect 27448 6072 27804 6100
rect 27798 6060 27804 6072
rect 27856 6060 27862 6112
rect 28534 6060 28540 6112
rect 28592 6100 28598 6112
rect 28813 6103 28871 6109
rect 28813 6100 28825 6103
rect 28592 6072 28825 6100
rect 28592 6060 28598 6072
rect 28813 6069 28825 6072
rect 28859 6069 28871 6103
rect 28813 6063 28871 6069
rect 29454 6060 29460 6112
rect 29512 6100 29518 6112
rect 30653 6103 30711 6109
rect 30653 6100 30665 6103
rect 29512 6072 30665 6100
rect 29512 6060 29518 6072
rect 30653 6069 30665 6072
rect 30699 6069 30711 6103
rect 30653 6063 30711 6069
rect 31113 6103 31171 6109
rect 31113 6069 31125 6103
rect 31159 6100 31171 6103
rect 31846 6100 31852 6112
rect 31159 6072 31852 6100
rect 31159 6069 31171 6072
rect 31113 6063 31171 6069
rect 31846 6060 31852 6072
rect 31904 6060 31910 6112
rect 33042 6060 33048 6112
rect 33100 6100 33106 6112
rect 33505 6103 33563 6109
rect 33505 6100 33517 6103
rect 33100 6072 33517 6100
rect 33100 6060 33106 6072
rect 33505 6069 33517 6072
rect 33551 6069 33563 6103
rect 35342 6100 35348 6112
rect 35303 6072 35348 6100
rect 33505 6063 33563 6069
rect 35342 6060 35348 6072
rect 35400 6060 35406 6112
rect 35986 6100 35992 6112
rect 35947 6072 35992 6100
rect 35986 6060 35992 6072
rect 36044 6060 36050 6112
rect 37277 6103 37335 6109
rect 37277 6069 37289 6103
rect 37323 6100 37335 6103
rect 37918 6100 37924 6112
rect 37323 6072 37924 6100
rect 37323 6069 37335 6072
rect 37277 6063 37335 6069
rect 37918 6060 37924 6072
rect 37976 6060 37982 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 1627 5868 3004 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 2976 5760 3004 5868
rect 3878 5856 3884 5908
rect 3936 5896 3942 5908
rect 4525 5899 4583 5905
rect 4525 5896 4537 5899
rect 3936 5868 4537 5896
rect 3936 5856 3942 5868
rect 4525 5865 4537 5868
rect 4571 5865 4583 5899
rect 4525 5859 4583 5865
rect 4614 5856 4620 5908
rect 4672 5896 4678 5908
rect 7742 5896 7748 5908
rect 4672 5868 7748 5896
rect 4672 5856 4678 5868
rect 7742 5856 7748 5868
rect 7800 5856 7806 5908
rect 8021 5899 8079 5905
rect 8021 5865 8033 5899
rect 8067 5896 8079 5899
rect 8202 5896 8208 5908
rect 8067 5868 8208 5896
rect 8067 5865 8079 5868
rect 8021 5859 8079 5865
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 11882 5896 11888 5908
rect 9232 5868 11888 5896
rect 3053 5831 3111 5837
rect 3053 5797 3065 5831
rect 3099 5828 3111 5831
rect 9232 5828 9260 5868
rect 11882 5856 11888 5868
rect 11940 5856 11946 5908
rect 11977 5899 12035 5905
rect 11977 5865 11989 5899
rect 12023 5896 12035 5899
rect 12250 5896 12256 5908
rect 12023 5868 12256 5896
rect 12023 5865 12035 5868
rect 11977 5859 12035 5865
rect 12250 5856 12256 5868
rect 12308 5856 12314 5908
rect 12342 5856 12348 5908
rect 12400 5896 12406 5908
rect 15286 5896 15292 5908
rect 12400 5868 15292 5896
rect 12400 5856 12406 5868
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 15473 5899 15531 5905
rect 15473 5865 15485 5899
rect 15519 5896 15531 5899
rect 15746 5896 15752 5908
rect 15519 5868 15752 5896
rect 15519 5865 15531 5868
rect 15473 5859 15531 5865
rect 15746 5856 15752 5868
rect 15804 5896 15810 5908
rect 16114 5896 16120 5908
rect 15804 5868 16120 5896
rect 15804 5856 15810 5868
rect 16114 5856 16120 5868
rect 16172 5856 16178 5908
rect 16574 5896 16580 5908
rect 16535 5868 16580 5896
rect 16574 5856 16580 5868
rect 16632 5856 16638 5908
rect 18046 5896 18052 5908
rect 17052 5868 18052 5896
rect 3099 5800 9260 5828
rect 3099 5797 3111 5800
rect 3053 5791 3111 5797
rect 10226 5788 10232 5840
rect 10284 5828 10290 5840
rect 10597 5831 10655 5837
rect 10597 5828 10609 5831
rect 10284 5800 10609 5828
rect 10284 5788 10290 5800
rect 10597 5797 10609 5800
rect 10643 5828 10655 5831
rect 11698 5828 11704 5840
rect 10643 5800 11704 5828
rect 10643 5797 10655 5800
rect 10597 5791 10655 5797
rect 11698 5788 11704 5800
rect 11756 5788 11762 5840
rect 12158 5788 12164 5840
rect 12216 5828 12222 5840
rect 12216 5800 12261 5828
rect 12216 5788 12222 5800
rect 12894 5788 12900 5840
rect 12952 5788 12958 5840
rect 13998 5788 14004 5840
rect 14056 5828 14062 5840
rect 15657 5831 15715 5837
rect 15657 5828 15669 5831
rect 14056 5800 15669 5828
rect 14056 5788 14062 5800
rect 15657 5797 15669 5800
rect 15703 5797 15715 5831
rect 15657 5791 15715 5797
rect 6178 5760 6184 5772
rect 2976 5732 6184 5760
rect 6178 5720 6184 5732
rect 6236 5720 6242 5772
rect 6270 5720 6276 5772
rect 6328 5760 6334 5772
rect 11514 5760 11520 5772
rect 6328 5732 9076 5760
rect 6328 5720 6334 5732
rect 1762 5692 1768 5704
rect 1723 5664 1768 5692
rect 1762 5652 1768 5664
rect 1820 5652 1826 5704
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5692 2191 5695
rect 2590 5692 2596 5704
rect 2179 5664 2596 5692
rect 2179 5661 2191 5664
rect 2133 5655 2191 5661
rect 2590 5652 2596 5664
rect 2648 5652 2654 5704
rect 4154 5692 4160 5704
rect 3237 5671 3295 5677
rect 3237 5637 3249 5671
rect 3283 5637 3295 5671
rect 4115 5664 4160 5692
rect 4154 5652 4160 5664
rect 4212 5652 4218 5704
rect 5721 5695 5779 5701
rect 5721 5661 5733 5695
rect 5767 5692 5779 5695
rect 6549 5695 6607 5701
rect 6549 5692 6561 5695
rect 5767 5664 6561 5692
rect 5767 5661 5779 5664
rect 5721 5655 5779 5661
rect 6549 5661 6561 5664
rect 6595 5661 6607 5695
rect 7837 5695 7895 5701
rect 7837 5692 7849 5695
rect 6549 5655 6607 5661
rect 7208 5664 7849 5692
rect 3237 5631 3295 5637
rect 2409 5559 2467 5565
rect 2409 5525 2421 5559
rect 2455 5556 2467 5559
rect 3050 5556 3056 5568
rect 2455 5528 3056 5556
rect 2455 5525 2467 5528
rect 2409 5519 2467 5525
rect 3050 5516 3056 5528
rect 3108 5516 3114 5568
rect 3252 5556 3280 5631
rect 4341 5627 4399 5633
rect 4341 5593 4353 5627
rect 4387 5624 4399 5627
rect 5074 5624 5080 5636
rect 4387 5596 5080 5624
rect 4387 5593 4399 5596
rect 4341 5587 4399 5593
rect 5074 5584 5080 5596
rect 5132 5584 5138 5636
rect 6086 5624 6092 5636
rect 5460 5596 6092 5624
rect 5460 5556 5488 5596
rect 6086 5584 6092 5596
rect 6144 5584 6150 5636
rect 6181 5627 6239 5633
rect 6181 5593 6193 5627
rect 6227 5593 6239 5627
rect 6181 5587 6239 5593
rect 6365 5627 6423 5633
rect 6365 5593 6377 5627
rect 6411 5624 6423 5627
rect 6454 5624 6460 5636
rect 6411 5596 6460 5624
rect 6411 5593 6423 5596
rect 6365 5587 6423 5593
rect 3252 5528 5488 5556
rect 5537 5559 5595 5565
rect 5537 5525 5549 5559
rect 5583 5556 5595 5559
rect 5902 5556 5908 5568
rect 5583 5528 5908 5556
rect 5583 5525 5595 5528
rect 5537 5519 5595 5525
rect 5902 5516 5908 5528
rect 5960 5516 5966 5568
rect 6196 5556 6224 5587
rect 6454 5584 6460 5596
rect 6512 5584 6518 5636
rect 7208 5633 7236 5664
rect 7837 5661 7849 5664
rect 7883 5692 7895 5695
rect 8938 5692 8944 5704
rect 7883 5664 8944 5692
rect 7883 5661 7895 5664
rect 7837 5655 7895 5661
rect 8938 5652 8944 5664
rect 8996 5652 9002 5704
rect 7193 5627 7251 5633
rect 7193 5593 7205 5627
rect 7239 5593 7251 5627
rect 7193 5587 7251 5593
rect 7006 5556 7012 5568
rect 6196 5528 7012 5556
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 7282 5556 7288 5568
rect 7243 5528 7288 5556
rect 7282 5516 7288 5528
rect 7340 5516 7346 5568
rect 9048 5556 9076 5732
rect 11072 5732 11520 5760
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5692 9275 5695
rect 9766 5692 9772 5704
rect 9263 5664 9772 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 9766 5652 9772 5664
rect 9824 5652 9830 5704
rect 9950 5652 9956 5704
rect 10008 5692 10014 5704
rect 11072 5692 11100 5732
rect 11514 5720 11520 5732
rect 11572 5720 11578 5772
rect 11790 5760 11796 5772
rect 11751 5732 11796 5760
rect 11790 5720 11796 5732
rect 11848 5720 11854 5772
rect 12802 5760 12808 5772
rect 11992 5732 12808 5760
rect 11238 5692 11244 5704
rect 10008 5664 11100 5692
rect 11199 5664 11244 5692
rect 10008 5652 10014 5664
rect 11238 5652 11244 5664
rect 11296 5652 11302 5704
rect 11330 5652 11336 5704
rect 11388 5692 11394 5704
rect 11992 5701 12020 5732
rect 12802 5720 12808 5732
rect 12860 5720 12866 5772
rect 12912 5701 12940 5788
rect 15102 5760 15108 5772
rect 13648 5732 15108 5760
rect 13648 5704 13676 5732
rect 15102 5720 15108 5732
rect 15160 5720 15166 5772
rect 15286 5760 15292 5772
rect 15247 5732 15292 5760
rect 15286 5720 15292 5732
rect 15344 5720 15350 5772
rect 16666 5760 16672 5772
rect 15396 5732 16672 5760
rect 11701 5695 11759 5701
rect 11701 5692 11713 5695
rect 11388 5664 11713 5692
rect 11388 5652 11394 5664
rect 11701 5661 11713 5664
rect 11747 5661 11759 5695
rect 11701 5655 11759 5661
rect 11977 5695 12035 5701
rect 11977 5661 11989 5695
rect 12023 5661 12035 5695
rect 11977 5655 12035 5661
rect 12897 5695 12955 5701
rect 12897 5661 12909 5695
rect 12943 5661 12955 5695
rect 12897 5655 12955 5661
rect 13541 5695 13599 5701
rect 13541 5661 13553 5695
rect 13587 5692 13599 5695
rect 13630 5692 13636 5704
rect 13587 5664 13636 5692
rect 13587 5661 13599 5664
rect 13541 5655 13599 5661
rect 13630 5652 13636 5664
rect 13688 5652 13694 5704
rect 14277 5695 14335 5701
rect 14277 5661 14289 5695
rect 14323 5692 14335 5695
rect 14461 5695 14519 5701
rect 14323 5664 14403 5692
rect 14323 5661 14335 5664
rect 14277 5655 14335 5661
rect 9484 5627 9542 5633
rect 9484 5593 9496 5627
rect 9530 5624 9542 5627
rect 9530 5596 11100 5624
rect 9530 5593 9542 5596
rect 9484 5587 9542 5593
rect 10870 5556 10876 5568
rect 9048 5528 10876 5556
rect 10870 5516 10876 5528
rect 10928 5516 10934 5568
rect 11072 5565 11100 5596
rect 13998 5584 14004 5636
rect 14056 5624 14062 5636
rect 14093 5627 14151 5633
rect 14093 5624 14105 5627
rect 14056 5596 14105 5624
rect 14056 5584 14062 5596
rect 14093 5593 14105 5596
rect 14139 5593 14151 5627
rect 14093 5587 14151 5593
rect 11057 5559 11115 5565
rect 11057 5525 11069 5559
rect 11103 5525 11115 5559
rect 11057 5519 11115 5525
rect 12713 5559 12771 5565
rect 12713 5525 12725 5559
rect 12759 5556 12771 5559
rect 12894 5556 12900 5568
rect 12759 5528 12900 5556
rect 12759 5525 12771 5528
rect 12713 5519 12771 5525
rect 12894 5516 12900 5528
rect 12952 5556 12958 5568
rect 13262 5556 13268 5568
rect 12952 5528 13268 5556
rect 12952 5516 12958 5528
rect 13262 5516 13268 5528
rect 13320 5516 13326 5568
rect 13357 5559 13415 5565
rect 13357 5525 13369 5559
rect 13403 5556 13415 5559
rect 13722 5556 13728 5568
rect 13403 5528 13728 5556
rect 13403 5525 13415 5528
rect 13357 5519 13415 5525
rect 13722 5516 13728 5528
rect 13780 5556 13786 5568
rect 14375 5556 14403 5664
rect 14461 5661 14473 5695
rect 14507 5692 14519 5695
rect 15396 5692 15424 5732
rect 16666 5720 16672 5732
rect 16724 5720 16730 5772
rect 17052 5760 17080 5868
rect 18046 5856 18052 5868
rect 18104 5856 18110 5908
rect 18414 5856 18420 5908
rect 18472 5896 18478 5908
rect 19150 5896 19156 5908
rect 18472 5868 19156 5896
rect 18472 5856 18478 5868
rect 19150 5856 19156 5868
rect 19208 5856 19214 5908
rect 19337 5899 19395 5905
rect 19337 5865 19349 5899
rect 19383 5896 19395 5899
rect 19426 5896 19432 5908
rect 19383 5868 19432 5896
rect 19383 5865 19395 5868
rect 19337 5859 19395 5865
rect 19426 5856 19432 5868
rect 19484 5856 19490 5908
rect 19610 5896 19616 5908
rect 19536 5868 19616 5896
rect 17126 5788 17132 5840
rect 17184 5828 17190 5840
rect 17865 5831 17923 5837
rect 17184 5800 17347 5828
rect 17184 5788 17190 5800
rect 17052 5732 17265 5760
rect 14507 5664 14872 5692
rect 14507 5661 14519 5664
rect 14461 5655 14519 5661
rect 14844 5624 14872 5664
rect 15089 5664 15424 5692
rect 15473 5695 15531 5701
rect 15089 5624 15117 5664
rect 15473 5661 15485 5695
rect 15519 5692 15531 5695
rect 16482 5692 16488 5704
rect 15519 5664 16488 5692
rect 15519 5661 15531 5664
rect 15473 5655 15531 5661
rect 16482 5652 16488 5664
rect 16540 5652 16546 5704
rect 17237 5701 17265 5732
rect 17130 5695 17188 5701
rect 17130 5661 17142 5695
rect 17176 5661 17188 5695
rect 17130 5655 17188 5661
rect 17222 5695 17280 5701
rect 17222 5661 17234 5695
rect 17268 5661 17280 5695
rect 17319 5692 17347 5800
rect 17865 5797 17877 5831
rect 17911 5828 17923 5831
rect 17911 5800 18736 5828
rect 17911 5797 17923 5800
rect 17865 5791 17923 5797
rect 17405 5763 17463 5769
rect 17405 5729 17417 5763
rect 17451 5760 17463 5763
rect 18598 5760 18604 5772
rect 17451 5732 18604 5760
rect 17451 5729 17463 5732
rect 17405 5723 17463 5729
rect 18598 5720 18604 5732
rect 18656 5720 18662 5772
rect 18708 5760 18736 5800
rect 19536 5760 19564 5868
rect 19610 5856 19616 5868
rect 19668 5856 19674 5908
rect 20898 5856 20904 5908
rect 20956 5896 20962 5908
rect 20993 5899 21051 5905
rect 20993 5896 21005 5899
rect 20956 5868 21005 5896
rect 20956 5856 20962 5868
rect 20993 5865 21005 5868
rect 21039 5865 21051 5899
rect 23842 5896 23848 5908
rect 23803 5868 23848 5896
rect 20993 5859 21051 5865
rect 23842 5856 23848 5868
rect 23900 5856 23906 5908
rect 26602 5896 26608 5908
rect 26563 5868 26608 5896
rect 26602 5856 26608 5868
rect 26660 5856 26666 5908
rect 26878 5856 26884 5908
rect 26936 5896 26942 5908
rect 30742 5896 30748 5908
rect 26936 5868 30748 5896
rect 26936 5856 26942 5868
rect 30742 5856 30748 5868
rect 30800 5856 30806 5908
rect 33410 5896 33416 5908
rect 33371 5868 33416 5896
rect 33410 5856 33416 5868
rect 33468 5856 33474 5908
rect 33594 5896 33600 5908
rect 33555 5868 33600 5896
rect 33594 5856 33600 5868
rect 33652 5856 33658 5908
rect 34606 5856 34612 5908
rect 34664 5896 34670 5908
rect 34885 5899 34943 5905
rect 34885 5896 34897 5899
rect 34664 5868 34897 5896
rect 34664 5856 34670 5868
rect 34885 5865 34897 5868
rect 34931 5865 34943 5899
rect 34885 5859 34943 5865
rect 35069 5899 35127 5905
rect 35069 5865 35081 5899
rect 35115 5896 35127 5899
rect 35802 5896 35808 5908
rect 35115 5868 35808 5896
rect 35115 5865 35127 5868
rect 35069 5859 35127 5865
rect 35802 5856 35808 5868
rect 35860 5856 35866 5908
rect 21266 5828 21272 5840
rect 18708 5732 19564 5760
rect 19720 5800 21272 5828
rect 17497 5695 17555 5701
rect 17497 5692 17509 5695
rect 17319 5664 17509 5692
rect 17222 5655 17280 5661
rect 17497 5661 17509 5664
rect 17543 5661 17555 5695
rect 17497 5655 17555 5661
rect 15194 5624 15200 5636
rect 14844 5596 15117 5624
rect 15155 5596 15200 5624
rect 15194 5584 15200 5596
rect 15252 5584 15258 5636
rect 16298 5624 16304 5636
rect 16211 5596 16304 5624
rect 16298 5584 16304 5596
rect 16356 5584 16362 5636
rect 17144 5624 17172 5655
rect 17678 5652 17684 5704
rect 17736 5692 17742 5704
rect 18325 5695 18383 5701
rect 18325 5692 18337 5695
rect 17736 5664 18337 5692
rect 17736 5652 17742 5664
rect 18325 5661 18337 5664
rect 18371 5661 18383 5695
rect 18325 5655 18383 5661
rect 17696 5624 17724 5652
rect 17144 5596 17724 5624
rect 18340 5624 18368 5655
rect 18414 5652 18420 5704
rect 18472 5692 18478 5704
rect 18708 5701 18736 5732
rect 18693 5695 18751 5701
rect 18472 5664 18517 5692
rect 18472 5652 18478 5664
rect 18693 5661 18705 5695
rect 18739 5661 18751 5695
rect 18693 5655 18751 5661
rect 19521 5695 19579 5701
rect 19521 5661 19533 5695
rect 19567 5661 19579 5695
rect 19521 5655 19579 5661
rect 19613 5695 19671 5701
rect 19613 5661 19625 5695
rect 19659 5688 19671 5695
rect 19720 5688 19748 5800
rect 21266 5788 21272 5800
rect 21324 5788 21330 5840
rect 21450 5788 21456 5840
rect 21508 5828 21514 5840
rect 22557 5831 22615 5837
rect 22557 5828 22569 5831
rect 21508 5800 22569 5828
rect 21508 5788 21514 5800
rect 22557 5797 22569 5800
rect 22603 5828 22615 5831
rect 24946 5828 24952 5840
rect 22603 5800 24952 5828
rect 22603 5797 22615 5800
rect 22557 5791 22615 5797
rect 24946 5788 24952 5800
rect 25004 5788 25010 5840
rect 28994 5788 29000 5840
rect 29052 5828 29058 5840
rect 29270 5828 29276 5840
rect 29052 5800 29276 5828
rect 29052 5788 29058 5800
rect 29270 5788 29276 5800
rect 29328 5788 29334 5840
rect 34422 5788 34428 5840
rect 34480 5828 34486 5840
rect 35986 5828 35992 5840
rect 34480 5800 35992 5828
rect 34480 5788 34486 5800
rect 35986 5788 35992 5800
rect 36044 5788 36050 5840
rect 36265 5831 36323 5837
rect 36265 5797 36277 5831
rect 36311 5828 36323 5831
rect 37366 5828 37372 5840
rect 36311 5800 37372 5828
rect 36311 5797 36323 5800
rect 36265 5791 36323 5797
rect 37366 5788 37372 5800
rect 37424 5788 37430 5840
rect 19797 5763 19855 5769
rect 19797 5729 19809 5763
rect 19843 5760 19855 5763
rect 19978 5760 19984 5772
rect 19843 5732 19984 5760
rect 19843 5729 19855 5732
rect 19797 5723 19855 5729
rect 19978 5720 19984 5732
rect 20036 5720 20042 5772
rect 27525 5763 27583 5769
rect 21192 5732 22324 5760
rect 19659 5661 19748 5688
rect 19613 5660 19748 5661
rect 19889 5695 19947 5701
rect 19889 5661 19901 5695
rect 19935 5692 19947 5695
rect 20438 5692 20444 5704
rect 19935 5664 20444 5692
rect 19935 5661 19947 5664
rect 19613 5655 19671 5660
rect 19889 5655 19947 5661
rect 19536 5624 19564 5655
rect 20438 5652 20444 5664
rect 20496 5652 20502 5704
rect 20533 5695 20591 5701
rect 20533 5661 20545 5695
rect 20579 5692 20591 5695
rect 20714 5692 20720 5704
rect 20579 5664 20720 5692
rect 20579 5661 20591 5664
rect 20533 5655 20591 5661
rect 20714 5652 20720 5664
rect 20772 5652 20778 5704
rect 21192 5701 21220 5732
rect 21177 5695 21235 5701
rect 21177 5661 21189 5695
rect 21223 5661 21235 5695
rect 21177 5655 21235 5661
rect 21269 5695 21327 5701
rect 21269 5661 21281 5695
rect 21315 5692 21327 5695
rect 21358 5692 21364 5704
rect 21315 5664 21364 5692
rect 21315 5661 21327 5664
rect 21269 5655 21327 5661
rect 21192 5624 21220 5655
rect 21358 5652 21364 5664
rect 21416 5652 21422 5704
rect 21545 5695 21603 5701
rect 21545 5661 21557 5695
rect 21591 5692 21603 5695
rect 21910 5692 21916 5704
rect 21591 5664 21916 5692
rect 21591 5661 21603 5664
rect 21545 5655 21603 5661
rect 21910 5652 21916 5664
rect 21968 5652 21974 5704
rect 22296 5701 22324 5732
rect 27525 5729 27537 5763
rect 27571 5760 27583 5763
rect 28258 5760 28264 5772
rect 27571 5732 28264 5760
rect 27571 5729 27583 5732
rect 27525 5723 27583 5729
rect 28258 5720 28264 5732
rect 28316 5720 28322 5772
rect 28350 5720 28356 5772
rect 28408 5760 28414 5772
rect 29546 5760 29552 5772
rect 28408 5732 29552 5760
rect 28408 5720 28414 5732
rect 29546 5720 29552 5732
rect 29604 5720 29610 5772
rect 31938 5760 31944 5772
rect 31899 5732 31944 5760
rect 31938 5720 31944 5732
rect 31996 5720 32002 5772
rect 32030 5720 32036 5772
rect 32088 5760 32094 5772
rect 32306 5760 32312 5772
rect 32088 5732 32312 5760
rect 32088 5720 32094 5732
rect 32306 5720 32312 5732
rect 32364 5720 32370 5772
rect 34054 5720 34060 5772
rect 34112 5760 34118 5772
rect 35802 5760 35808 5772
rect 34112 5732 35808 5760
rect 34112 5720 34118 5732
rect 35802 5720 35808 5732
rect 35860 5720 35866 5772
rect 22281 5695 22339 5701
rect 22281 5661 22293 5695
rect 22327 5661 22339 5695
rect 22281 5655 22339 5661
rect 22373 5695 22431 5701
rect 22373 5661 22385 5695
rect 22419 5661 22431 5695
rect 22373 5655 22431 5661
rect 22094 5624 22100 5636
rect 18340 5596 21220 5624
rect 22055 5596 22100 5624
rect 22094 5584 22100 5596
rect 22152 5584 22158 5636
rect 22388 5624 22416 5655
rect 22646 5652 22652 5704
rect 22704 5692 22710 5704
rect 23477 5695 23535 5701
rect 22704 5664 22749 5692
rect 22704 5652 22710 5664
rect 23477 5661 23489 5695
rect 23523 5692 23535 5695
rect 24118 5692 24124 5704
rect 23523 5664 24124 5692
rect 23523 5661 23535 5664
rect 23477 5655 23535 5661
rect 24118 5652 24124 5664
rect 24176 5652 24182 5704
rect 24394 5692 24400 5704
rect 24355 5664 24400 5692
rect 24394 5652 24400 5664
rect 24452 5652 24458 5704
rect 25225 5695 25283 5701
rect 25225 5661 25237 5695
rect 25271 5692 25283 5695
rect 26234 5692 26240 5704
rect 25271 5664 26240 5692
rect 25271 5661 25283 5664
rect 25225 5655 25283 5661
rect 26234 5652 26240 5664
rect 26292 5652 26298 5704
rect 27706 5652 27712 5704
rect 27764 5692 27770 5704
rect 27801 5695 27859 5701
rect 27801 5692 27813 5695
rect 27764 5664 27813 5692
rect 27764 5652 27770 5664
rect 27801 5661 27813 5664
rect 27847 5661 27859 5695
rect 28997 5695 29055 5701
rect 28997 5692 29009 5695
rect 27801 5655 27859 5661
rect 27908 5664 29009 5692
rect 23290 5624 23296 5636
rect 22388 5596 23296 5624
rect 23290 5584 23296 5596
rect 23348 5584 23354 5636
rect 23382 5584 23388 5636
rect 23440 5624 23446 5636
rect 23661 5627 23719 5633
rect 23661 5624 23673 5627
rect 23440 5596 23673 5624
rect 23440 5584 23446 5596
rect 23661 5593 23673 5596
rect 23707 5624 23719 5627
rect 24302 5624 24308 5636
rect 23707 5596 24308 5624
rect 23707 5593 23719 5596
rect 23661 5587 23719 5593
rect 24302 5584 24308 5596
rect 24360 5624 24366 5636
rect 24581 5627 24639 5633
rect 24581 5624 24593 5627
rect 24360 5596 24593 5624
rect 24360 5584 24366 5596
rect 24581 5593 24593 5596
rect 24627 5593 24639 5627
rect 24762 5624 24768 5636
rect 24723 5596 24768 5624
rect 24581 5587 24639 5593
rect 24762 5584 24768 5596
rect 24820 5584 24826 5636
rect 25492 5627 25550 5633
rect 25492 5593 25504 5627
rect 25538 5624 25550 5627
rect 26694 5624 26700 5636
rect 25538 5596 26700 5624
rect 25538 5593 25550 5596
rect 25492 5587 25550 5593
rect 26694 5584 26700 5596
rect 26752 5584 26758 5636
rect 13780 5528 14403 5556
rect 13780 5516 13786 5528
rect 15102 5516 15108 5568
rect 15160 5556 15166 5568
rect 16316 5556 16344 5584
rect 16942 5556 16948 5568
rect 15160 5528 16344 5556
rect 16903 5528 16948 5556
rect 15160 5516 15166 5528
rect 16942 5516 16948 5528
rect 17000 5516 17006 5568
rect 18138 5556 18144 5568
rect 18099 5528 18144 5556
rect 18138 5516 18144 5528
rect 18196 5516 18202 5568
rect 18598 5516 18604 5568
rect 18656 5556 18662 5568
rect 19978 5556 19984 5568
rect 18656 5528 19984 5556
rect 18656 5516 18662 5528
rect 19978 5516 19984 5528
rect 20036 5516 20042 5568
rect 20349 5559 20407 5565
rect 20349 5525 20361 5559
rect 20395 5556 20407 5559
rect 21818 5556 21824 5568
rect 20395 5528 21824 5556
rect 20395 5525 20407 5528
rect 20349 5519 20407 5525
rect 21818 5516 21824 5528
rect 21876 5516 21882 5568
rect 22370 5516 22376 5568
rect 22428 5556 22434 5568
rect 27908 5556 27936 5664
rect 28997 5661 29009 5664
rect 29043 5692 29055 5695
rect 29730 5692 29736 5704
rect 29043 5664 29736 5692
rect 29043 5661 29055 5664
rect 28997 5655 29055 5661
rect 29730 5652 29736 5664
rect 29788 5652 29794 5704
rect 30101 5695 30159 5701
rect 30101 5661 30113 5695
rect 30147 5692 30159 5695
rect 32217 5695 32275 5701
rect 30147 5664 31754 5692
rect 30147 5661 30159 5664
rect 30101 5655 30159 5661
rect 30374 5633 30380 5636
rect 30368 5587 30380 5633
rect 30432 5624 30438 5636
rect 31726 5624 31754 5664
rect 32217 5661 32229 5695
rect 32263 5661 32275 5695
rect 32217 5655 32275 5661
rect 32122 5624 32128 5636
rect 30432 5596 30468 5624
rect 31726 5596 32128 5624
rect 30374 5584 30380 5587
rect 30432 5584 30438 5596
rect 32122 5584 32128 5596
rect 32180 5584 32186 5636
rect 22428 5528 27936 5556
rect 28813 5559 28871 5565
rect 22428 5516 22434 5528
rect 28813 5525 28825 5559
rect 28859 5556 28871 5559
rect 28902 5556 28908 5568
rect 28859 5528 28908 5556
rect 28859 5525 28871 5528
rect 28813 5519 28871 5525
rect 28902 5516 28908 5528
rect 28960 5516 28966 5568
rect 30006 5516 30012 5568
rect 30064 5556 30070 5568
rect 30282 5556 30288 5568
rect 30064 5528 30288 5556
rect 30064 5516 30070 5528
rect 30282 5516 30288 5528
rect 30340 5516 30346 5568
rect 31481 5559 31539 5565
rect 31481 5525 31493 5559
rect 31527 5556 31539 5559
rect 31570 5556 31576 5568
rect 31527 5528 31576 5556
rect 31527 5525 31539 5528
rect 31481 5519 31539 5525
rect 31570 5516 31576 5528
rect 31628 5516 31634 5568
rect 32232 5556 32260 5655
rect 34146 5652 34152 5704
rect 34204 5692 34210 5704
rect 35713 5695 35771 5701
rect 35713 5692 35725 5695
rect 34204 5664 35725 5692
rect 34204 5652 34210 5664
rect 35713 5661 35725 5664
rect 35759 5661 35771 5695
rect 35713 5655 35771 5661
rect 36449 5695 36507 5701
rect 36449 5661 36461 5695
rect 36495 5692 36507 5695
rect 36906 5692 36912 5704
rect 36495 5664 36912 5692
rect 36495 5661 36507 5664
rect 36449 5655 36507 5661
rect 36906 5652 36912 5664
rect 36964 5652 36970 5704
rect 37090 5692 37096 5704
rect 37051 5664 37096 5692
rect 37090 5652 37096 5664
rect 37148 5652 37154 5704
rect 37734 5692 37740 5704
rect 37695 5664 37740 5692
rect 37734 5652 37740 5664
rect 37792 5652 37798 5704
rect 32398 5584 32404 5636
rect 32456 5624 32462 5636
rect 33042 5624 33048 5636
rect 32456 5596 33048 5624
rect 32456 5584 32462 5596
rect 33042 5584 33048 5596
rect 33100 5624 33106 5636
rect 33229 5627 33287 5633
rect 33229 5624 33241 5627
rect 33100 5596 33241 5624
rect 33100 5584 33106 5596
rect 33229 5593 33241 5596
rect 33275 5593 33287 5627
rect 33229 5587 33287 5593
rect 33445 5627 33503 5633
rect 33445 5593 33457 5627
rect 33491 5624 33503 5627
rect 34606 5624 34612 5636
rect 33491 5596 34612 5624
rect 33491 5593 33503 5596
rect 33445 5587 33503 5593
rect 32950 5556 32956 5568
rect 32232 5528 32956 5556
rect 32950 5516 32956 5528
rect 33008 5556 33014 5568
rect 33460 5556 33488 5587
rect 34606 5584 34612 5596
rect 34664 5584 34670 5636
rect 34701 5627 34759 5633
rect 34701 5593 34713 5627
rect 34747 5624 34759 5627
rect 35342 5624 35348 5636
rect 34747 5596 35348 5624
rect 34747 5593 34759 5596
rect 34701 5587 34759 5593
rect 35342 5584 35348 5596
rect 35400 5584 35406 5636
rect 33008 5528 33488 5556
rect 33008 5516 33014 5528
rect 34514 5516 34520 5568
rect 34572 5556 34578 5568
rect 34790 5556 34796 5568
rect 34572 5528 34796 5556
rect 34572 5516 34578 5528
rect 34790 5516 34796 5528
rect 34848 5556 34854 5568
rect 34901 5559 34959 5565
rect 34901 5556 34913 5559
rect 34848 5528 34913 5556
rect 34848 5516 34854 5528
rect 34901 5525 34913 5528
rect 34947 5525 34959 5559
rect 35526 5556 35532 5568
rect 35487 5528 35532 5556
rect 34901 5519 34959 5525
rect 35526 5516 35532 5528
rect 35584 5516 35590 5568
rect 36909 5559 36967 5565
rect 36909 5525 36921 5559
rect 36955 5556 36967 5559
rect 37458 5556 37464 5568
rect 36955 5528 37464 5556
rect 36955 5525 36967 5528
rect 36909 5519 36967 5525
rect 37458 5516 37464 5528
rect 37516 5516 37522 5568
rect 37553 5559 37611 5565
rect 37553 5525 37565 5559
rect 37599 5556 37611 5559
rect 37826 5556 37832 5568
rect 37599 5528 37832 5556
rect 37599 5525 37611 5528
rect 37553 5519 37611 5525
rect 37826 5516 37832 5528
rect 37884 5516 37890 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 4614 5352 4620 5364
rect 3108 5324 4620 5352
rect 3108 5312 3114 5324
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 4985 5355 5043 5361
rect 4985 5321 4997 5355
rect 5031 5352 5043 5355
rect 5074 5352 5080 5364
rect 5031 5324 5080 5352
rect 5031 5321 5043 5324
rect 4985 5315 5043 5321
rect 5074 5312 5080 5324
rect 5132 5352 5138 5364
rect 5350 5352 5356 5364
rect 5132 5324 5356 5352
rect 5132 5312 5138 5324
rect 5350 5312 5356 5324
rect 5408 5312 5414 5364
rect 5445 5355 5503 5361
rect 5445 5321 5457 5355
rect 5491 5321 5503 5355
rect 5445 5315 5503 5321
rect 2225 5287 2283 5293
rect 2225 5284 2237 5287
rect 1872 5256 2237 5284
rect 1872 5225 1900 5256
rect 2225 5253 2237 5256
rect 2271 5284 2283 5287
rect 2866 5284 2872 5296
rect 2271 5256 2872 5284
rect 2271 5253 2283 5256
rect 2225 5247 2283 5253
rect 2866 5244 2872 5256
rect 2924 5244 2930 5296
rect 3872 5287 3930 5293
rect 3872 5253 3884 5287
rect 3918 5284 3930 5287
rect 5460 5284 5488 5315
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 6914 5352 6920 5364
rect 5684 5324 6920 5352
rect 5684 5312 5690 5324
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 7837 5355 7895 5361
rect 7837 5321 7849 5355
rect 7883 5352 7895 5355
rect 7926 5352 7932 5364
rect 7883 5324 7932 5352
rect 7883 5321 7895 5324
rect 7837 5315 7895 5321
rect 7926 5312 7932 5324
rect 7984 5312 7990 5364
rect 8018 5312 8024 5364
rect 8076 5352 8082 5364
rect 9766 5352 9772 5364
rect 8076 5324 9772 5352
rect 8076 5312 8082 5324
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 9861 5355 9919 5361
rect 9861 5321 9873 5355
rect 9907 5352 9919 5355
rect 10318 5352 10324 5364
rect 9907 5324 10324 5352
rect 9907 5321 9919 5324
rect 9861 5315 9919 5321
rect 10318 5312 10324 5324
rect 10376 5312 10382 5364
rect 10873 5355 10931 5361
rect 10612 5324 10824 5352
rect 6365 5287 6423 5293
rect 3918 5256 5488 5284
rect 5543 5256 5764 5284
rect 3918 5253 3930 5256
rect 3872 5247 3930 5253
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5185 1915 5219
rect 1857 5179 1915 5185
rect 2501 5219 2559 5225
rect 2501 5185 2513 5219
rect 2547 5216 2559 5219
rect 2774 5216 2780 5228
rect 2547 5188 2780 5216
rect 2547 5185 2559 5188
rect 2501 5179 2559 5185
rect 2774 5176 2780 5188
rect 2832 5176 2838 5228
rect 3145 5219 3203 5225
rect 3145 5185 3157 5219
rect 3191 5216 3203 5219
rect 3418 5216 3424 5228
rect 3191 5188 3424 5216
rect 3191 5185 3203 5188
rect 3145 5179 3203 5185
rect 3418 5176 3424 5188
rect 3476 5176 3482 5228
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5216 3663 5219
rect 3694 5216 3700 5228
rect 3651 5188 3700 5216
rect 3651 5185 3663 5188
rect 3605 5179 3663 5185
rect 3694 5176 3700 5188
rect 3752 5176 3758 5228
rect 4614 5176 4620 5228
rect 4672 5216 4678 5228
rect 5543 5216 5571 5256
rect 4672 5188 5571 5216
rect 5637 5219 5695 5225
rect 5637 5212 5649 5219
rect 5683 5212 5695 5219
rect 4672 5176 4678 5188
rect 5626 5160 5632 5212
rect 5684 5179 5695 5212
rect 5736 5216 5764 5256
rect 6365 5253 6377 5287
rect 6411 5284 6423 5287
rect 7098 5284 7104 5296
rect 6411 5256 7104 5284
rect 6411 5253 6423 5256
rect 6365 5247 6423 5253
rect 7098 5244 7104 5256
rect 7156 5244 7162 5296
rect 10042 5284 10048 5296
rect 7208 5256 10048 5284
rect 6454 5216 6460 5228
rect 5736 5188 6460 5216
rect 5684 5160 5690 5179
rect 6454 5176 6460 5188
rect 6512 5216 6518 5228
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 6512 5188 6561 5216
rect 6512 5176 6518 5188
rect 6549 5185 6561 5188
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 5810 5108 5816 5160
rect 5868 5148 5874 5160
rect 7208 5148 7236 5256
rect 10042 5244 10048 5256
rect 10100 5244 10106 5296
rect 10612 5293 10640 5324
rect 10597 5287 10655 5293
rect 10597 5253 10609 5287
rect 10643 5253 10655 5287
rect 10796 5284 10824 5324
rect 10873 5321 10885 5355
rect 10919 5352 10931 5355
rect 10962 5352 10968 5364
rect 10919 5324 10968 5352
rect 10919 5321 10931 5324
rect 10873 5315 10931 5321
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 11330 5312 11336 5364
rect 11388 5352 11394 5364
rect 12805 5355 12863 5361
rect 11388 5324 12434 5352
rect 11388 5312 11394 5324
rect 11054 5284 11060 5296
rect 10796 5256 11060 5284
rect 10597 5247 10655 5253
rect 11054 5244 11060 5256
rect 11112 5244 11118 5296
rect 12406 5284 12434 5324
rect 12805 5321 12817 5355
rect 12851 5352 12863 5355
rect 15102 5352 15108 5364
rect 12851 5324 15108 5352
rect 12851 5321 12863 5324
rect 12805 5315 12863 5321
rect 15102 5312 15108 5324
rect 15160 5312 15166 5364
rect 17405 5355 17463 5361
rect 17405 5321 17417 5355
rect 17451 5352 17463 5355
rect 17494 5352 17500 5364
rect 17451 5324 17500 5352
rect 17451 5321 17463 5324
rect 17405 5315 17463 5321
rect 17494 5312 17500 5324
rect 17552 5312 17558 5364
rect 18509 5355 18567 5361
rect 18509 5321 18521 5355
rect 18555 5352 18567 5355
rect 18966 5352 18972 5364
rect 18555 5324 18972 5352
rect 18555 5321 18567 5324
rect 18509 5315 18567 5321
rect 18966 5312 18972 5324
rect 19024 5312 19030 5364
rect 20346 5312 20352 5364
rect 20404 5352 20410 5364
rect 20717 5355 20775 5361
rect 20717 5352 20729 5355
rect 20404 5324 20729 5352
rect 20404 5312 20410 5324
rect 20717 5321 20729 5324
rect 20763 5321 20775 5355
rect 20717 5315 20775 5321
rect 24210 5312 24216 5364
rect 24268 5352 24274 5364
rect 24673 5355 24731 5361
rect 24673 5352 24685 5355
rect 24268 5324 24685 5352
rect 24268 5312 24274 5324
rect 24673 5321 24685 5324
rect 24719 5321 24731 5355
rect 24673 5315 24731 5321
rect 24854 5312 24860 5364
rect 24912 5352 24918 5364
rect 25133 5355 25191 5361
rect 25133 5352 25145 5355
rect 24912 5324 25145 5352
rect 24912 5312 24918 5324
rect 25133 5321 25145 5324
rect 25179 5321 25191 5355
rect 27890 5352 27896 5364
rect 25133 5315 25191 5321
rect 25332 5324 27896 5352
rect 15197 5287 15255 5293
rect 15197 5284 15209 5287
rect 12406 5256 15209 5284
rect 15197 5253 15209 5256
rect 15243 5253 15255 5287
rect 15197 5247 15255 5253
rect 16942 5244 16948 5296
rect 17000 5284 17006 5296
rect 17037 5287 17095 5293
rect 17037 5284 17049 5287
rect 17000 5256 17049 5284
rect 17000 5244 17006 5256
rect 17037 5253 17049 5256
rect 17083 5253 17095 5287
rect 17037 5247 17095 5253
rect 17221 5287 17279 5293
rect 17221 5253 17233 5287
rect 17267 5284 17279 5287
rect 18138 5284 18144 5296
rect 17267 5256 17448 5284
rect 18099 5256 18144 5284
rect 17267 5253 17279 5256
rect 17221 5247 17279 5253
rect 17420 5228 17448 5256
rect 18138 5244 18144 5256
rect 18196 5244 18202 5296
rect 19604 5287 19662 5293
rect 19604 5253 19616 5287
rect 19650 5284 19662 5287
rect 20254 5284 20260 5296
rect 19650 5256 20260 5284
rect 19650 5253 19662 5256
rect 19604 5247 19662 5253
rect 20254 5244 20260 5256
rect 20312 5244 20318 5296
rect 23566 5293 23572 5296
rect 23560 5284 23572 5293
rect 23527 5256 23572 5284
rect 23560 5247 23572 5256
rect 23566 5244 23572 5247
rect 23624 5244 23630 5296
rect 25332 5284 25360 5324
rect 27890 5312 27896 5324
rect 27948 5312 27954 5364
rect 29454 5352 29460 5364
rect 28828 5324 29460 5352
rect 26602 5284 26608 5296
rect 24596 5256 25360 5284
rect 25424 5256 26608 5284
rect 7374 5216 7380 5228
rect 7335 5188 7380 5216
rect 7374 5176 7380 5188
rect 7432 5176 7438 5228
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5216 7711 5219
rect 8018 5216 8024 5228
rect 7699 5188 8024 5216
rect 7699 5185 7711 5188
rect 7653 5179 7711 5185
rect 8018 5176 8024 5188
rect 8076 5176 8082 5228
rect 8849 5219 8907 5225
rect 8849 5185 8861 5219
rect 8895 5216 8907 5219
rect 9122 5216 9128 5228
rect 8895 5188 9128 5216
rect 8895 5185 8907 5188
rect 8849 5179 8907 5185
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 9582 5216 9588 5228
rect 9543 5188 9588 5216
rect 9582 5176 9588 5188
rect 9640 5176 9646 5228
rect 9677 5219 9735 5225
rect 9677 5185 9689 5219
rect 9723 5185 9735 5219
rect 9677 5179 9735 5185
rect 7466 5148 7472 5160
rect 5868 5120 7236 5148
rect 7427 5120 7472 5148
rect 5868 5108 5874 5120
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 9692 5148 9720 5179
rect 10226 5176 10232 5228
rect 10284 5214 10290 5228
rect 10321 5219 10379 5225
rect 10321 5214 10333 5219
rect 10284 5186 10333 5214
rect 10284 5176 10290 5186
rect 10321 5185 10333 5186
rect 10367 5185 10379 5219
rect 10502 5216 10508 5228
rect 10463 5188 10508 5216
rect 10321 5179 10379 5185
rect 10502 5176 10508 5188
rect 10560 5176 10566 5228
rect 10713 5219 10771 5225
rect 10713 5216 10725 5219
rect 10704 5185 10725 5216
rect 10759 5185 10771 5219
rect 10704 5179 10771 5185
rect 10704 5148 10732 5179
rect 10870 5176 10876 5228
rect 10928 5216 10934 5228
rect 11701 5219 11759 5225
rect 10928 5188 11652 5216
rect 10928 5176 10934 5188
rect 9692 5120 10272 5148
rect 10704 5120 10885 5148
rect 1673 5083 1731 5089
rect 1673 5049 1685 5083
rect 1719 5080 1731 5083
rect 3602 5080 3608 5092
rect 1719 5052 3608 5080
rect 1719 5049 1731 5052
rect 1673 5043 1731 5049
rect 3602 5040 3608 5052
rect 3660 5040 3666 5092
rect 9766 5080 9772 5092
rect 4908 5052 5580 5080
rect 2314 5012 2320 5024
rect 2275 4984 2320 5012
rect 2314 4972 2320 4984
rect 2372 4972 2378 5024
rect 2961 5015 3019 5021
rect 2961 4981 2973 5015
rect 3007 5012 3019 5015
rect 4908 5012 4936 5052
rect 3007 4984 4936 5012
rect 3007 4981 3019 4984
rect 2961 4975 3019 4981
rect 4982 4972 4988 5024
rect 5040 5012 5046 5024
rect 5258 5012 5264 5024
rect 5040 4984 5264 5012
rect 5040 4972 5046 4984
rect 5258 4972 5264 4984
rect 5316 4972 5322 5024
rect 5552 5012 5580 5052
rect 5920 5052 9772 5080
rect 5920 5012 5948 5052
rect 9766 5040 9772 5052
rect 9824 5040 9830 5092
rect 10244 5080 10272 5120
rect 10594 5080 10600 5092
rect 10244 5052 10600 5080
rect 10594 5040 10600 5052
rect 10652 5040 10658 5092
rect 5552 4984 5948 5012
rect 5994 4972 6000 5024
rect 6052 5012 6058 5024
rect 6733 5015 6791 5021
rect 6733 5012 6745 5015
rect 6052 4984 6745 5012
rect 6052 4972 6058 4984
rect 6733 4981 6745 4984
rect 6779 4981 6791 5015
rect 7650 5012 7656 5024
rect 7611 4984 7656 5012
rect 6733 4975 6791 4981
rect 7650 4972 7656 4984
rect 7708 4972 7714 5024
rect 8665 5015 8723 5021
rect 8665 4981 8677 5015
rect 8711 5012 8723 5015
rect 8938 5012 8944 5024
rect 8711 4984 8944 5012
rect 8711 4981 8723 4984
rect 8665 4975 8723 4981
rect 8938 4972 8944 4984
rect 8996 5012 9002 5024
rect 9214 5012 9220 5024
rect 8996 4984 9220 5012
rect 8996 4972 9002 4984
rect 9214 4972 9220 4984
rect 9272 5012 9278 5024
rect 9582 5012 9588 5024
rect 9272 4984 9588 5012
rect 9272 4972 9278 4984
rect 9582 4972 9588 4984
rect 9640 5012 9646 5024
rect 10686 5012 10692 5024
rect 9640 4984 10692 5012
rect 9640 4972 9646 4984
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 10857 5012 10885 5120
rect 10962 5108 10968 5160
rect 11020 5148 11026 5160
rect 11517 5151 11575 5157
rect 11517 5148 11529 5151
rect 11020 5120 11529 5148
rect 11020 5108 11026 5120
rect 11517 5117 11529 5120
rect 11563 5117 11575 5151
rect 11624 5148 11652 5188
rect 11701 5185 11713 5219
rect 11747 5216 11759 5219
rect 12158 5216 12164 5228
rect 11747 5188 12164 5216
rect 11747 5185 11759 5188
rect 11701 5179 11759 5185
rect 12158 5176 12164 5188
rect 12216 5176 12222 5228
rect 12989 5219 13047 5225
rect 12989 5185 13001 5219
rect 13035 5185 13047 5219
rect 12989 5179 13047 5185
rect 12802 5148 12808 5160
rect 11624 5120 12808 5148
rect 11517 5111 11575 5117
rect 12802 5108 12808 5120
rect 12860 5108 12866 5160
rect 13004 5080 13032 5179
rect 13262 5176 13268 5228
rect 13320 5216 13326 5228
rect 13449 5219 13507 5225
rect 13449 5216 13461 5219
rect 13320 5188 13461 5216
rect 13320 5176 13326 5188
rect 13449 5185 13461 5188
rect 13495 5185 13507 5219
rect 13449 5179 13507 5185
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5216 13691 5219
rect 14642 5216 14648 5228
rect 13679 5188 14648 5216
rect 13679 5185 13691 5188
rect 13633 5179 13691 5185
rect 13464 5148 13492 5179
rect 14642 5176 14648 5188
rect 14700 5176 14706 5228
rect 15013 5219 15071 5225
rect 15013 5185 15025 5219
rect 15059 5216 15071 5219
rect 15562 5216 15568 5228
rect 15059 5188 15568 5216
rect 15059 5185 15071 5188
rect 15013 5179 15071 5185
rect 15562 5176 15568 5188
rect 15620 5176 15626 5228
rect 15838 5216 15844 5228
rect 15799 5188 15844 5216
rect 15838 5176 15844 5188
rect 15896 5176 15902 5228
rect 17402 5176 17408 5228
rect 17460 5216 17466 5228
rect 18325 5219 18383 5225
rect 18325 5216 18337 5219
rect 17460 5188 18337 5216
rect 17460 5176 17466 5188
rect 18325 5185 18337 5188
rect 18371 5185 18383 5219
rect 19334 5216 19340 5228
rect 19295 5188 19340 5216
rect 18325 5179 18383 5185
rect 19334 5176 19340 5188
rect 19392 5176 19398 5228
rect 21818 5216 21824 5228
rect 21779 5188 21824 5216
rect 21818 5176 21824 5188
rect 21876 5176 21882 5228
rect 22557 5219 22615 5225
rect 22557 5185 22569 5219
rect 22603 5216 22615 5219
rect 24596 5216 24624 5256
rect 22603 5188 24624 5216
rect 22603 5185 22615 5188
rect 22557 5179 22615 5185
rect 24670 5176 24676 5228
rect 24728 5216 24734 5228
rect 25424 5225 25452 5256
rect 26602 5244 26608 5256
rect 26660 5244 26666 5296
rect 28828 5293 28856 5324
rect 29454 5312 29460 5324
rect 29512 5312 29518 5364
rect 30374 5352 30380 5364
rect 30335 5324 30380 5352
rect 30374 5312 30380 5324
rect 30432 5312 30438 5364
rect 32769 5355 32827 5361
rect 32769 5352 32781 5355
rect 30484 5324 32781 5352
rect 28813 5287 28871 5293
rect 27172 5256 27936 5284
rect 25317 5219 25375 5225
rect 25317 5216 25329 5219
rect 24728 5188 25329 5216
rect 24728 5176 24734 5188
rect 25317 5185 25329 5188
rect 25363 5185 25375 5219
rect 25317 5179 25375 5185
rect 25409 5219 25467 5225
rect 25409 5185 25421 5219
rect 25455 5185 25467 5219
rect 25409 5179 25467 5185
rect 25685 5219 25743 5225
rect 25685 5185 25697 5219
rect 25731 5185 25743 5219
rect 25685 5179 25743 5185
rect 14829 5151 14887 5157
rect 14829 5148 14841 5151
rect 13464 5120 14841 5148
rect 14829 5117 14841 5120
rect 14875 5148 14887 5151
rect 15657 5151 15715 5157
rect 15657 5148 15669 5151
rect 14875 5120 15669 5148
rect 14875 5117 14887 5120
rect 14829 5111 14887 5117
rect 15657 5117 15669 5120
rect 15703 5117 15715 5151
rect 15657 5111 15715 5117
rect 22278 5108 22284 5160
rect 22336 5148 22342 5160
rect 23293 5151 23351 5157
rect 23293 5148 23305 5151
rect 22336 5120 23305 5148
rect 22336 5108 22342 5120
rect 23293 5117 23305 5120
rect 23339 5117 23351 5151
rect 23293 5111 23351 5117
rect 24946 5108 24952 5160
rect 25004 5148 25010 5160
rect 25593 5151 25651 5157
rect 25593 5148 25605 5151
rect 25004 5120 25605 5148
rect 25004 5108 25010 5120
rect 25593 5117 25605 5120
rect 25639 5117 25651 5151
rect 25700 5148 25728 5179
rect 25774 5176 25780 5228
rect 25832 5216 25838 5228
rect 27172 5225 27200 5256
rect 26329 5219 26387 5225
rect 26329 5216 26341 5219
rect 25832 5188 26341 5216
rect 25832 5176 25838 5188
rect 26329 5185 26341 5188
rect 26375 5216 26387 5219
rect 27157 5219 27215 5225
rect 27157 5216 27169 5219
rect 26375 5188 27169 5216
rect 26375 5185 26387 5188
rect 26329 5179 26387 5185
rect 27157 5185 27169 5188
rect 27203 5185 27215 5219
rect 27157 5179 27215 5185
rect 27338 5176 27344 5228
rect 27396 5216 27402 5228
rect 27801 5219 27859 5225
rect 27801 5216 27813 5219
rect 27396 5188 27813 5216
rect 27396 5176 27402 5188
rect 27801 5185 27813 5188
rect 27847 5185 27859 5219
rect 27908 5216 27936 5256
rect 28813 5253 28825 5287
rect 28859 5253 28871 5287
rect 28813 5247 28871 5253
rect 28994 5244 29000 5296
rect 29052 5293 29058 5296
rect 29052 5287 29071 5293
rect 29059 5253 29071 5287
rect 30484 5284 30512 5324
rect 32769 5321 32781 5324
rect 32815 5352 32827 5355
rect 34514 5352 34520 5364
rect 32815 5324 34520 5352
rect 32815 5321 32827 5324
rect 32769 5315 32827 5321
rect 34514 5312 34520 5324
rect 34572 5312 34578 5364
rect 34793 5355 34851 5361
rect 34793 5321 34805 5355
rect 34839 5352 34851 5355
rect 37274 5352 37280 5364
rect 34839 5324 37280 5352
rect 34839 5321 34851 5324
rect 34793 5315 34851 5321
rect 37274 5312 37280 5324
rect 37332 5312 37338 5364
rect 29052 5247 29071 5253
rect 29104 5256 30512 5284
rect 30745 5287 30803 5293
rect 29052 5244 29058 5247
rect 29104 5216 29132 5256
rect 30745 5253 30757 5287
rect 30791 5284 30803 5287
rect 31570 5284 31576 5296
rect 30791 5256 31576 5284
rect 30791 5253 30803 5256
rect 30745 5247 30803 5253
rect 31570 5244 31576 5256
rect 31628 5244 31634 5296
rect 32490 5284 32496 5296
rect 31726 5256 32496 5284
rect 27908 5188 29132 5216
rect 27801 5179 27859 5185
rect 29270 5176 29276 5228
rect 29328 5216 29334 5228
rect 29825 5219 29883 5225
rect 29825 5216 29837 5219
rect 29328 5188 29837 5216
rect 29328 5176 29334 5188
rect 29825 5185 29837 5188
rect 29871 5185 29883 5219
rect 30282 5216 30288 5228
rect 29825 5179 29883 5185
rect 29932 5188 30288 5216
rect 25866 5148 25872 5160
rect 25700 5120 25872 5148
rect 25593 5111 25651 5117
rect 25866 5108 25872 5120
rect 25924 5108 25930 5160
rect 27706 5108 27712 5160
rect 27764 5148 27770 5160
rect 28718 5148 28724 5160
rect 27764 5120 28724 5148
rect 27764 5108 27770 5120
rect 28718 5108 28724 5120
rect 28776 5148 28782 5160
rect 29932 5148 29960 5188
rect 30282 5176 30288 5188
rect 30340 5216 30346 5228
rect 30561 5219 30619 5225
rect 30561 5216 30573 5219
rect 30340 5188 30573 5216
rect 30340 5176 30346 5188
rect 30561 5185 30573 5188
rect 30607 5185 30619 5219
rect 30561 5179 30619 5185
rect 30837 5219 30895 5225
rect 30837 5185 30849 5219
rect 30883 5185 30895 5219
rect 30837 5179 30895 5185
rect 31481 5219 31539 5225
rect 31481 5185 31493 5219
rect 31527 5216 31539 5219
rect 31726 5216 31754 5256
rect 32490 5244 32496 5256
rect 32548 5244 32554 5296
rect 34425 5287 34483 5293
rect 34425 5253 34437 5287
rect 34471 5253 34483 5287
rect 34606 5284 34612 5296
rect 34664 5293 34670 5296
rect 34664 5287 34699 5293
rect 34551 5256 34612 5284
rect 34425 5247 34483 5253
rect 31527 5188 31754 5216
rect 32677 5219 32735 5225
rect 31527 5185 31539 5188
rect 31481 5179 31539 5185
rect 32677 5185 32689 5219
rect 32723 5216 32735 5219
rect 32766 5216 32772 5228
rect 32723 5188 32772 5216
rect 32723 5185 32735 5188
rect 32677 5179 32735 5185
rect 28776 5120 29960 5148
rect 28776 5108 28782 5120
rect 30190 5108 30196 5160
rect 30248 5148 30254 5160
rect 30852 5148 30880 5179
rect 32766 5176 32772 5188
rect 32824 5176 32830 5228
rect 33410 5176 33416 5228
rect 33468 5216 33474 5228
rect 33505 5219 33563 5225
rect 33505 5216 33517 5219
rect 33468 5188 33517 5216
rect 33468 5176 33474 5188
rect 33505 5185 33517 5188
rect 33551 5185 33563 5219
rect 34440 5216 34468 5247
rect 34606 5244 34612 5256
rect 34687 5284 34699 5287
rect 35894 5284 35900 5296
rect 34687 5256 35900 5284
rect 34687 5253 34699 5256
rect 34664 5247 34699 5253
rect 34664 5244 34670 5247
rect 35894 5244 35900 5256
rect 35952 5244 35958 5296
rect 34790 5216 34796 5228
rect 34440 5188 34796 5216
rect 33505 5179 33563 5185
rect 34790 5176 34796 5188
rect 34848 5176 34854 5228
rect 35342 5176 35348 5228
rect 35400 5216 35406 5228
rect 35437 5219 35495 5225
rect 35437 5216 35449 5219
rect 35400 5188 35449 5216
rect 35400 5176 35406 5188
rect 35437 5185 35449 5188
rect 35483 5185 35495 5219
rect 35437 5179 35495 5185
rect 36081 5219 36139 5225
rect 36081 5185 36093 5219
rect 36127 5185 36139 5219
rect 36081 5179 36139 5185
rect 30248 5120 30880 5148
rect 30248 5108 30254 5120
rect 34514 5108 34520 5160
rect 34572 5148 34578 5160
rect 36096 5148 36124 5179
rect 36262 5176 36268 5228
rect 36320 5216 36326 5228
rect 36725 5219 36783 5225
rect 36725 5216 36737 5219
rect 36320 5188 36737 5216
rect 36320 5176 36326 5188
rect 36725 5185 36737 5188
rect 36771 5185 36783 5219
rect 36725 5179 36783 5185
rect 37642 5176 37648 5228
rect 37700 5216 37706 5228
rect 37829 5219 37887 5225
rect 37829 5216 37841 5219
rect 37700 5188 37841 5216
rect 37700 5176 37706 5188
rect 37829 5185 37841 5188
rect 37875 5185 37887 5219
rect 37829 5179 37887 5185
rect 34572 5120 36124 5148
rect 34572 5108 34578 5120
rect 18598 5080 18604 5092
rect 13004 5052 18604 5080
rect 18598 5040 18604 5052
rect 18656 5040 18662 5092
rect 24394 5040 24400 5092
rect 24452 5080 24458 5092
rect 24452 5052 25728 5080
rect 24452 5040 24458 5052
rect 11330 5012 11336 5024
rect 10857 4984 11336 5012
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 11885 5015 11943 5021
rect 11885 4981 11897 5015
rect 11931 5012 11943 5015
rect 12434 5012 12440 5024
rect 11931 4984 12440 5012
rect 11931 4981 11943 4984
rect 11885 4975 11943 4981
rect 12434 4972 12440 4984
rect 12492 4972 12498 5024
rect 13817 5015 13875 5021
rect 13817 4981 13829 5015
rect 13863 5012 13875 5015
rect 13998 5012 14004 5024
rect 13863 4984 14004 5012
rect 13863 4981 13875 4984
rect 13817 4975 13875 4981
rect 13998 4972 14004 4984
rect 14056 4972 14062 5024
rect 14274 4972 14280 5024
rect 14332 5012 14338 5024
rect 15194 5012 15200 5024
rect 14332 4984 15200 5012
rect 14332 4972 14338 4984
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 15378 4972 15384 5024
rect 15436 5012 15442 5024
rect 16025 5015 16083 5021
rect 16025 5012 16037 5015
rect 15436 4984 16037 5012
rect 15436 4972 15442 4984
rect 16025 4981 16037 4984
rect 16071 4981 16083 5015
rect 16025 4975 16083 4981
rect 20898 4972 20904 5024
rect 20956 5012 20962 5024
rect 22005 5015 22063 5021
rect 22005 5012 22017 5015
rect 20956 4984 22017 5012
rect 20956 4972 20962 4984
rect 22005 4981 22017 4984
rect 22051 4981 22063 5015
rect 22005 4975 22063 4981
rect 22186 4972 22192 5024
rect 22244 5012 22250 5024
rect 22741 5015 22799 5021
rect 22741 5012 22753 5015
rect 22244 4984 22753 5012
rect 22244 4972 22250 4984
rect 22741 4981 22753 4984
rect 22787 4981 22799 5015
rect 22741 4975 22799 4981
rect 23934 4972 23940 5024
rect 23992 5012 23998 5024
rect 24210 5012 24216 5024
rect 23992 4984 24216 5012
rect 23992 4972 23998 4984
rect 24210 4972 24216 4984
rect 24268 4972 24274 5024
rect 25700 5012 25728 5052
rect 26050 5040 26056 5092
rect 26108 5080 26114 5092
rect 26973 5083 27031 5089
rect 26973 5080 26985 5083
rect 26108 5052 26985 5080
rect 26108 5040 26114 5052
rect 26973 5049 26985 5052
rect 27019 5049 27031 5083
rect 26973 5043 27031 5049
rect 29181 5083 29239 5089
rect 29181 5049 29193 5083
rect 29227 5080 29239 5083
rect 31018 5080 31024 5092
rect 29227 5052 31024 5080
rect 29227 5049 29239 5052
rect 29181 5043 29239 5049
rect 31018 5040 31024 5052
rect 31076 5040 31082 5092
rect 34698 5040 34704 5092
rect 34756 5080 34762 5092
rect 35253 5083 35311 5089
rect 35253 5080 35265 5083
rect 34756 5052 35265 5080
rect 34756 5040 34762 5052
rect 35253 5049 35265 5052
rect 35299 5049 35311 5083
rect 35253 5043 35311 5049
rect 26145 5015 26203 5021
rect 26145 5012 26157 5015
rect 25700 4984 26157 5012
rect 26145 4981 26157 4984
rect 26191 4981 26203 5015
rect 27614 5012 27620 5024
rect 27575 4984 27620 5012
rect 26145 4975 26203 4981
rect 27614 4972 27620 4984
rect 27672 4972 27678 5024
rect 28997 5015 29055 5021
rect 28997 4981 29009 5015
rect 29043 5012 29055 5015
rect 29086 5012 29092 5024
rect 29043 4984 29092 5012
rect 29043 4981 29055 4984
rect 28997 4975 29055 4981
rect 29086 4972 29092 4984
rect 29144 4972 29150 5024
rect 29546 4972 29552 5024
rect 29604 5012 29610 5024
rect 29641 5015 29699 5021
rect 29641 5012 29653 5015
rect 29604 4984 29653 5012
rect 29604 4972 29610 4984
rect 29641 4981 29653 4984
rect 29687 4981 29699 5015
rect 29641 4975 29699 4981
rect 29730 4972 29736 5024
rect 29788 5012 29794 5024
rect 31297 5015 31355 5021
rect 31297 5012 31309 5015
rect 29788 4984 31309 5012
rect 29788 4972 29794 4984
rect 31297 4981 31309 4984
rect 31343 4981 31355 5015
rect 31297 4975 31355 4981
rect 31386 4972 31392 5024
rect 31444 5012 31450 5024
rect 32214 5012 32220 5024
rect 31444 4984 32220 5012
rect 31444 4972 31450 4984
rect 32214 4972 32220 4984
rect 32272 4972 32278 5024
rect 33318 5012 33324 5024
rect 33279 4984 33324 5012
rect 33318 4972 33324 4984
rect 33376 4972 33382 5024
rect 34422 4972 34428 5024
rect 34480 5012 34486 5024
rect 34609 5015 34667 5021
rect 34609 5012 34621 5015
rect 34480 4984 34621 5012
rect 34480 4972 34486 4984
rect 34609 4981 34621 4984
rect 34655 4981 34667 5015
rect 35894 5012 35900 5024
rect 35855 4984 35900 5012
rect 34609 4975 34667 4981
rect 35894 4972 35900 4984
rect 35952 4972 35958 5024
rect 36541 5015 36599 5021
rect 36541 4981 36553 5015
rect 36587 5012 36599 5015
rect 37274 5012 37280 5024
rect 36587 4984 37280 5012
rect 36587 4981 36599 4984
rect 36541 4975 36599 4981
rect 37274 4972 37280 4984
rect 37332 4972 37338 5024
rect 38013 5015 38071 5021
rect 38013 4981 38025 5015
rect 38059 5012 38071 5015
rect 39758 5012 39764 5024
rect 38059 4984 39764 5012
rect 38059 4981 38071 4984
rect 38013 4975 38071 4981
rect 39758 4972 39764 4984
rect 39816 4972 39822 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 2314 4768 2320 4820
rect 2372 4808 2378 4820
rect 4341 4811 4399 4817
rect 2372 4780 4292 4808
rect 2372 4768 2378 4780
rect 2409 4743 2467 4749
rect 2409 4709 2421 4743
rect 2455 4740 2467 4743
rect 3050 4740 3056 4752
rect 2455 4712 2912 4740
rect 3011 4712 3056 4740
rect 2455 4709 2467 4712
rect 2409 4703 2467 4709
rect 2682 4672 2688 4684
rect 1964 4644 2688 4672
rect 1964 4613 1992 4644
rect 2682 4632 2688 4644
rect 2740 4632 2746 4684
rect 1949 4607 2007 4613
rect 1949 4573 1961 4607
rect 1995 4573 2007 4607
rect 1949 4567 2007 4573
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4573 2651 4607
rect 2884 4604 2912 4712
rect 3050 4700 3056 4712
rect 3108 4700 3114 4752
rect 4154 4740 4160 4752
rect 3160 4712 4160 4740
rect 3160 4604 3188 4712
rect 4154 4700 4160 4712
rect 4212 4700 4218 4752
rect 4264 4672 4292 4780
rect 4341 4777 4353 4811
rect 4387 4808 4399 4811
rect 5626 4808 5632 4820
rect 4387 4780 5632 4808
rect 4387 4777 4399 4780
rect 4341 4771 4399 4777
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 7006 4768 7012 4820
rect 7064 4808 7070 4820
rect 7653 4811 7711 4817
rect 7653 4808 7665 4811
rect 7064 4780 7665 4808
rect 7064 4768 7070 4780
rect 7653 4777 7665 4780
rect 7699 4777 7711 4811
rect 7653 4771 7711 4777
rect 7926 4768 7932 4820
rect 7984 4808 7990 4820
rect 8110 4808 8116 4820
rect 7984 4780 8116 4808
rect 7984 4768 7990 4780
rect 8110 4768 8116 4780
rect 8168 4768 8174 4820
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 9306 4808 9312 4820
rect 8260 4780 9312 4808
rect 8260 4768 8266 4780
rect 9306 4768 9312 4780
rect 9364 4768 9370 4820
rect 11790 4808 11796 4820
rect 11751 4780 11796 4808
rect 11790 4768 11796 4780
rect 11848 4768 11854 4820
rect 14642 4808 14648 4820
rect 14603 4780 14648 4808
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 18598 4808 18604 4820
rect 18559 4780 18604 4808
rect 18598 4768 18604 4780
rect 18656 4768 18662 4820
rect 21726 4768 21732 4820
rect 21784 4808 21790 4820
rect 22005 4811 22063 4817
rect 22005 4808 22017 4811
rect 21784 4780 22017 4808
rect 21784 4768 21790 4780
rect 22005 4777 22017 4780
rect 22051 4777 22063 4811
rect 22005 4771 22063 4777
rect 22094 4768 22100 4820
rect 22152 4808 22158 4820
rect 22462 4808 22468 4820
rect 22152 4780 22468 4808
rect 22152 4768 22158 4780
rect 22462 4768 22468 4780
rect 22520 4768 22526 4820
rect 22646 4768 22652 4820
rect 22704 4808 22710 4820
rect 28442 4808 28448 4820
rect 22704 4780 28448 4808
rect 22704 4768 22710 4780
rect 28442 4768 28448 4780
rect 28500 4768 28506 4820
rect 29730 4808 29736 4820
rect 29691 4780 29736 4808
rect 29730 4768 29736 4780
rect 29788 4768 29794 4820
rect 30558 4808 30564 4820
rect 29840 4780 30564 4808
rect 5261 4743 5319 4749
rect 5261 4709 5273 4743
rect 5307 4740 5319 4743
rect 5534 4740 5540 4752
rect 5307 4712 5540 4740
rect 5307 4709 5319 4712
rect 5261 4703 5319 4709
rect 5534 4700 5540 4712
rect 5592 4700 5598 4752
rect 7193 4743 7251 4749
rect 7193 4709 7205 4743
rect 7239 4709 7251 4743
rect 9490 4740 9496 4752
rect 7193 4703 7251 4709
rect 8036 4712 9496 4740
rect 7208 4672 7236 4703
rect 7650 4672 7656 4684
rect 4264 4644 5672 4672
rect 7208 4644 7656 4672
rect 2884 4576 3188 4604
rect 3237 4607 3295 4613
rect 2593 4567 2651 4573
rect 3237 4573 3249 4607
rect 3283 4604 3295 4607
rect 3878 4604 3884 4616
rect 3283 4576 3884 4604
rect 3283 4573 3295 4576
rect 3237 4567 3295 4573
rect 2608 4536 2636 4567
rect 3878 4564 3884 4576
rect 3936 4564 3942 4616
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4604 4031 4607
rect 4801 4607 4859 4613
rect 4801 4604 4813 4607
rect 4019 4576 4813 4604
rect 4019 4573 4031 4576
rect 3973 4567 4031 4573
rect 4801 4573 4813 4576
rect 4847 4573 4859 4607
rect 4982 4604 4988 4616
rect 4943 4576 4988 4604
rect 4801 4567 4859 4573
rect 4982 4564 4988 4576
rect 5040 4564 5046 4616
rect 5074 4564 5080 4616
rect 5132 4604 5138 4616
rect 5132 4576 5177 4604
rect 5132 4564 5138 4576
rect 5258 4564 5264 4616
rect 5316 4604 5322 4616
rect 5353 4607 5411 4613
rect 5353 4604 5365 4607
rect 5316 4576 5365 4604
rect 5316 4564 5322 4576
rect 5353 4573 5365 4576
rect 5399 4573 5411 4607
rect 5353 4567 5411 4573
rect 2866 4536 2872 4548
rect 2608 4508 2872 4536
rect 2866 4496 2872 4508
rect 2924 4496 2930 4548
rect 2976 4508 3280 4536
rect 1765 4471 1823 4477
rect 1765 4437 1777 4471
rect 1811 4468 1823 4471
rect 2976 4468 3004 4508
rect 1811 4440 3004 4468
rect 3252 4468 3280 4508
rect 4062 4496 4068 4548
rect 4120 4536 4126 4548
rect 4157 4539 4215 4545
rect 4157 4536 4169 4539
rect 4120 4508 4169 4536
rect 4120 4496 4126 4508
rect 4157 4505 4169 4508
rect 4203 4536 4215 4539
rect 4614 4536 4620 4548
rect 4203 4508 4620 4536
rect 4203 4505 4215 4508
rect 4157 4499 4215 4505
rect 4614 4496 4620 4508
rect 4672 4496 4678 4548
rect 5644 4536 5672 4644
rect 7650 4632 7656 4644
rect 7708 4672 7714 4684
rect 7708 4644 7972 4672
rect 7708 4632 7714 4644
rect 5810 4604 5816 4616
rect 5771 4576 5816 4604
rect 5810 4564 5816 4576
rect 5868 4564 5874 4616
rect 5902 4564 5908 4616
rect 5960 4604 5966 4616
rect 6069 4607 6127 4613
rect 6069 4604 6081 4607
rect 5960 4576 6081 4604
rect 5960 4564 5966 4576
rect 6069 4573 6081 4576
rect 6115 4573 6127 4607
rect 6069 4567 6127 4573
rect 6546 4564 6552 4616
rect 6604 4604 6610 4616
rect 7282 4604 7288 4616
rect 6604 4576 7288 4604
rect 6604 4564 6610 4576
rect 7282 4564 7288 4576
rect 7340 4604 7346 4616
rect 7944 4613 7972 4644
rect 7837 4607 7895 4613
rect 7837 4604 7849 4607
rect 7340 4576 7849 4604
rect 7340 4564 7346 4576
rect 7837 4573 7849 4576
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 7929 4607 7987 4613
rect 7929 4573 7941 4607
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 8036 4536 8064 4712
rect 9490 4700 9496 4712
rect 9548 4700 9554 4752
rect 9766 4700 9772 4752
rect 9824 4740 9830 4752
rect 20530 4740 20536 4752
rect 9824 4712 9869 4740
rect 19536 4712 20536 4740
rect 9824 4700 9830 4712
rect 8938 4672 8944 4684
rect 8899 4644 8944 4672
rect 8938 4632 8944 4644
rect 8996 4632 9002 4684
rect 9140 4644 10272 4672
rect 8202 4604 8208 4616
rect 8163 4576 8208 4604
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 9140 4613 9168 4644
rect 9125 4607 9183 4613
rect 9125 4573 9137 4607
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 9309 4607 9367 4613
rect 9309 4573 9321 4607
rect 9355 4604 9367 4607
rect 9953 4607 10011 4613
rect 9692 4604 9812 4606
rect 9953 4604 9965 4607
rect 9355 4578 9965 4604
rect 9355 4576 9720 4578
rect 9784 4576 9965 4578
rect 9355 4573 9367 4576
rect 9309 4567 9367 4573
rect 9953 4573 9965 4576
rect 9999 4573 10011 4607
rect 9953 4567 10011 4573
rect 5644 4508 8064 4536
rect 9398 4468 9404 4480
rect 3252 4440 9404 4468
rect 1811 4437 1823 4440
rect 1765 4431 1823 4437
rect 9398 4428 9404 4440
rect 9456 4428 9462 4480
rect 10244 4468 10272 4644
rect 10318 4632 10324 4684
rect 10376 4672 10382 4684
rect 10413 4675 10471 4681
rect 10413 4672 10425 4675
rect 10376 4644 10425 4672
rect 10376 4632 10382 4644
rect 10413 4641 10425 4644
rect 10459 4641 10471 4675
rect 10413 4635 10471 4641
rect 13906 4632 13912 4684
rect 13964 4672 13970 4684
rect 13964 4644 14412 4672
rect 13964 4632 13970 4644
rect 12434 4564 12440 4616
rect 12492 4604 12498 4616
rect 12492 4576 12537 4604
rect 12492 4564 12498 4576
rect 12618 4564 12624 4616
rect 12676 4604 12682 4616
rect 12894 4604 12900 4616
rect 12676 4576 12900 4604
rect 12676 4564 12682 4576
rect 12894 4564 12900 4576
rect 12952 4564 12958 4616
rect 13078 4604 13084 4616
rect 13039 4576 13084 4604
rect 13078 4564 13084 4576
rect 13136 4564 13142 4616
rect 14090 4604 14096 4616
rect 14051 4576 14096 4604
rect 14090 4564 14096 4576
rect 14148 4564 14154 4616
rect 14384 4613 14412 4644
rect 14734 4632 14740 4684
rect 14792 4672 14798 4684
rect 15105 4675 15163 4681
rect 15105 4672 15117 4675
rect 14792 4644 15117 4672
rect 14792 4632 14798 4644
rect 15105 4641 15117 4644
rect 15151 4641 15163 4675
rect 15105 4635 15163 4641
rect 17126 4632 17132 4684
rect 17184 4672 17190 4684
rect 17221 4675 17279 4681
rect 17221 4672 17233 4675
rect 17184 4644 17233 4672
rect 17184 4632 17190 4644
rect 17221 4641 17233 4644
rect 17267 4641 17279 4675
rect 17221 4635 17279 4641
rect 18233 4675 18291 4681
rect 18233 4641 18245 4675
rect 18279 4672 18291 4675
rect 19334 4672 19340 4684
rect 18279 4644 19340 4672
rect 18279 4641 18291 4644
rect 18233 4635 18291 4641
rect 19334 4632 19340 4644
rect 19392 4672 19398 4684
rect 19536 4681 19564 4712
rect 20530 4700 20536 4712
rect 20588 4700 20594 4752
rect 21818 4700 21824 4752
rect 21876 4740 21882 4752
rect 23385 4743 23443 4749
rect 23385 4740 23397 4743
rect 21876 4712 23397 4740
rect 21876 4700 21882 4712
rect 23385 4709 23397 4712
rect 23431 4709 23443 4743
rect 23385 4703 23443 4709
rect 23566 4700 23572 4752
rect 23624 4740 23630 4752
rect 25317 4743 25375 4749
rect 25317 4740 25329 4743
rect 23624 4712 25329 4740
rect 23624 4700 23630 4712
rect 25317 4709 25329 4712
rect 25363 4709 25375 4743
rect 25317 4703 25375 4709
rect 25866 4700 25872 4752
rect 25924 4740 25930 4752
rect 29840 4740 29868 4780
rect 30558 4768 30564 4780
rect 30616 4768 30622 4820
rect 31386 4808 31392 4820
rect 31347 4780 31392 4808
rect 31386 4768 31392 4780
rect 31444 4768 31450 4820
rect 31573 4811 31631 4817
rect 31573 4777 31585 4811
rect 31619 4808 31631 4811
rect 31754 4808 31760 4820
rect 31619 4780 31760 4808
rect 31619 4777 31631 4780
rect 31573 4771 31631 4777
rect 31754 4768 31760 4780
rect 31812 4768 31818 4820
rect 32214 4808 32220 4820
rect 32175 4780 32220 4808
rect 32214 4768 32220 4780
rect 32272 4768 32278 4820
rect 33042 4808 33048 4820
rect 33003 4780 33048 4808
rect 33042 4768 33048 4780
rect 33100 4768 33106 4820
rect 33134 4768 33140 4820
rect 33192 4808 33198 4820
rect 33229 4811 33287 4817
rect 33229 4808 33241 4811
rect 33192 4780 33241 4808
rect 33192 4768 33198 4780
rect 33229 4777 33241 4780
rect 33275 4777 33287 4811
rect 34885 4811 34943 4817
rect 34885 4808 34897 4811
rect 33229 4771 33287 4777
rect 34532 4780 34897 4808
rect 25924 4712 29868 4740
rect 29917 4743 29975 4749
rect 25924 4700 25930 4712
rect 29917 4709 29929 4743
rect 29963 4740 29975 4743
rect 32401 4743 32459 4749
rect 29963 4712 31754 4740
rect 29963 4709 29975 4712
rect 29917 4703 29975 4709
rect 19521 4675 19579 4681
rect 19521 4672 19533 4675
rect 19392 4644 19533 4672
rect 19392 4632 19398 4644
rect 19521 4641 19533 4644
rect 19567 4641 19579 4675
rect 19521 4635 19579 4641
rect 19889 4675 19947 4681
rect 19889 4641 19901 4675
rect 19935 4672 19947 4675
rect 23658 4672 23664 4684
rect 19935 4644 23664 4672
rect 19935 4641 19947 4644
rect 19889 4635 19947 4641
rect 23658 4632 23664 4644
rect 23716 4632 23722 4684
rect 27614 4672 27620 4684
rect 24412 4644 27620 4672
rect 14369 4607 14427 4613
rect 14369 4573 14381 4607
rect 14415 4573 14427 4607
rect 14369 4567 14427 4573
rect 14458 4564 14464 4616
rect 14516 4604 14522 4616
rect 14516 4576 14561 4604
rect 14516 4564 14522 4576
rect 14642 4564 14648 4616
rect 14700 4604 14706 4616
rect 16945 4607 17003 4613
rect 16945 4604 16957 4607
rect 14700 4576 16957 4604
rect 14700 4564 14706 4576
rect 16945 4573 16957 4576
rect 16991 4604 17003 4607
rect 17586 4604 17592 4616
rect 16991 4576 17592 4604
rect 16991 4573 17003 4576
rect 16945 4567 17003 4573
rect 17586 4564 17592 4576
rect 17644 4564 17650 4616
rect 18414 4604 18420 4616
rect 18375 4576 18420 4604
rect 18414 4564 18420 4576
rect 18472 4564 18478 4616
rect 19705 4607 19763 4613
rect 19705 4573 19717 4607
rect 19751 4604 19763 4607
rect 19978 4604 19984 4616
rect 19751 4576 19984 4604
rect 19751 4573 19763 4576
rect 19705 4567 19763 4573
rect 19978 4564 19984 4576
rect 20036 4564 20042 4616
rect 20349 4607 20407 4613
rect 20349 4573 20361 4607
rect 20395 4573 20407 4607
rect 20349 4567 20407 4573
rect 10680 4539 10738 4545
rect 10680 4505 10692 4539
rect 10726 4536 10738 4539
rect 14274 4536 14280 4548
rect 10726 4508 12296 4536
rect 14235 4508 14280 4536
rect 10726 4505 10738 4508
rect 10680 4499 10738 4505
rect 10594 4468 10600 4480
rect 10244 4440 10600 4468
rect 10594 4428 10600 4440
rect 10652 4428 10658 4480
rect 12268 4477 12296 4508
rect 14274 4496 14280 4508
rect 14332 4496 14338 4548
rect 15350 4539 15408 4545
rect 15350 4536 15362 4539
rect 14384 4508 15362 4536
rect 12253 4471 12311 4477
rect 12253 4437 12265 4471
rect 12299 4437 12311 4471
rect 13262 4468 13268 4480
rect 13223 4440 13268 4468
rect 12253 4431 12311 4437
rect 13262 4428 13268 4440
rect 13320 4428 13326 4480
rect 13630 4428 13636 4480
rect 13688 4468 13694 4480
rect 14384 4468 14412 4508
rect 15350 4505 15362 4508
rect 15396 4505 15408 4539
rect 15350 4499 15408 4505
rect 16574 4496 16580 4548
rect 16632 4536 16638 4548
rect 20364 4536 20392 4567
rect 20530 4564 20536 4616
rect 20588 4604 20594 4616
rect 21637 4607 21695 4613
rect 21637 4604 21649 4607
rect 20588 4576 21649 4604
rect 20588 4564 20594 4576
rect 21637 4573 21649 4576
rect 21683 4573 21695 4607
rect 21637 4567 21695 4573
rect 21821 4607 21879 4613
rect 21821 4573 21833 4607
rect 21867 4604 21879 4607
rect 22370 4604 22376 4616
rect 21867 4576 22376 4604
rect 21867 4573 21879 4576
rect 21821 4567 21879 4573
rect 22370 4564 22376 4576
rect 22428 4564 22434 4616
rect 22465 4607 22523 4613
rect 22465 4573 22477 4607
rect 22511 4573 22523 4607
rect 23198 4604 23204 4616
rect 23159 4576 23204 4604
rect 22465 4567 22523 4573
rect 16632 4508 20392 4536
rect 22480 4536 22508 4567
rect 23198 4564 23204 4576
rect 23256 4564 23262 4616
rect 24412 4613 24440 4644
rect 27614 4632 27620 4644
rect 27672 4632 27678 4684
rect 28089 4644 29040 4672
rect 24397 4607 24455 4613
rect 24397 4573 24409 4607
rect 24443 4573 24455 4607
rect 25130 4604 25136 4616
rect 25091 4576 25136 4604
rect 24397 4567 24455 4573
rect 25130 4564 25136 4576
rect 25188 4564 25194 4616
rect 26050 4564 26056 4616
rect 26108 4604 26114 4616
rect 26237 4607 26295 4613
rect 26237 4604 26249 4607
rect 26108 4576 26249 4604
rect 26108 4564 26114 4576
rect 26237 4573 26249 4576
rect 26283 4573 26295 4607
rect 26237 4567 26295 4573
rect 26421 4607 26479 4613
rect 26421 4573 26433 4607
rect 26467 4604 26479 4607
rect 26786 4604 26792 4616
rect 26467 4576 26792 4604
rect 26467 4573 26479 4576
rect 26421 4567 26479 4573
rect 26786 4564 26792 4576
rect 26844 4564 26850 4616
rect 27706 4564 27712 4616
rect 27764 4604 27770 4616
rect 28089 4613 28117 4644
rect 29012 4616 29040 4644
rect 27801 4607 27859 4613
rect 27801 4604 27813 4607
rect 27764 4576 27813 4604
rect 27764 4564 27770 4576
rect 27801 4573 27813 4576
rect 27847 4573 27859 4607
rect 27801 4567 27859 4573
rect 28077 4607 28135 4613
rect 28077 4573 28089 4607
rect 28123 4573 28135 4607
rect 28718 4604 28724 4616
rect 28679 4576 28724 4604
rect 28077 4567 28135 4573
rect 28718 4564 28724 4576
rect 28776 4564 28782 4616
rect 28994 4604 29000 4616
rect 28955 4576 29000 4604
rect 28994 4564 29000 4576
rect 29052 4564 29058 4616
rect 30561 4607 30619 4613
rect 30561 4604 30573 4607
rect 29104 4576 30573 4604
rect 24762 4536 24768 4548
rect 22480 4508 24768 4536
rect 16632 4496 16638 4508
rect 24762 4496 24768 4508
rect 24820 4496 24826 4548
rect 26605 4539 26663 4545
rect 26605 4505 26617 4539
rect 26651 4536 26663 4539
rect 29104 4536 29132 4576
rect 30561 4573 30573 4576
rect 30607 4573 30619 4607
rect 31726 4604 31754 4712
rect 32401 4709 32413 4743
rect 32447 4709 32459 4743
rect 33060 4740 33088 4768
rect 34422 4740 34428 4752
rect 33060 4712 34428 4740
rect 32401 4703 32459 4709
rect 32416 4672 32444 4703
rect 34422 4700 34428 4712
rect 34480 4740 34486 4752
rect 34532 4740 34560 4780
rect 34885 4777 34897 4780
rect 34931 4777 34943 4811
rect 34885 4771 34943 4777
rect 35069 4811 35127 4817
rect 35069 4777 35081 4811
rect 35115 4808 35127 4811
rect 35710 4808 35716 4820
rect 35115 4780 35716 4808
rect 35115 4777 35127 4780
rect 35069 4771 35127 4777
rect 35710 4768 35716 4780
rect 35768 4768 35774 4820
rect 34480 4712 34560 4740
rect 34480 4700 34486 4712
rect 34606 4700 34612 4752
rect 34664 4740 34670 4752
rect 35342 4740 35348 4752
rect 34664 4712 35348 4740
rect 34664 4700 34670 4712
rect 35342 4700 35348 4712
rect 35400 4700 35406 4752
rect 35802 4700 35808 4752
rect 35860 4740 35866 4752
rect 35860 4712 37044 4740
rect 35860 4700 35866 4712
rect 32416 4644 36400 4672
rect 33873 4607 33931 4613
rect 33873 4604 33885 4607
rect 31726 4576 33885 4604
rect 30561 4567 30619 4573
rect 33873 4573 33885 4576
rect 33919 4573 33931 4607
rect 33873 4567 33931 4573
rect 33962 4564 33968 4616
rect 34020 4604 34026 4616
rect 35710 4604 35716 4616
rect 34020 4576 35572 4604
rect 35671 4576 35716 4604
rect 34020 4564 34026 4576
rect 26651 4508 29132 4536
rect 26651 4505 26663 4508
rect 26605 4499 26663 4505
rect 29454 4496 29460 4548
rect 29512 4536 29518 4548
rect 29549 4539 29607 4545
rect 29549 4536 29561 4539
rect 29512 4508 29561 4536
rect 29512 4496 29518 4508
rect 29549 4505 29561 4508
rect 29595 4505 29607 4539
rect 31202 4536 31208 4548
rect 31163 4508 31208 4536
rect 29549 4499 29607 4505
rect 31202 4496 31208 4508
rect 31260 4496 31266 4548
rect 31421 4539 31479 4545
rect 31421 4505 31433 4539
rect 31467 4536 31479 4539
rect 31467 4508 31616 4536
rect 31467 4505 31479 4508
rect 31421 4499 31479 4505
rect 16482 4468 16488 4480
rect 13688 4440 14412 4468
rect 16443 4440 16488 4468
rect 13688 4428 13694 4440
rect 16482 4428 16488 4440
rect 16540 4428 16546 4480
rect 18138 4428 18144 4480
rect 18196 4468 18202 4480
rect 20533 4471 20591 4477
rect 20533 4468 20545 4471
rect 18196 4440 20545 4468
rect 18196 4428 18202 4440
rect 20533 4437 20545 4440
rect 20579 4437 20591 4471
rect 20533 4431 20591 4437
rect 20622 4428 20628 4480
rect 20680 4468 20686 4480
rect 22649 4471 22707 4477
rect 22649 4468 22661 4471
rect 20680 4440 22661 4468
rect 20680 4428 20686 4440
rect 22649 4437 22661 4440
rect 22695 4437 22707 4471
rect 22649 4431 22707 4437
rect 23474 4428 23480 4480
rect 23532 4468 23538 4480
rect 24581 4471 24639 4477
rect 24581 4468 24593 4471
rect 23532 4440 24593 4468
rect 23532 4428 23538 4440
rect 24581 4437 24593 4440
rect 24627 4437 24639 4471
rect 27614 4468 27620 4480
rect 27575 4440 27620 4468
rect 24581 4431 24639 4437
rect 27614 4428 27620 4440
rect 27672 4428 27678 4480
rect 27985 4471 28043 4477
rect 27985 4437 27997 4471
rect 28031 4468 28043 4471
rect 28350 4468 28356 4480
rect 28031 4440 28356 4468
rect 28031 4437 28043 4440
rect 27985 4431 28043 4437
rect 28350 4428 28356 4440
rect 28408 4428 28414 4480
rect 28442 4428 28448 4480
rect 28500 4468 28506 4480
rect 28537 4471 28595 4477
rect 28537 4468 28549 4471
rect 28500 4440 28549 4468
rect 28500 4428 28506 4440
rect 28537 4437 28549 4440
rect 28583 4437 28595 4471
rect 28537 4431 28595 4437
rect 28810 4428 28816 4480
rect 28868 4468 28874 4480
rect 28905 4471 28963 4477
rect 28905 4468 28917 4471
rect 28868 4440 28917 4468
rect 28868 4428 28874 4440
rect 28905 4437 28917 4440
rect 28951 4437 28963 4471
rect 28905 4431 28963 4437
rect 29086 4428 29092 4480
rect 29144 4468 29150 4480
rect 29749 4471 29807 4477
rect 29749 4468 29761 4471
rect 29144 4440 29761 4468
rect 29144 4428 29150 4440
rect 29749 4437 29761 4440
rect 29795 4437 29807 4471
rect 30374 4468 30380 4480
rect 30335 4440 30380 4468
rect 29749 4431 29807 4437
rect 30374 4428 30380 4440
rect 30432 4428 30438 4480
rect 31588 4468 31616 4508
rect 31662 4496 31668 4548
rect 31720 4536 31726 4548
rect 32033 4539 32091 4545
rect 32033 4536 32045 4539
rect 31720 4508 32045 4536
rect 31720 4496 31726 4508
rect 32033 4505 32045 4508
rect 32079 4505 32091 4539
rect 32033 4499 32091 4505
rect 32861 4539 32919 4545
rect 32861 4505 32873 4539
rect 32907 4536 32919 4539
rect 33502 4536 33508 4548
rect 32907 4508 33508 4536
rect 32907 4505 32919 4508
rect 32861 4499 32919 4505
rect 33502 4496 33508 4508
rect 33560 4496 33566 4548
rect 34330 4496 34336 4548
rect 34388 4536 34394 4548
rect 34701 4539 34759 4545
rect 34701 4536 34713 4539
rect 34388 4508 34713 4536
rect 34388 4496 34394 4508
rect 34701 4505 34713 4508
rect 34747 4505 34759 4539
rect 34701 4499 34759 4505
rect 32214 4468 32220 4480
rect 32272 4477 32278 4480
rect 32272 4471 32291 4477
rect 31588 4440 32220 4468
rect 32214 4428 32220 4440
rect 32279 4437 32291 4471
rect 32272 4431 32291 4437
rect 32272 4428 32278 4431
rect 32950 4428 32956 4480
rect 33008 4468 33014 4480
rect 33061 4471 33119 4477
rect 33061 4468 33073 4471
rect 33008 4440 33073 4468
rect 33008 4428 33014 4440
rect 33061 4437 33073 4440
rect 33107 4437 33119 4471
rect 33061 4431 33119 4437
rect 33226 4428 33232 4480
rect 33284 4468 33290 4480
rect 33689 4471 33747 4477
rect 33689 4468 33701 4471
rect 33284 4440 33701 4468
rect 33284 4428 33290 4440
rect 33689 4437 33701 4440
rect 33735 4437 33747 4471
rect 33689 4431 33747 4437
rect 34882 4428 34888 4480
rect 34940 4477 34946 4480
rect 35544 4477 35572 4576
rect 35710 4564 35716 4576
rect 35768 4564 35774 4616
rect 36372 4613 36400 4644
rect 37016 4613 37044 4712
rect 36357 4607 36415 4613
rect 36357 4573 36369 4607
rect 36403 4573 36415 4607
rect 36357 4567 36415 4573
rect 37001 4607 37059 4613
rect 37001 4573 37013 4607
rect 37047 4573 37059 4607
rect 37001 4567 37059 4573
rect 37550 4564 37556 4616
rect 37608 4604 37614 4616
rect 37829 4607 37887 4613
rect 37829 4604 37841 4607
rect 37608 4576 37841 4604
rect 37608 4564 37614 4576
rect 37829 4573 37841 4576
rect 37875 4573 37887 4607
rect 37829 4567 37887 4573
rect 34940 4471 34959 4477
rect 34947 4437 34959 4471
rect 34940 4431 34959 4437
rect 35529 4471 35587 4477
rect 35529 4437 35541 4471
rect 35575 4437 35587 4471
rect 36170 4468 36176 4480
rect 36131 4440 36176 4468
rect 35529 4431 35587 4437
rect 34940 4428 34946 4431
rect 36170 4428 36176 4440
rect 36228 4428 36234 4480
rect 36446 4428 36452 4480
rect 36504 4468 36510 4480
rect 36817 4471 36875 4477
rect 36817 4468 36829 4471
rect 36504 4440 36829 4468
rect 36504 4428 36510 4440
rect 36817 4437 36829 4440
rect 36863 4437 36875 4471
rect 36817 4431 36875 4437
rect 38013 4471 38071 4477
rect 38013 4437 38025 4471
rect 38059 4468 38071 4471
rect 39022 4468 39028 4480
rect 38059 4440 39028 4468
rect 38059 4437 38071 4440
rect 38013 4431 38071 4437
rect 39022 4428 39028 4440
rect 39080 4428 39086 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 1949 4267 2007 4273
rect 1949 4233 1961 4267
rect 1995 4264 2007 4267
rect 2038 4264 2044 4276
rect 1995 4236 2044 4264
rect 1995 4233 2007 4236
rect 1949 4227 2007 4233
rect 2038 4224 2044 4236
rect 2096 4224 2102 4276
rect 3234 4264 3240 4276
rect 2148 4236 2774 4264
rect 3195 4236 3240 4264
rect 2148 4137 2176 4236
rect 2746 4196 2774 4236
rect 3234 4224 3240 4236
rect 3292 4224 3298 4276
rect 3418 4224 3424 4276
rect 3476 4264 3482 4276
rect 12250 4264 12256 4276
rect 3476 4236 12256 4264
rect 3476 4224 3482 4236
rect 12250 4224 12256 4236
rect 12308 4224 12314 4276
rect 14090 4224 14096 4276
rect 14148 4264 14154 4276
rect 15013 4267 15071 4273
rect 15013 4264 15025 4267
rect 14148 4236 15025 4264
rect 14148 4224 14154 4236
rect 15013 4233 15025 4236
rect 15059 4233 15071 4267
rect 15013 4227 15071 4233
rect 15562 4224 15568 4276
rect 15620 4264 15626 4276
rect 16025 4267 16083 4273
rect 16025 4264 16037 4267
rect 15620 4236 16037 4264
rect 15620 4224 15626 4236
rect 16025 4233 16037 4236
rect 16071 4233 16083 4267
rect 16025 4227 16083 4233
rect 18322 4224 18328 4276
rect 18380 4264 18386 4276
rect 19797 4267 19855 4273
rect 18380 4236 19647 4264
rect 18380 4224 18386 4236
rect 3694 4196 3700 4208
rect 2746 4168 3700 4196
rect 3694 4156 3700 4168
rect 3752 4156 3758 4208
rect 3786 4156 3792 4208
rect 3844 4196 3850 4208
rect 5902 4196 5908 4208
rect 3844 4168 5908 4196
rect 3844 4156 3850 4168
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4097 2191 4131
rect 2133 4091 2191 4097
rect 2777 4131 2835 4137
rect 2777 4097 2789 4131
rect 2823 4128 2835 4131
rect 3234 4128 3240 4140
rect 2823 4100 3240 4128
rect 2823 4097 2835 4100
rect 2777 4091 2835 4097
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 3896 4137 3924 4168
rect 5902 4156 5908 4168
rect 5960 4196 5966 4208
rect 10318 4196 10324 4208
rect 5960 4168 10324 4196
rect 5960 4156 5966 4168
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4097 3479 4131
rect 3421 4091 3479 4097
rect 3881 4131 3939 4137
rect 3881 4097 3893 4131
rect 3927 4097 3939 4131
rect 3881 4091 3939 4097
rect 4148 4131 4206 4137
rect 4148 4097 4160 4131
rect 4194 4128 4206 4131
rect 4614 4128 4620 4140
rect 4194 4100 4620 4128
rect 4194 4097 4206 4100
rect 4148 4091 4206 4097
rect 3436 4060 3464 4091
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 4982 4088 4988 4140
rect 5040 4128 5046 4140
rect 6546 4128 6552 4140
rect 5040 4100 6552 4128
rect 5040 4088 5046 4100
rect 6546 4088 6552 4100
rect 6604 4088 6610 4140
rect 6638 4088 6644 4140
rect 6696 4128 6702 4140
rect 6914 4128 6920 4140
rect 6696 4100 6741 4128
rect 6875 4100 6920 4128
rect 6696 4088 6702 4100
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 7392 4137 7420 4168
rect 9232 4137 9260 4168
rect 10318 4156 10324 4168
rect 10376 4156 10382 4208
rect 11238 4156 11244 4208
rect 11296 4196 11302 4208
rect 12038 4199 12096 4205
rect 12038 4196 12050 4199
rect 11296 4168 12050 4196
rect 11296 4156 11302 4168
rect 12038 4165 12050 4168
rect 12084 4165 12096 4199
rect 14734 4196 14740 4208
rect 12038 4159 12096 4165
rect 13832 4168 14740 4196
rect 9490 4137 9496 4140
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 7644 4131 7702 4137
rect 7644 4097 7656 4131
rect 7690 4128 7702 4131
rect 9217 4131 9275 4137
rect 7690 4100 8892 4128
rect 7690 4097 7702 4100
rect 7644 4091 7702 4097
rect 3786 4060 3792 4072
rect 3436 4032 3792 4060
rect 3786 4020 3792 4032
rect 3844 4020 3850 4072
rect 7190 4060 7196 4072
rect 5000 4032 7196 4060
rect 2593 3927 2651 3933
rect 2593 3893 2605 3927
rect 2639 3924 2651 3927
rect 5000 3924 5028 4032
rect 7190 4020 7196 4032
rect 7248 4020 7254 4072
rect 5074 3952 5080 4004
rect 5132 3992 5138 4004
rect 6365 3995 6423 4001
rect 6365 3992 6377 3995
rect 5132 3964 6377 3992
rect 5132 3952 5138 3964
rect 6365 3961 6377 3964
rect 6411 3961 6423 3995
rect 6822 3992 6828 4004
rect 6783 3964 6828 3992
rect 6365 3955 6423 3961
rect 6822 3952 6828 3964
rect 6880 3952 6886 4004
rect 2639 3896 5028 3924
rect 5261 3927 5319 3933
rect 2639 3893 2651 3896
rect 2593 3887 2651 3893
rect 5261 3893 5273 3927
rect 5307 3924 5319 3927
rect 5718 3924 5724 3936
rect 5307 3896 5724 3924
rect 5307 3893 5319 3896
rect 5261 3887 5319 3893
rect 5718 3884 5724 3896
rect 5776 3924 5782 3936
rect 6638 3924 6644 3936
rect 5776 3896 6644 3924
rect 5776 3884 5782 3896
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 8754 3924 8760 3936
rect 8715 3896 8760 3924
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 8864 3924 8892 4100
rect 9217 4097 9229 4131
rect 9263 4097 9275 4131
rect 9217 4091 9275 4097
rect 9484 4091 9496 4137
rect 9548 4128 9554 4140
rect 10336 4128 10364 4156
rect 11422 4128 11428 4140
rect 9548 4100 9584 4128
rect 10336 4100 11428 4128
rect 9490 4088 9496 4091
rect 9548 4088 9554 4100
rect 11422 4088 11428 4100
rect 11480 4128 11486 4140
rect 11793 4131 11851 4137
rect 11793 4128 11805 4131
rect 11480 4100 11805 4128
rect 11480 4088 11486 4100
rect 11793 4097 11805 4100
rect 11839 4097 11851 4131
rect 13538 4128 13544 4140
rect 11793 4091 11851 4097
rect 11900 4100 13544 4128
rect 10410 4020 10416 4072
rect 10468 4060 10474 4072
rect 11900 4060 11928 4100
rect 13538 4088 13544 4100
rect 13596 4088 13602 4140
rect 13633 4131 13691 4137
rect 13633 4097 13645 4131
rect 13679 4128 13691 4131
rect 13832 4128 13860 4168
rect 14734 4156 14740 4168
rect 14792 4156 14798 4208
rect 15657 4199 15715 4205
rect 15657 4196 15669 4199
rect 14844 4168 15669 4196
rect 14844 4140 14872 4168
rect 15657 4165 15669 4168
rect 15703 4165 15715 4199
rect 19426 4196 19432 4208
rect 19387 4168 19432 4196
rect 15657 4159 15715 4165
rect 19426 4156 19432 4168
rect 19484 4156 19490 4208
rect 19619 4140 19647 4236
rect 19797 4233 19809 4267
rect 19843 4264 19855 4267
rect 19978 4264 19984 4276
rect 19843 4236 19984 4264
rect 19843 4233 19855 4236
rect 19797 4227 19855 4233
rect 19978 4224 19984 4236
rect 20036 4224 20042 4276
rect 21836 4236 22416 4264
rect 20346 4196 20352 4208
rect 20114 4168 20352 4196
rect 13906 4137 13912 4140
rect 13679 4100 13860 4128
rect 13679 4097 13691 4100
rect 13633 4091 13691 4097
rect 13900 4091 13912 4137
rect 13964 4128 13970 4140
rect 13964 4100 14000 4128
rect 13906 4088 13912 4091
rect 13964 4088 13970 4100
rect 14274 4088 14280 4140
rect 14332 4128 14338 4140
rect 14826 4128 14832 4140
rect 14332 4100 14832 4128
rect 14332 4088 14338 4100
rect 14826 4088 14832 4100
rect 14884 4088 14890 4140
rect 15286 4088 15292 4140
rect 15344 4128 15350 4140
rect 15470 4128 15476 4140
rect 15344 4100 15476 4128
rect 15344 4088 15350 4100
rect 15470 4088 15476 4100
rect 15528 4088 15534 4140
rect 15746 4128 15752 4140
rect 15707 4100 15752 4128
rect 15746 4088 15752 4100
rect 15804 4088 15810 4140
rect 15841 4131 15899 4137
rect 15841 4097 15853 4131
rect 15887 4097 15899 4131
rect 15841 4091 15899 4097
rect 10468 4032 11928 4060
rect 10468 4020 10474 4032
rect 10597 3995 10655 4001
rect 10597 3961 10609 3995
rect 10643 3992 10655 3995
rect 11054 3992 11060 4004
rect 10643 3964 11060 3992
rect 10643 3961 10655 3964
rect 10597 3955 10655 3961
rect 11054 3952 11060 3964
rect 11112 3992 11118 4004
rect 11606 3992 11612 4004
rect 11112 3964 11612 3992
rect 11112 3952 11118 3964
rect 11606 3952 11612 3964
rect 11664 3952 11670 4004
rect 13630 3992 13636 4004
rect 13096 3964 13636 3992
rect 9858 3924 9864 3936
rect 8864 3896 9864 3924
rect 9858 3884 9864 3896
rect 9916 3884 9922 3936
rect 9950 3884 9956 3936
rect 10008 3924 10014 3936
rect 13096 3924 13124 3964
rect 13630 3952 13636 3964
rect 13688 3952 13694 4004
rect 15654 3952 15660 4004
rect 15712 3992 15718 4004
rect 15856 3992 15884 4091
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 17293 4131 17351 4137
rect 17293 4128 17305 4131
rect 15988 4100 17305 4128
rect 15988 4088 15994 4100
rect 17293 4097 17305 4100
rect 17339 4097 17351 4131
rect 17293 4091 17351 4097
rect 19245 4131 19303 4137
rect 19245 4097 19257 4131
rect 19291 4097 19303 4131
rect 19245 4091 19303 4097
rect 19521 4131 19579 4137
rect 19521 4097 19533 4131
rect 19567 4097 19579 4131
rect 19521 4091 19579 4097
rect 17034 4060 17040 4072
rect 15712 3964 15884 3992
rect 16040 4032 17040 4060
rect 15712 3952 15718 3964
rect 10008 3896 13124 3924
rect 13173 3927 13231 3933
rect 10008 3884 10014 3896
rect 13173 3893 13185 3927
rect 13219 3924 13231 3927
rect 13814 3924 13820 3936
rect 13219 3896 13820 3924
rect 13219 3893 13231 3896
rect 13173 3887 13231 3893
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 16040 3924 16068 4032
rect 17034 4020 17040 4032
rect 17092 4020 17098 4072
rect 19260 4060 19288 4091
rect 19536 4060 19564 4091
rect 19610 4088 19616 4140
rect 19668 4128 19674 4140
rect 19668 4100 19761 4128
rect 19668 4088 19674 4100
rect 20114 4060 20142 4168
rect 20346 4156 20352 4168
rect 20404 4156 20410 4208
rect 20806 4196 20812 4208
rect 20456 4168 20812 4196
rect 20456 4137 20484 4168
rect 20806 4156 20812 4168
rect 20864 4156 20870 4208
rect 21836 4196 21864 4236
rect 22278 4196 22284 4208
rect 21744 4168 21864 4196
rect 22020 4168 22284 4196
rect 20441 4131 20499 4137
rect 20441 4097 20453 4131
rect 20487 4097 20499 4131
rect 20441 4091 20499 4097
rect 20530 4088 20536 4140
rect 20588 4128 20594 4140
rect 21269 4131 21327 4137
rect 21269 4128 21281 4131
rect 20588 4100 21281 4128
rect 20588 4088 20594 4100
rect 21269 4097 21281 4100
rect 21315 4097 21327 4131
rect 21269 4091 21327 4097
rect 20254 4060 20260 4072
rect 19260 4032 19472 4060
rect 19536 4032 20142 4060
rect 20215 4032 20260 4060
rect 19444 3992 19472 4032
rect 20254 4020 20260 4032
rect 20312 4020 20318 4072
rect 20346 4020 20352 4072
rect 20404 4060 20410 4072
rect 21744 4060 21772 4168
rect 21821 4131 21879 4137
rect 21821 4097 21833 4131
rect 21867 4128 21879 4131
rect 22020 4128 22048 4168
rect 22278 4156 22284 4168
rect 22336 4156 22342 4208
rect 22094 4137 22100 4140
rect 21867 4100 22048 4128
rect 21867 4097 21879 4100
rect 21821 4091 21879 4097
rect 22088 4091 22100 4137
rect 22152 4128 22158 4140
rect 22388 4128 22416 4236
rect 22462 4224 22468 4276
rect 22520 4264 22526 4276
rect 22646 4264 22652 4276
rect 22520 4236 22652 4264
rect 22520 4224 22526 4236
rect 22646 4224 22652 4236
rect 22704 4224 22710 4276
rect 23845 4267 23903 4273
rect 23845 4264 23857 4267
rect 23584 4236 23857 4264
rect 23584 4128 23612 4236
rect 23845 4233 23857 4236
rect 23891 4233 23903 4267
rect 33502 4264 33508 4276
rect 33463 4236 33508 4264
rect 23845 4227 23903 4233
rect 33502 4224 33508 4236
rect 33560 4224 33566 4276
rect 34790 4224 34796 4276
rect 34848 4264 34854 4276
rect 35802 4264 35808 4276
rect 34848 4236 35808 4264
rect 34848 4224 34854 4236
rect 35802 4224 35808 4236
rect 35860 4224 35866 4276
rect 25682 4196 25688 4208
rect 24780 4168 25688 4196
rect 22152 4100 22188 4128
rect 22388 4100 23612 4128
rect 23661 4131 23719 4137
rect 22094 4088 22100 4091
rect 22152 4088 22158 4100
rect 23661 4097 23673 4131
rect 23707 4128 23719 4131
rect 24673 4131 24731 4137
rect 23707 4100 24624 4128
rect 23707 4097 23719 4100
rect 23661 4091 23719 4097
rect 20404 4032 21772 4060
rect 20404 4020 20410 4032
rect 24394 4020 24400 4072
rect 24452 4060 24458 4072
rect 24489 4063 24547 4069
rect 24489 4060 24501 4063
rect 24452 4032 24501 4060
rect 24452 4020 24458 4032
rect 24489 4029 24501 4032
rect 24535 4029 24547 4063
rect 24596 4060 24624 4100
rect 24673 4097 24685 4131
rect 24719 4128 24731 4131
rect 24780 4128 24808 4168
rect 25682 4156 25688 4168
rect 25740 4156 25746 4208
rect 30006 4196 30012 4208
rect 27172 4168 27752 4196
rect 24719 4100 24808 4128
rect 24857 4131 24915 4137
rect 24719 4097 24731 4100
rect 24673 4091 24731 4097
rect 24857 4097 24869 4131
rect 24903 4128 24915 4131
rect 25314 4128 25320 4140
rect 24903 4100 25320 4128
rect 24903 4097 24915 4100
rect 24857 4091 24915 4097
rect 25314 4088 25320 4100
rect 25372 4088 25378 4140
rect 25501 4131 25559 4137
rect 25501 4097 25513 4131
rect 25547 4128 25559 4131
rect 25774 4128 25780 4140
rect 25547 4100 25780 4128
rect 25547 4097 25559 4100
rect 25501 4091 25559 4097
rect 25774 4088 25780 4100
rect 25832 4088 25838 4140
rect 26050 4128 26056 4140
rect 26011 4100 26056 4128
rect 26050 4088 26056 4100
rect 26108 4088 26114 4140
rect 26142 4088 26148 4140
rect 26200 4128 26206 4140
rect 26326 4128 26332 4140
rect 26200 4100 26245 4128
rect 26287 4100 26332 4128
rect 26200 4088 26206 4100
rect 26326 4088 26332 4100
rect 26384 4088 26390 4140
rect 27172 4128 27200 4168
rect 26436 4100 27200 4128
rect 27240 4131 27298 4137
rect 24946 4060 24952 4072
rect 24596 4032 24952 4060
rect 24489 4023 24547 4029
rect 24946 4020 24952 4032
rect 25004 4020 25010 4072
rect 19518 3992 19524 4004
rect 17972 3964 19334 3992
rect 19444 3964 19524 3992
rect 14792 3896 16068 3924
rect 14792 3884 14798 3896
rect 16114 3884 16120 3936
rect 16172 3924 16178 3936
rect 17972 3924 18000 3964
rect 16172 3896 18000 3924
rect 16172 3884 16178 3896
rect 18046 3884 18052 3936
rect 18104 3924 18110 3936
rect 18417 3927 18475 3933
rect 18417 3924 18429 3927
rect 18104 3896 18429 3924
rect 18104 3884 18110 3896
rect 18417 3893 18429 3896
rect 18463 3893 18475 3927
rect 19306 3924 19334 3964
rect 19518 3952 19524 3964
rect 19576 3952 19582 4004
rect 20625 3995 20683 4001
rect 20625 3992 20637 3995
rect 19812 3964 20637 3992
rect 19812 3924 19840 3964
rect 20625 3961 20637 3964
rect 20671 3961 20683 3995
rect 21266 3992 21272 4004
rect 20625 3955 20683 3961
rect 20732 3964 21272 3992
rect 19306 3896 19840 3924
rect 18417 3887 18475 3893
rect 20162 3884 20168 3936
rect 20220 3924 20226 3936
rect 20732 3924 20760 3964
rect 21266 3952 21272 3964
rect 21324 3952 21330 4004
rect 25317 3995 25375 4001
rect 25317 3992 25329 3995
rect 22756 3964 25329 3992
rect 20220 3896 20760 3924
rect 20220 3884 20226 3896
rect 20806 3884 20812 3936
rect 20864 3924 20870 3936
rect 21085 3927 21143 3933
rect 21085 3924 21097 3927
rect 20864 3896 21097 3924
rect 20864 3884 20870 3896
rect 21085 3893 21097 3896
rect 21131 3893 21143 3927
rect 21085 3887 21143 3893
rect 22094 3884 22100 3936
rect 22152 3924 22158 3936
rect 22756 3924 22784 3964
rect 25317 3961 25329 3964
rect 25363 3961 25375 3995
rect 26436 3992 26464 4100
rect 27240 4097 27252 4131
rect 27286 4128 27298 4131
rect 27614 4128 27620 4140
rect 27286 4100 27620 4128
rect 27286 4097 27298 4100
rect 27240 4091 27298 4097
rect 27614 4088 27620 4100
rect 27672 4088 27678 4140
rect 27724 4128 27752 4168
rect 28736 4168 30012 4196
rect 28736 4128 28764 4168
rect 30006 4156 30012 4168
rect 30064 4156 30070 4208
rect 30300 4168 31248 4196
rect 30300 4140 30328 4168
rect 27724 4100 28764 4128
rect 28813 4131 28871 4137
rect 28813 4097 28825 4131
rect 28859 4128 28871 4131
rect 29454 4128 29460 4140
rect 28859 4100 29460 4128
rect 28859 4097 28871 4100
rect 28813 4091 28871 4097
rect 29454 4088 29460 4100
rect 29512 4128 29518 4140
rect 29730 4128 29736 4140
rect 29512 4100 29736 4128
rect 29512 4088 29518 4100
rect 29730 4088 29736 4100
rect 29788 4088 29794 4140
rect 30282 4128 30288 4140
rect 30243 4100 30288 4128
rect 30282 4088 30288 4100
rect 30340 4088 30346 4140
rect 30466 4128 30472 4140
rect 30427 4100 30472 4128
rect 30466 4088 30472 4100
rect 30524 4088 30530 4140
rect 31220 4137 31248 4168
rect 36078 4156 36084 4208
rect 36136 4196 36142 4208
rect 36265 4199 36323 4205
rect 36265 4196 36277 4199
rect 36136 4168 36277 4196
rect 36136 4156 36142 4168
rect 36265 4165 36277 4168
rect 36311 4165 36323 4199
rect 36265 4159 36323 4165
rect 36354 4156 36360 4208
rect 36412 4196 36418 4208
rect 36465 4199 36523 4205
rect 36465 4196 36477 4199
rect 36412 4168 36477 4196
rect 36412 4156 36418 4168
rect 36465 4165 36477 4168
rect 36511 4165 36523 4199
rect 36465 4159 36523 4165
rect 30561 4131 30619 4137
rect 30561 4097 30573 4131
rect 30607 4097 30619 4131
rect 30561 4091 30619 4097
rect 31205 4131 31263 4137
rect 31205 4097 31217 4131
rect 31251 4097 31263 4131
rect 31386 4128 31392 4140
rect 31347 4100 31392 4128
rect 31205 4091 31263 4097
rect 26970 4060 26976 4072
rect 26931 4032 26976 4060
rect 26970 4020 26976 4032
rect 27028 4020 27034 4072
rect 28074 4020 28080 4072
rect 28132 4060 28138 4072
rect 28718 4060 28724 4072
rect 28132 4032 28724 4060
rect 28132 4020 28138 4032
rect 28718 4020 28724 4032
rect 28776 4020 28782 4072
rect 28994 4020 29000 4072
rect 29052 4060 29058 4072
rect 29089 4063 29147 4069
rect 29089 4060 29101 4063
rect 29052 4032 29101 4060
rect 29052 4020 29058 4032
rect 29089 4029 29101 4032
rect 29135 4060 29147 4063
rect 30190 4060 30196 4072
rect 29135 4032 30196 4060
rect 29135 4029 29147 4032
rect 29089 4023 29147 4029
rect 30190 4020 30196 4032
rect 30248 4060 30254 4072
rect 30576 4060 30604 4091
rect 31386 4088 31392 4100
rect 31444 4088 31450 4140
rect 31481 4131 31539 4137
rect 31481 4097 31493 4131
rect 31527 4097 31539 4131
rect 31481 4091 31539 4097
rect 32392 4131 32450 4137
rect 32392 4097 32404 4131
rect 32438 4128 32450 4131
rect 32674 4128 32680 4140
rect 32438 4100 32680 4128
rect 32438 4097 32450 4100
rect 32392 4091 32450 4097
rect 31496 4060 31524 4091
rect 32674 4088 32680 4100
rect 32732 4088 32738 4140
rect 34692 4131 34750 4137
rect 34692 4097 34704 4131
rect 34738 4128 34750 4131
rect 37826 4128 37832 4140
rect 34738 4100 36032 4128
rect 37787 4100 37832 4128
rect 34738 4097 34750 4100
rect 34692 4091 34750 4097
rect 30248 4032 31524 4060
rect 32125 4063 32183 4069
rect 30248 4020 30254 4032
rect 32125 4029 32137 4063
rect 32171 4029 32183 4063
rect 34422 4060 34428 4072
rect 34383 4032 34428 4060
rect 32125 4023 32183 4029
rect 30650 3992 30656 4004
rect 25317 3955 25375 3961
rect 25424 3964 26464 3992
rect 27908 3964 30656 3992
rect 23198 3924 23204 3936
rect 22152 3896 22784 3924
rect 23159 3896 23204 3924
rect 22152 3884 22158 3896
rect 23198 3884 23204 3896
rect 23256 3884 23262 3936
rect 23290 3884 23296 3936
rect 23348 3924 23354 3936
rect 25424 3924 25452 3964
rect 23348 3896 25452 3924
rect 23348 3884 23354 3896
rect 25866 3884 25872 3936
rect 25924 3924 25930 3936
rect 27908 3924 27936 3964
rect 30650 3952 30656 3964
rect 30708 3952 30714 4004
rect 32140 3936 32168 4023
rect 34422 4020 34428 4032
rect 34480 4020 34486 4072
rect 36004 4060 36032 4100
rect 37826 4088 37832 4100
rect 37884 4088 37890 4140
rect 37918 4060 37924 4072
rect 36004 4032 37924 4060
rect 37918 4020 37924 4032
rect 37976 4020 37982 4072
rect 34440 3992 34468 4020
rect 33060 3964 34468 3992
rect 36633 3995 36691 4001
rect 28350 3924 28356 3936
rect 25924 3896 27936 3924
rect 28311 3896 28356 3924
rect 25924 3884 25930 3896
rect 28350 3884 28356 3896
rect 28408 3884 28414 3936
rect 30098 3924 30104 3936
rect 30059 3896 30104 3924
rect 30098 3884 30104 3896
rect 30156 3884 30162 3936
rect 31018 3924 31024 3936
rect 30979 3896 31024 3924
rect 31018 3884 31024 3896
rect 31076 3884 31082 3936
rect 32122 3924 32128 3936
rect 32035 3896 32128 3924
rect 32122 3884 32128 3896
rect 32180 3924 32186 3936
rect 33060 3924 33088 3964
rect 36633 3961 36645 3995
rect 36679 3992 36691 3995
rect 37734 3992 37740 4004
rect 36679 3964 37740 3992
rect 36679 3961 36691 3964
rect 36633 3955 36691 3961
rect 37734 3952 37740 3964
rect 37792 3952 37798 4004
rect 36446 3924 36452 3936
rect 32180 3896 33088 3924
rect 36407 3896 36452 3924
rect 32180 3884 32186 3896
rect 36446 3884 36452 3896
rect 36504 3884 36510 3936
rect 38013 3927 38071 3933
rect 38013 3893 38025 3927
rect 38059 3924 38071 3927
rect 38286 3924 38292 3936
rect 38059 3896 38292 3924
rect 38059 3893 38071 3896
rect 38013 3887 38071 3893
rect 38286 3884 38292 3896
rect 38344 3884 38350 3936
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 2409 3723 2467 3729
rect 2409 3689 2421 3723
rect 2455 3720 2467 3723
rect 3694 3720 3700 3732
rect 2455 3692 3700 3720
rect 2455 3689 2467 3692
rect 2409 3683 2467 3689
rect 3694 3680 3700 3692
rect 3752 3680 3758 3732
rect 3789 3723 3847 3729
rect 3789 3689 3801 3723
rect 3835 3720 3847 3723
rect 7098 3720 7104 3732
rect 3835 3692 6592 3720
rect 7059 3692 7104 3720
rect 3835 3689 3847 3692
rect 3789 3683 3847 3689
rect 5258 3652 5264 3664
rect 3252 3624 5264 3652
rect 2608 3556 3188 3584
rect 1946 3516 1952 3528
rect 1907 3488 1952 3516
rect 1946 3476 1952 3488
rect 2004 3476 2010 3528
rect 2608 3525 2636 3556
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3485 2651 3519
rect 2593 3479 2651 3485
rect 2958 3448 2964 3460
rect 1780 3420 2964 3448
rect 1780 3389 1808 3420
rect 2958 3408 2964 3420
rect 3016 3408 3022 3460
rect 3160 3448 3188 3556
rect 3252 3525 3280 3624
rect 5258 3612 5264 3624
rect 5316 3612 5322 3664
rect 6564 3584 6592 3692
rect 7098 3680 7104 3692
rect 7156 3680 7162 3732
rect 7190 3680 7196 3732
rect 7248 3720 7254 3732
rect 8110 3720 8116 3732
rect 7248 3692 8116 3720
rect 7248 3680 7254 3692
rect 8110 3680 8116 3692
rect 8168 3680 8174 3732
rect 8205 3723 8263 3729
rect 8205 3689 8217 3723
rect 8251 3720 8263 3723
rect 9490 3720 9496 3732
rect 8251 3692 9496 3720
rect 8251 3689 8263 3692
rect 8205 3683 8263 3689
rect 9490 3680 9496 3692
rect 9548 3680 9554 3732
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 9916 3692 10456 3720
rect 9916 3680 9922 3692
rect 6641 3655 6699 3661
rect 6641 3621 6653 3655
rect 6687 3652 6699 3655
rect 7374 3652 7380 3664
rect 6687 3624 7380 3652
rect 6687 3621 6699 3624
rect 6641 3615 6699 3621
rect 7374 3612 7380 3624
rect 7432 3612 7438 3664
rect 9950 3652 9956 3664
rect 7484 3624 9956 3652
rect 7484 3584 7512 3624
rect 9950 3612 9956 3624
rect 10008 3612 10014 3664
rect 3988 3556 5212 3584
rect 6564 3556 7512 3584
rect 7561 3587 7619 3593
rect 3988 3525 4016 3556
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3485 3295 3519
rect 3237 3479 3295 3485
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 4433 3519 4491 3525
rect 4433 3485 4445 3519
rect 4479 3516 4491 3519
rect 5074 3516 5080 3528
rect 4479 3488 5080 3516
rect 4479 3485 4491 3488
rect 4433 3479 4491 3485
rect 5074 3476 5080 3488
rect 5132 3476 5138 3528
rect 4338 3448 4344 3460
rect 3160 3420 4344 3448
rect 4338 3408 4344 3420
rect 4396 3408 4402 3460
rect 4617 3451 4675 3457
rect 4617 3417 4629 3451
rect 4663 3417 4675 3451
rect 4617 3411 4675 3417
rect 1765 3383 1823 3389
rect 1765 3349 1777 3383
rect 1811 3349 1823 3383
rect 1765 3343 1823 3349
rect 3053 3383 3111 3389
rect 3053 3349 3065 3383
rect 3099 3380 3111 3383
rect 3970 3380 3976 3392
rect 3099 3352 3976 3380
rect 3099 3349 3111 3352
rect 3053 3343 3111 3349
rect 3970 3340 3976 3352
rect 4028 3340 4034 3392
rect 4062 3340 4068 3392
rect 4120 3380 4126 3392
rect 4632 3380 4660 3411
rect 4120 3352 4660 3380
rect 4801 3383 4859 3389
rect 4120 3340 4126 3352
rect 4801 3349 4813 3383
rect 4847 3380 4859 3383
rect 4890 3380 4896 3392
rect 4847 3352 4896 3380
rect 4847 3349 4859 3352
rect 4801 3343 4859 3349
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 5184 3380 5212 3556
rect 7561 3553 7573 3587
rect 7607 3584 7619 3587
rect 7926 3584 7932 3596
rect 7607 3556 7932 3584
rect 7607 3553 7619 3556
rect 7561 3547 7619 3553
rect 7926 3544 7932 3556
rect 7984 3544 7990 3596
rect 9030 3544 9036 3596
rect 9088 3584 9094 3596
rect 10428 3584 10456 3692
rect 10594 3680 10600 3732
rect 10652 3720 10658 3732
rect 10965 3723 11023 3729
rect 10965 3720 10977 3723
rect 10652 3692 10977 3720
rect 10652 3680 10658 3692
rect 10965 3689 10977 3692
rect 11011 3689 11023 3723
rect 10965 3683 11023 3689
rect 11330 3680 11336 3732
rect 11388 3720 11394 3732
rect 11977 3723 12035 3729
rect 11388 3692 11920 3720
rect 11388 3680 11394 3692
rect 11790 3612 11796 3664
rect 11848 3612 11854 3664
rect 11808 3584 11836 3612
rect 9088 3556 10364 3584
rect 10428 3556 10640 3584
rect 9088 3544 9094 3556
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3516 5319 3519
rect 5902 3516 5908 3528
rect 5307 3488 5908 3516
rect 5307 3485 5319 3488
rect 5261 3479 5319 3485
rect 5902 3476 5908 3488
rect 5960 3476 5966 3528
rect 7282 3516 7288 3528
rect 7243 3488 7288 3516
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 7374 3476 7380 3528
rect 7432 3516 7438 3528
rect 7653 3519 7711 3525
rect 7432 3488 7477 3516
rect 7432 3476 7438 3488
rect 7653 3485 7665 3519
rect 7699 3485 7711 3519
rect 7653 3479 7711 3485
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 5528 3451 5586 3457
rect 5528 3417 5540 3451
rect 5574 3448 5586 3451
rect 5626 3448 5632 3460
rect 5574 3420 5632 3448
rect 5574 3417 5586 3420
rect 5528 3411 5586 3417
rect 5626 3408 5632 3420
rect 5684 3408 5690 3460
rect 5718 3408 5724 3460
rect 5776 3448 5782 3460
rect 6454 3448 6460 3460
rect 5776 3420 6460 3448
rect 5776 3408 5782 3420
rect 6454 3408 6460 3420
rect 6512 3408 6518 3460
rect 6638 3408 6644 3460
rect 6696 3448 6702 3460
rect 7668 3448 7696 3479
rect 6696 3420 7696 3448
rect 8404 3448 8432 3479
rect 8570 3476 8576 3528
rect 8628 3516 8634 3528
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 8628 3488 9137 3516
rect 8628 3476 8634 3488
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9398 3516 9404 3528
rect 9359 3488 9404 3516
rect 9125 3479 9183 3485
rect 9398 3476 9404 3488
rect 9456 3516 9462 3528
rect 10226 3516 10232 3528
rect 9456 3488 10232 3516
rect 9456 3476 9462 3488
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 10336 3512 10364 3556
rect 10413 3519 10471 3525
rect 10413 3512 10425 3519
rect 10336 3485 10425 3512
rect 10459 3485 10471 3519
rect 10612 3516 10640 3556
rect 11532 3556 11836 3584
rect 10689 3519 10747 3525
rect 10689 3516 10701 3519
rect 10612 3488 10701 3516
rect 10336 3484 10471 3485
rect 10413 3479 10471 3484
rect 10689 3485 10701 3488
rect 10735 3485 10747 3519
rect 10689 3479 10747 3485
rect 10781 3519 10839 3525
rect 10781 3485 10793 3519
rect 10827 3516 10839 3519
rect 11330 3516 11336 3528
rect 10827 3488 11336 3516
rect 10827 3485 10839 3488
rect 10781 3479 10839 3485
rect 11330 3476 11336 3488
rect 11388 3476 11394 3528
rect 11445 3519 11503 3525
rect 11445 3485 11457 3519
rect 11491 3516 11503 3519
rect 11532 3516 11560 3556
rect 11698 3516 11704 3528
rect 11491 3488 11560 3516
rect 11659 3488 11704 3516
rect 11491 3485 11503 3488
rect 11445 3479 11503 3485
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 11793 3519 11851 3525
rect 11793 3485 11805 3519
rect 11839 3516 11851 3519
rect 11892 3516 11920 3692
rect 11977 3689 11989 3723
rect 12023 3720 12035 3723
rect 12158 3720 12164 3732
rect 12023 3692 12164 3720
rect 12023 3689 12035 3692
rect 11977 3683 12035 3689
rect 12158 3680 12164 3692
rect 12216 3680 12222 3732
rect 13078 3680 13084 3732
rect 13136 3720 13142 3732
rect 13541 3723 13599 3729
rect 13541 3720 13553 3723
rect 13136 3692 13553 3720
rect 13136 3680 13142 3692
rect 13541 3689 13553 3692
rect 13587 3689 13599 3723
rect 13541 3683 13599 3689
rect 13630 3680 13636 3732
rect 13688 3720 13694 3732
rect 15010 3720 15016 3732
rect 13688 3692 15016 3720
rect 13688 3680 13694 3692
rect 15010 3680 15016 3692
rect 15068 3680 15074 3732
rect 15470 3680 15476 3732
rect 15528 3720 15534 3732
rect 16209 3723 16267 3729
rect 16209 3720 16221 3723
rect 15528 3692 16221 3720
rect 15528 3680 15534 3692
rect 16209 3689 16221 3692
rect 16255 3689 16267 3723
rect 16209 3683 16267 3689
rect 17954 3680 17960 3732
rect 18012 3720 18018 3732
rect 18693 3723 18751 3729
rect 18693 3720 18705 3723
rect 18012 3692 18705 3720
rect 18012 3680 18018 3692
rect 18693 3689 18705 3692
rect 18739 3689 18751 3723
rect 18693 3683 18751 3689
rect 19610 3680 19616 3732
rect 19668 3720 19674 3732
rect 19668 3692 20760 3720
rect 19668 3680 19674 3692
rect 18874 3612 18880 3664
rect 18932 3652 18938 3664
rect 20622 3652 20628 3664
rect 18932 3624 20628 3652
rect 18932 3612 18938 3624
rect 20622 3612 20628 3624
rect 20680 3612 20686 3664
rect 20732 3652 20760 3692
rect 21266 3680 21272 3732
rect 21324 3720 21330 3732
rect 23198 3720 23204 3732
rect 21324 3692 23204 3720
rect 21324 3680 21330 3692
rect 23198 3680 23204 3692
rect 23256 3680 23262 3732
rect 25130 3680 25136 3732
rect 25188 3720 25194 3732
rect 25498 3720 25504 3732
rect 25188 3692 25504 3720
rect 25188 3680 25194 3692
rect 25498 3680 25504 3692
rect 25556 3680 25562 3732
rect 25961 3723 26019 3729
rect 25961 3689 25973 3723
rect 26007 3720 26019 3723
rect 27338 3720 27344 3732
rect 26007 3692 27344 3720
rect 26007 3689 26019 3692
rect 25961 3683 26019 3689
rect 27338 3680 27344 3692
rect 27396 3680 27402 3732
rect 27522 3680 27528 3732
rect 27580 3720 27586 3732
rect 30006 3720 30012 3732
rect 27580 3692 30012 3720
rect 27580 3680 27586 3692
rect 30006 3680 30012 3692
rect 30064 3680 30070 3732
rect 30466 3680 30472 3732
rect 30524 3720 30530 3732
rect 31113 3723 31171 3729
rect 31113 3720 31125 3723
rect 30524 3692 31125 3720
rect 30524 3680 30530 3692
rect 31113 3689 31125 3692
rect 31159 3689 31171 3723
rect 31113 3683 31171 3689
rect 31757 3723 31815 3729
rect 31757 3689 31769 3723
rect 31803 3689 31815 3723
rect 31757 3683 31815 3689
rect 31941 3723 31999 3729
rect 31941 3689 31953 3723
rect 31987 3720 31999 3723
rect 32030 3720 32036 3732
rect 31987 3692 32036 3720
rect 31987 3689 31999 3692
rect 31941 3683 31999 3689
rect 22186 3652 22192 3664
rect 20732 3624 22192 3652
rect 14090 3584 14096 3596
rect 13372 3556 14096 3584
rect 11839 3488 11920 3516
rect 12989 3519 13047 3525
rect 11839 3485 11851 3488
rect 11793 3479 11851 3485
rect 12989 3485 13001 3519
rect 13035 3485 13047 3519
rect 12989 3479 13047 3485
rect 10042 3448 10048 3460
rect 8404 3420 10048 3448
rect 6696 3408 6702 3420
rect 10042 3408 10048 3420
rect 10100 3408 10106 3460
rect 10594 3448 10600 3460
rect 10555 3420 10600 3448
rect 10594 3408 10600 3420
rect 10652 3448 10658 3460
rect 11609 3451 11667 3457
rect 11609 3448 11621 3451
rect 10652 3420 11621 3448
rect 10652 3408 10658 3420
rect 11609 3417 11621 3420
rect 11655 3417 11667 3451
rect 11609 3411 11667 3417
rect 11974 3408 11980 3460
rect 12032 3448 12038 3460
rect 12032 3420 12434 3448
rect 12032 3408 12038 3420
rect 12158 3380 12164 3392
rect 5184 3352 12164 3380
rect 12158 3340 12164 3352
rect 12216 3340 12222 3392
rect 12406 3380 12434 3420
rect 12894 3380 12900 3392
rect 12406 3352 12900 3380
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 13004 3380 13032 3479
rect 13078 3476 13084 3528
rect 13136 3516 13142 3528
rect 13372 3525 13400 3556
rect 14090 3544 14096 3556
rect 14148 3584 14154 3596
rect 14458 3584 14464 3596
rect 14148 3556 14464 3584
rect 14148 3544 14154 3556
rect 14458 3544 14464 3556
rect 14516 3544 14522 3596
rect 14734 3544 14740 3596
rect 14792 3584 14798 3596
rect 14829 3587 14887 3593
rect 14829 3584 14841 3587
rect 14792 3556 14841 3584
rect 14792 3544 14798 3556
rect 14829 3553 14841 3556
rect 14875 3553 14887 3587
rect 14829 3547 14887 3553
rect 17034 3544 17040 3596
rect 17092 3584 17098 3596
rect 17313 3587 17371 3593
rect 17313 3584 17325 3587
rect 17092 3556 17325 3584
rect 17092 3544 17098 3556
rect 17313 3553 17325 3556
rect 17359 3553 17371 3587
rect 17313 3547 17371 3553
rect 19245 3587 19303 3593
rect 19245 3553 19257 3587
rect 19291 3584 19303 3587
rect 20254 3584 20260 3596
rect 19291 3556 20260 3584
rect 19291 3553 19303 3556
rect 19245 3547 19303 3553
rect 20254 3544 20260 3556
rect 20312 3544 20318 3596
rect 13265 3519 13323 3525
rect 13265 3516 13277 3519
rect 13136 3488 13277 3516
rect 13136 3476 13142 3488
rect 13265 3485 13277 3488
rect 13311 3485 13323 3519
rect 13265 3479 13323 3485
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3485 13415 3519
rect 14274 3516 14280 3528
rect 13357 3479 13415 3485
rect 13464 3488 14280 3516
rect 13173 3451 13231 3457
rect 13173 3417 13185 3451
rect 13219 3448 13231 3451
rect 13464 3448 13492 3488
rect 14274 3476 14280 3488
rect 14332 3476 14338 3528
rect 14369 3519 14427 3525
rect 14369 3485 14381 3519
rect 14415 3516 14427 3519
rect 16022 3516 16028 3528
rect 14415 3488 16028 3516
rect 14415 3485 14427 3488
rect 14369 3479 14427 3485
rect 16022 3476 16028 3488
rect 16080 3476 16086 3528
rect 16853 3519 16911 3525
rect 16853 3485 16865 3519
rect 16899 3516 16911 3519
rect 19426 3516 19432 3528
rect 16899 3488 18276 3516
rect 19387 3488 19432 3516
rect 16899 3485 16911 3488
rect 16853 3479 16911 3485
rect 13538 3448 13544 3460
rect 13219 3420 13544 3448
rect 13219 3417 13231 3420
rect 13173 3411 13231 3417
rect 13538 3408 13544 3420
rect 13596 3408 13602 3460
rect 13722 3408 13728 3460
rect 13780 3448 13786 3460
rect 15074 3451 15132 3457
rect 15074 3448 15086 3451
rect 13780 3420 15086 3448
rect 13780 3408 13786 3420
rect 15074 3417 15086 3420
rect 15120 3417 15132 3451
rect 15074 3411 15132 3417
rect 15194 3408 15200 3460
rect 15252 3448 15258 3460
rect 17558 3451 17616 3457
rect 17558 3448 17570 3451
rect 15252 3420 17570 3448
rect 15252 3408 15258 3420
rect 17558 3417 17570 3420
rect 17604 3417 17616 3451
rect 18248 3448 18276 3488
rect 19426 3476 19432 3488
rect 19484 3476 19490 3528
rect 20162 3476 20168 3528
rect 20220 3516 20226 3528
rect 20533 3519 20591 3525
rect 20533 3516 20545 3519
rect 20220 3488 20545 3516
rect 20220 3476 20226 3488
rect 20533 3485 20545 3488
rect 20579 3485 20591 3519
rect 20732 3516 20760 3624
rect 22186 3612 22192 3624
rect 22244 3612 22250 3664
rect 25869 3655 25927 3661
rect 23492 3624 25636 3652
rect 21637 3587 21695 3593
rect 21637 3553 21649 3587
rect 21683 3584 21695 3587
rect 21910 3584 21916 3596
rect 21683 3556 21916 3584
rect 21683 3553 21695 3556
rect 21637 3547 21695 3553
rect 21910 3544 21916 3556
rect 21968 3544 21974 3596
rect 22278 3544 22284 3596
rect 22336 3584 22342 3596
rect 22465 3587 22523 3593
rect 22465 3584 22477 3587
rect 22336 3556 22477 3584
rect 22336 3544 22342 3556
rect 22465 3553 22477 3556
rect 22511 3553 22523 3587
rect 22465 3547 22523 3553
rect 20901 3519 20959 3525
rect 20901 3516 20913 3519
rect 20732 3488 20913 3516
rect 20533 3479 20591 3485
rect 20901 3485 20913 3488
rect 20947 3485 20959 3519
rect 20901 3479 20959 3485
rect 21082 3476 21088 3528
rect 21140 3516 21146 3528
rect 21726 3516 21732 3528
rect 21140 3488 21732 3516
rect 21140 3476 21146 3488
rect 21726 3476 21732 3488
rect 21784 3476 21790 3528
rect 21821 3519 21879 3525
rect 21821 3485 21833 3519
rect 21867 3516 21879 3519
rect 22002 3516 22008 3528
rect 21867 3488 22008 3516
rect 21867 3485 21879 3488
rect 21821 3479 21879 3485
rect 22002 3476 22008 3488
rect 22060 3476 22066 3528
rect 22664 3516 22784 3518
rect 23492 3516 23520 3624
rect 24394 3584 24400 3596
rect 24355 3556 24400 3584
rect 24394 3544 24400 3556
rect 24452 3544 24458 3596
rect 25038 3544 25044 3596
rect 25096 3584 25102 3596
rect 25501 3587 25559 3593
rect 25501 3584 25513 3587
rect 25096 3556 25513 3584
rect 25096 3544 25102 3556
rect 25501 3553 25513 3556
rect 25547 3553 25559 3587
rect 25608 3584 25636 3624
rect 25869 3621 25881 3655
rect 25915 3652 25927 3655
rect 26050 3652 26056 3664
rect 25915 3624 26056 3652
rect 25915 3621 25927 3624
rect 25869 3615 25927 3621
rect 26050 3612 26056 3624
rect 26108 3612 26114 3664
rect 31772 3652 31800 3683
rect 32030 3680 32036 3692
rect 32088 3680 32094 3732
rect 32585 3723 32643 3729
rect 32585 3720 32597 3723
rect 32324 3692 32597 3720
rect 32324 3664 32352 3692
rect 32585 3689 32597 3692
rect 32631 3720 32643 3723
rect 33413 3723 33471 3729
rect 33413 3720 33425 3723
rect 32631 3692 33425 3720
rect 32631 3689 32643 3692
rect 32585 3683 32643 3689
rect 33413 3689 33425 3692
rect 33459 3689 33471 3723
rect 33413 3683 33471 3689
rect 33597 3723 33655 3729
rect 33597 3689 33609 3723
rect 33643 3720 33655 3723
rect 34514 3720 34520 3732
rect 33643 3692 34520 3720
rect 33643 3689 33655 3692
rect 33597 3683 33655 3689
rect 34514 3680 34520 3692
rect 34572 3680 34578 3732
rect 36446 3680 36452 3732
rect 36504 3720 36510 3732
rect 36725 3723 36783 3729
rect 36725 3720 36737 3723
rect 36504 3692 36737 3720
rect 36504 3680 36510 3692
rect 36725 3689 36737 3692
rect 36771 3689 36783 3723
rect 36906 3720 36912 3732
rect 36867 3692 36912 3720
rect 36725 3683 36783 3689
rect 36906 3680 36912 3692
rect 36964 3680 36970 3732
rect 32306 3652 32312 3664
rect 31772 3624 32312 3652
rect 32306 3612 32312 3624
rect 32364 3612 32370 3664
rect 32769 3655 32827 3661
rect 32769 3621 32781 3655
rect 32815 3652 32827 3655
rect 34606 3652 34612 3664
rect 32815 3624 34612 3652
rect 32815 3621 32827 3624
rect 32769 3615 32827 3621
rect 34606 3612 34612 3624
rect 34664 3612 34670 3664
rect 26878 3584 26884 3596
rect 25608 3556 26884 3584
rect 25501 3547 25559 3553
rect 26878 3544 26884 3556
rect 26936 3544 26942 3596
rect 26970 3544 26976 3596
rect 27028 3584 27034 3596
rect 27157 3587 27215 3593
rect 27157 3584 27169 3587
rect 27028 3556 27169 3584
rect 27028 3544 27034 3556
rect 27157 3553 27169 3556
rect 27203 3553 27215 3587
rect 27157 3547 27215 3553
rect 24578 3516 24584 3528
rect 22664 3510 22876 3516
rect 22940 3510 23520 3516
rect 22664 3490 23520 3510
rect 19613 3451 19671 3457
rect 19613 3448 19625 3451
rect 18248 3420 19625 3448
rect 17558 3411 17616 3417
rect 19613 3417 19625 3420
rect 19659 3417 19671 3451
rect 19613 3411 19671 3417
rect 19794 3408 19800 3460
rect 19852 3448 19858 3460
rect 20622 3448 20628 3460
rect 19852 3420 20628 3448
rect 19852 3408 19858 3420
rect 20622 3408 20628 3420
rect 20680 3448 20686 3460
rect 20717 3451 20775 3457
rect 20717 3448 20729 3451
rect 20680 3420 20729 3448
rect 20680 3408 20686 3420
rect 20717 3417 20729 3420
rect 20763 3417 20775 3451
rect 20717 3411 20775 3417
rect 20809 3451 20867 3457
rect 20809 3417 20821 3451
rect 20855 3448 20867 3451
rect 22664 3448 22692 3490
rect 22756 3488 23520 3490
rect 24539 3488 24584 3516
rect 22848 3482 22968 3488
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 24765 3519 24823 3525
rect 24765 3485 24777 3519
rect 24811 3516 24823 3519
rect 26234 3516 26240 3528
rect 24811 3488 26240 3516
rect 24811 3485 24823 3488
rect 24765 3479 24823 3485
rect 26234 3476 26240 3488
rect 26292 3476 26298 3528
rect 26418 3516 26424 3528
rect 26379 3488 26424 3516
rect 26418 3476 26424 3488
rect 26476 3476 26482 3528
rect 27172 3516 27200 3547
rect 30742 3544 30748 3596
rect 30800 3584 30806 3596
rect 33410 3584 33416 3596
rect 30800 3556 33416 3584
rect 30800 3544 30806 3556
rect 33410 3544 33416 3556
rect 33468 3544 33474 3596
rect 34422 3544 34428 3596
rect 34480 3584 34486 3596
rect 34701 3587 34759 3593
rect 34701 3584 34713 3587
rect 34480 3556 34713 3584
rect 34480 3544 34486 3556
rect 34701 3553 34713 3556
rect 34747 3553 34759 3587
rect 34701 3547 34759 3553
rect 29730 3516 29736 3528
rect 27172 3488 29736 3516
rect 29730 3476 29736 3488
rect 29788 3516 29794 3528
rect 32122 3516 32128 3528
rect 29788 3488 32128 3516
rect 29788 3476 29794 3488
rect 32122 3476 32128 3488
rect 32180 3476 32186 3528
rect 33502 3476 33508 3528
rect 33560 3476 33566 3528
rect 34968 3519 35026 3525
rect 34968 3485 34980 3519
rect 35014 3516 35026 3519
rect 35434 3516 35440 3528
rect 35014 3488 35440 3516
rect 35014 3485 35026 3488
rect 34968 3479 35026 3485
rect 35434 3476 35440 3488
rect 35492 3476 35498 3528
rect 37458 3476 37464 3528
rect 37516 3516 37522 3528
rect 37645 3519 37703 3525
rect 37645 3516 37657 3519
rect 37516 3488 37657 3516
rect 37516 3476 37522 3488
rect 37645 3485 37657 3488
rect 37691 3485 37703 3519
rect 37645 3479 37703 3485
rect 22738 3457 22744 3460
rect 20855 3420 22692 3448
rect 20855 3417 20867 3420
rect 20809 3411 20867 3417
rect 22732 3411 22744 3457
rect 22796 3448 22802 3460
rect 22796 3420 22832 3448
rect 22738 3408 22744 3411
rect 22796 3408 22802 3420
rect 23106 3408 23112 3460
rect 23164 3448 23170 3460
rect 27424 3451 27482 3457
rect 23164 3420 26740 3448
rect 23164 3408 23170 3420
rect 13814 3380 13820 3392
rect 13004 3352 13820 3380
rect 13814 3340 13820 3352
rect 13872 3340 13878 3392
rect 14185 3383 14243 3389
rect 14185 3349 14197 3383
rect 14231 3380 14243 3383
rect 15930 3380 15936 3392
rect 14231 3352 15936 3380
rect 14231 3349 14243 3352
rect 14185 3343 14243 3349
rect 15930 3340 15936 3352
rect 15988 3340 15994 3392
rect 16669 3383 16727 3389
rect 16669 3349 16681 3383
rect 16715 3380 16727 3383
rect 18598 3380 18604 3392
rect 16715 3352 18604 3380
rect 16715 3349 16727 3352
rect 16669 3343 16727 3349
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 20898 3380 20904 3392
rect 19484 3352 20904 3380
rect 19484 3340 19490 3352
rect 20898 3340 20904 3352
rect 20956 3340 20962 3392
rect 21085 3383 21143 3389
rect 21085 3349 21097 3383
rect 21131 3380 21143 3383
rect 21266 3380 21272 3392
rect 21131 3352 21272 3380
rect 21131 3349 21143 3352
rect 21085 3343 21143 3349
rect 21266 3340 21272 3352
rect 21324 3340 21330 3392
rect 22005 3383 22063 3389
rect 22005 3349 22017 3383
rect 22051 3380 22063 3383
rect 23658 3380 23664 3392
rect 22051 3352 23664 3380
rect 22051 3349 22063 3352
rect 22005 3343 22063 3349
rect 23658 3340 23664 3352
rect 23716 3340 23722 3392
rect 23842 3380 23848 3392
rect 23803 3352 23848 3380
rect 23842 3340 23848 3352
rect 23900 3340 23906 3392
rect 26326 3340 26332 3392
rect 26384 3380 26390 3392
rect 26605 3383 26663 3389
rect 26605 3380 26617 3383
rect 26384 3352 26617 3380
rect 26384 3340 26390 3352
rect 26605 3349 26617 3352
rect 26651 3349 26663 3383
rect 26712 3380 26740 3420
rect 27424 3417 27436 3451
rect 27470 3448 27482 3451
rect 28442 3448 28448 3460
rect 27470 3420 28448 3448
rect 27470 3417 27482 3420
rect 27424 3411 27482 3417
rect 28442 3408 28448 3420
rect 28500 3408 28506 3460
rect 30000 3451 30058 3457
rect 30000 3417 30012 3451
rect 30046 3448 30058 3451
rect 30098 3448 30104 3460
rect 30046 3420 30104 3448
rect 30046 3417 30058 3420
rect 30000 3411 30058 3417
rect 30098 3408 30104 3420
rect 30156 3408 30162 3460
rect 30466 3408 30472 3460
rect 30524 3448 30530 3460
rect 31573 3451 31631 3457
rect 31573 3448 31585 3451
rect 30524 3420 31585 3448
rect 30524 3408 30530 3420
rect 31573 3417 31585 3420
rect 31619 3417 31631 3451
rect 32398 3448 32404 3460
rect 32359 3420 32404 3448
rect 31573 3411 31631 3417
rect 32398 3408 32404 3420
rect 32456 3408 32462 3460
rect 33229 3451 33287 3457
rect 33229 3417 33241 3451
rect 33275 3448 33287 3451
rect 33520 3448 33548 3476
rect 33275 3420 33548 3448
rect 33275 3417 33287 3420
rect 33229 3411 33287 3417
rect 35618 3408 35624 3460
rect 35676 3448 35682 3460
rect 36541 3451 36599 3457
rect 36541 3448 36553 3451
rect 35676 3420 36553 3448
rect 35676 3408 35682 3420
rect 36541 3417 36553 3420
rect 36587 3417 36599 3451
rect 36541 3411 36599 3417
rect 27522 3380 27528 3392
rect 26712 3352 27528 3380
rect 26605 3343 26663 3349
rect 27522 3340 27528 3352
rect 27580 3340 27586 3392
rect 28537 3383 28595 3389
rect 28537 3349 28549 3383
rect 28583 3380 28595 3383
rect 28810 3380 28816 3392
rect 28583 3352 28816 3380
rect 28583 3349 28595 3352
rect 28537 3343 28595 3349
rect 28810 3340 28816 3352
rect 28868 3340 28874 3392
rect 29362 3340 29368 3392
rect 29420 3380 29426 3392
rect 31294 3380 31300 3392
rect 29420 3352 31300 3380
rect 29420 3340 29426 3352
rect 31294 3340 31300 3352
rect 31352 3340 31358 3392
rect 31783 3383 31841 3389
rect 31783 3349 31795 3383
rect 31829 3380 31841 3383
rect 32214 3380 32220 3392
rect 31829 3352 32220 3380
rect 31829 3349 31841 3352
rect 31783 3343 31841 3349
rect 32214 3340 32220 3352
rect 32272 3380 32278 3392
rect 32611 3383 32669 3389
rect 32611 3380 32623 3383
rect 32272 3352 32623 3380
rect 32272 3340 32278 3352
rect 32611 3349 32623 3352
rect 32657 3380 32669 3383
rect 33439 3383 33497 3389
rect 33439 3380 33451 3383
rect 32657 3352 33451 3380
rect 32657 3349 32669 3352
rect 32611 3343 32669 3349
rect 33439 3349 33451 3352
rect 33485 3380 33497 3383
rect 33962 3380 33968 3392
rect 33485 3352 33968 3380
rect 33485 3349 33497 3352
rect 33439 3343 33497 3349
rect 33962 3340 33968 3352
rect 34020 3340 34026 3392
rect 34330 3340 34336 3392
rect 34388 3380 34394 3392
rect 35342 3380 35348 3392
rect 34388 3352 35348 3380
rect 34388 3340 34394 3352
rect 35342 3340 35348 3352
rect 35400 3380 35406 3392
rect 36081 3383 36139 3389
rect 36081 3380 36093 3383
rect 35400 3352 36093 3380
rect 35400 3340 35406 3352
rect 36081 3349 36093 3352
rect 36127 3349 36139 3383
rect 36081 3343 36139 3349
rect 36354 3340 36360 3392
rect 36412 3380 36418 3392
rect 36741 3383 36799 3389
rect 36741 3380 36753 3383
rect 36412 3352 36753 3380
rect 36412 3340 36418 3352
rect 36741 3349 36753 3352
rect 36787 3349 36799 3383
rect 36741 3343 36799 3349
rect 37550 3340 37556 3392
rect 37608 3380 37614 3392
rect 37829 3383 37887 3389
rect 37829 3380 37841 3383
rect 37608 3352 37841 3380
rect 37608 3340 37614 3352
rect 37829 3349 37841 3352
rect 37875 3349 37887 3383
rect 37829 3343 37887 3349
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 1765 3179 1823 3185
rect 1765 3145 1777 3179
rect 1811 3145 1823 3179
rect 1765 3139 1823 3145
rect 1780 3108 1808 3139
rect 2958 3136 2964 3188
rect 3016 3176 3022 3188
rect 4246 3176 4252 3188
rect 3016 3148 4252 3176
rect 3016 3136 3022 3148
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 4341 3179 4399 3185
rect 4341 3145 4353 3179
rect 4387 3176 4399 3179
rect 4614 3176 4620 3188
rect 4387 3148 4620 3176
rect 4387 3145 4399 3148
rect 4341 3139 4399 3145
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 5626 3176 5632 3188
rect 5587 3148 5632 3176
rect 5626 3136 5632 3148
rect 5684 3136 5690 3188
rect 8018 3176 8024 3188
rect 7979 3148 8024 3176
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 8168 3148 10456 3176
rect 8168 3136 8174 3148
rect 9950 3108 9956 3120
rect 1780 3080 6408 3108
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3009 2007 3043
rect 1949 3003 2007 3009
rect 2593 3043 2651 3049
rect 2593 3009 2605 3043
rect 2639 3040 2651 3043
rect 3050 3040 3056 3052
rect 2639 3012 3056 3040
rect 2639 3009 2651 3012
rect 2593 3003 2651 3009
rect 1964 2972 1992 3003
rect 3050 3000 3056 3012
rect 3108 3000 3114 3052
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3040 3295 3043
rect 3786 3040 3792 3052
rect 3283 3012 3792 3040
rect 3283 3009 3295 3012
rect 3237 3003 3295 3009
rect 3786 3000 3792 3012
rect 3844 3000 3850 3052
rect 3881 3043 3939 3049
rect 3881 3009 3893 3043
rect 3927 3040 3939 3043
rect 4154 3040 4160 3052
rect 3927 3012 4160 3040
rect 3927 3009 3939 3012
rect 3881 3003 3939 3009
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 4525 3043 4583 3049
rect 4525 3009 4537 3043
rect 4571 3040 4583 3043
rect 4890 3040 4896 3052
rect 4571 3012 4896 3040
rect 4571 3009 4583 3012
rect 4525 3003 4583 3009
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 5169 3043 5227 3049
rect 5169 3009 5181 3043
rect 5215 3040 5227 3043
rect 5718 3040 5724 3052
rect 5215 3012 5724 3040
rect 5215 3009 5227 3012
rect 5169 3003 5227 3009
rect 5718 3000 5724 3012
rect 5776 3000 5782 3052
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 5994 3040 6000 3052
rect 5859 3012 6000 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 5994 3000 6000 3012
rect 6052 3000 6058 3052
rect 6380 3040 6408 3080
rect 6564 3080 9956 3108
rect 6564 3040 6592 3080
rect 9950 3068 9956 3080
rect 10008 3068 10014 3120
rect 10428 3117 10456 3148
rect 12894 3136 12900 3188
rect 12952 3176 12958 3188
rect 15746 3176 15752 3188
rect 12952 3148 15752 3176
rect 12952 3136 12958 3148
rect 15746 3136 15752 3148
rect 15804 3136 15810 3188
rect 15933 3179 15991 3185
rect 15933 3145 15945 3179
rect 15979 3176 15991 3179
rect 16574 3176 16580 3188
rect 15979 3148 16580 3176
rect 15979 3145 15991 3148
rect 15933 3139 15991 3145
rect 16574 3136 16580 3148
rect 16632 3136 16638 3188
rect 18414 3136 18420 3188
rect 18472 3176 18478 3188
rect 18509 3179 18567 3185
rect 18509 3176 18521 3179
rect 18472 3148 18521 3176
rect 18472 3136 18478 3148
rect 18509 3145 18521 3148
rect 18555 3145 18567 3179
rect 18509 3139 18567 3145
rect 19889 3179 19947 3185
rect 19889 3145 19901 3179
rect 19935 3176 19947 3179
rect 20530 3176 20536 3188
rect 19935 3148 20536 3176
rect 19935 3145 19947 3148
rect 19889 3139 19947 3145
rect 20530 3136 20536 3148
rect 20588 3136 20594 3188
rect 20714 3176 20720 3188
rect 20675 3148 20720 3176
rect 20714 3136 20720 3148
rect 20772 3136 20778 3188
rect 21726 3136 21732 3188
rect 21784 3176 21790 3188
rect 23842 3176 23848 3188
rect 21784 3148 23848 3176
rect 21784 3136 21790 3148
rect 23842 3136 23848 3148
rect 23900 3136 23906 3188
rect 24486 3176 24492 3188
rect 24447 3148 24492 3176
rect 24486 3136 24492 3148
rect 24544 3136 24550 3188
rect 25590 3136 25596 3188
rect 25648 3176 25654 3188
rect 25777 3179 25835 3185
rect 25777 3176 25789 3179
rect 25648 3148 25789 3176
rect 25648 3136 25654 3148
rect 25777 3145 25789 3148
rect 25823 3145 25835 3179
rect 27798 3176 27804 3188
rect 27759 3148 27804 3176
rect 25777 3139 25835 3145
rect 27798 3136 27804 3148
rect 27856 3136 27862 3188
rect 28074 3136 28080 3188
rect 28132 3176 28138 3188
rect 28655 3179 28713 3185
rect 28655 3176 28667 3179
rect 28132 3148 28667 3176
rect 28132 3136 28138 3148
rect 28655 3145 28667 3148
rect 28701 3176 28713 3179
rect 28902 3176 28908 3188
rect 28701 3148 28908 3176
rect 28701 3145 28713 3148
rect 28655 3139 28713 3145
rect 28902 3136 28908 3148
rect 28960 3176 28966 3188
rect 29473 3179 29531 3185
rect 29473 3176 29485 3179
rect 28960 3148 29485 3176
rect 28960 3136 28966 3148
rect 29473 3145 29485 3148
rect 29519 3145 29531 3179
rect 29473 3139 29531 3145
rect 29641 3179 29699 3185
rect 29641 3145 29653 3179
rect 29687 3176 29699 3179
rect 30742 3176 30748 3188
rect 29687 3148 30748 3176
rect 29687 3145 29699 3148
rect 29641 3139 29699 3145
rect 30742 3136 30748 3148
rect 30800 3136 30806 3188
rect 31386 3136 31392 3188
rect 31444 3176 31450 3188
rect 31481 3179 31539 3185
rect 31481 3176 31493 3179
rect 31444 3148 31493 3176
rect 31444 3136 31450 3148
rect 31481 3145 31493 3148
rect 31527 3176 31539 3179
rect 31527 3148 31754 3176
rect 31527 3145 31539 3148
rect 31481 3139 31539 3145
rect 10413 3111 10471 3117
rect 10413 3077 10425 3111
rect 10459 3077 10471 3111
rect 10413 3071 10471 3077
rect 10778 3068 10784 3120
rect 10836 3108 10842 3120
rect 14734 3108 14740 3120
rect 10836 3080 14740 3108
rect 10836 3068 10842 3080
rect 14734 3068 14740 3080
rect 14792 3068 14798 3120
rect 15286 3068 15292 3120
rect 15344 3108 15350 3120
rect 15562 3108 15568 3120
rect 15344 3080 15568 3108
rect 15344 3068 15350 3080
rect 15562 3068 15568 3080
rect 15620 3068 15626 3120
rect 18230 3108 18236 3120
rect 18191 3080 18236 3108
rect 18230 3068 18236 3080
rect 18288 3068 18294 3120
rect 20622 3108 20628 3120
rect 19076 3080 20628 3108
rect 6380 3012 6592 3040
rect 6641 3043 6699 3049
rect 6641 3009 6653 3043
rect 6687 3009 6699 3043
rect 6641 3003 6699 3009
rect 6908 3043 6966 3049
rect 6908 3009 6920 3043
rect 6954 3040 6966 3043
rect 7374 3040 7380 3052
rect 6954 3012 7380 3040
rect 6954 3009 6966 3012
rect 6908 3003 6966 3009
rect 2958 2972 2964 2984
rect 1964 2944 2964 2972
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 5902 2932 5908 2984
rect 5960 2972 5966 2984
rect 6656 2972 6684 3003
rect 7374 3000 7380 3012
rect 7432 3000 7438 3052
rect 10042 3040 10048 3052
rect 7668 3012 10048 3040
rect 5960 2944 6684 2972
rect 5960 2932 5966 2944
rect 3053 2907 3111 2913
rect 3053 2873 3065 2907
rect 3099 2904 3111 2907
rect 6638 2904 6644 2916
rect 3099 2876 6644 2904
rect 3099 2873 3111 2876
rect 3053 2867 3111 2873
rect 6638 2864 6644 2876
rect 6696 2864 6702 2916
rect 2409 2839 2467 2845
rect 2409 2805 2421 2839
rect 2455 2836 2467 2839
rect 3418 2836 3424 2848
rect 2455 2808 3424 2836
rect 2455 2805 2467 2808
rect 2409 2799 2467 2805
rect 3418 2796 3424 2808
rect 3476 2796 3482 2848
rect 3697 2839 3755 2845
rect 3697 2805 3709 2839
rect 3743 2836 3755 2839
rect 4798 2836 4804 2848
rect 3743 2808 4804 2836
rect 3743 2805 3755 2808
rect 3697 2799 3755 2805
rect 4798 2796 4804 2808
rect 4856 2796 4862 2848
rect 4985 2839 5043 2845
rect 4985 2805 4997 2839
rect 5031 2836 5043 2839
rect 6914 2836 6920 2848
rect 5031 2808 6920 2836
rect 5031 2805 5043 2808
rect 4985 2799 5043 2805
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 7006 2796 7012 2848
rect 7064 2836 7070 2848
rect 7668 2836 7696 3012
rect 10042 3000 10048 3012
rect 10100 3000 10106 3052
rect 10137 3043 10195 3049
rect 10137 3009 10149 3043
rect 10183 3009 10195 3043
rect 10137 3003 10195 3009
rect 8846 2972 8852 2984
rect 8807 2944 8852 2972
rect 8846 2932 8852 2944
rect 8904 2932 8910 2984
rect 9030 2932 9036 2984
rect 9088 2972 9094 2984
rect 9125 2975 9183 2981
rect 9125 2972 9137 2975
rect 9088 2944 9137 2972
rect 9088 2932 9094 2944
rect 9125 2941 9137 2944
rect 9171 2972 9183 2975
rect 10152 2972 10180 3003
rect 10226 3000 10232 3052
rect 10284 3040 10290 3052
rect 10321 3043 10379 3049
rect 10321 3040 10333 3043
rect 10284 3012 10333 3040
rect 10284 3000 10290 3012
rect 10321 3009 10333 3012
rect 10367 3009 10379 3043
rect 10321 3003 10379 3009
rect 10502 3000 10508 3052
rect 10560 3040 10566 3052
rect 11330 3040 11336 3052
rect 10560 3012 11336 3040
rect 10560 3000 10566 3012
rect 11330 3000 11336 3012
rect 11388 3000 11394 3052
rect 11422 3000 11428 3052
rect 11480 3040 11486 3052
rect 11790 3049 11796 3052
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11480 3012 11529 3040
rect 11480 3000 11486 3012
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 11784 3003 11796 3049
rect 11848 3040 11854 3052
rect 11848 3012 11884 3040
rect 11790 3000 11796 3003
rect 11848 3000 11854 3012
rect 12986 3000 12992 3052
rect 13044 3040 13050 3052
rect 13357 3043 13415 3049
rect 13357 3040 13369 3043
rect 13044 3012 13369 3040
rect 13044 3000 13050 3012
rect 13357 3009 13369 3012
rect 13403 3009 13415 3043
rect 13538 3040 13544 3052
rect 13499 3012 13544 3040
rect 13357 3003 13415 3009
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 13633 3043 13691 3049
rect 13633 3009 13645 3043
rect 13679 3009 13691 3043
rect 13633 3003 13691 3009
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3040 13783 3043
rect 14090 3040 14096 3052
rect 13771 3012 14096 3040
rect 13771 3009 13783 3012
rect 13725 3003 13783 3009
rect 11054 2972 11060 2984
rect 9171 2944 9674 2972
rect 10152 2944 11060 2972
rect 9171 2941 9183 2944
rect 9125 2935 9183 2941
rect 9646 2904 9674 2944
rect 11054 2932 11060 2944
rect 11112 2932 11118 2984
rect 12710 2932 12716 2984
rect 12768 2972 12774 2984
rect 13648 2972 13676 3003
rect 14090 3000 14096 3012
rect 14148 3040 14154 3052
rect 16114 3040 16120 3052
rect 14148 3012 14964 3040
rect 16075 3012 16120 3040
rect 14148 3000 14154 3012
rect 14642 2972 14648 2984
rect 12768 2944 13676 2972
rect 14603 2944 14648 2972
rect 12768 2932 12774 2944
rect 14642 2932 14648 2944
rect 14700 2932 14706 2984
rect 14936 2981 14964 3012
rect 16114 3000 16120 3012
rect 16172 3000 16178 3052
rect 17954 3040 17960 3052
rect 17915 3012 17960 3040
rect 17954 3000 17960 3012
rect 18012 3000 18018 3052
rect 18141 3043 18199 3049
rect 18141 3009 18153 3043
rect 18187 3009 18199 3043
rect 18322 3040 18328 3052
rect 18283 3012 18328 3040
rect 18141 3003 18199 3009
rect 14921 2975 14979 2981
rect 14921 2941 14933 2975
rect 14967 2972 14979 2975
rect 15746 2972 15752 2984
rect 14967 2944 15752 2972
rect 14967 2941 14979 2944
rect 14921 2935 14979 2941
rect 15746 2932 15752 2944
rect 15804 2932 15810 2984
rect 16298 2932 16304 2984
rect 16356 2972 16362 2984
rect 16669 2975 16727 2981
rect 16669 2972 16681 2975
rect 16356 2944 16681 2972
rect 16356 2932 16362 2944
rect 16669 2941 16681 2944
rect 16715 2941 16727 2975
rect 16942 2972 16948 2984
rect 16855 2944 16948 2972
rect 16669 2935 16727 2941
rect 16942 2932 16948 2944
rect 17000 2972 17006 2984
rect 18156 2972 18184 3003
rect 18322 3000 18328 3012
rect 18380 3000 18386 3052
rect 19076 2972 19104 3080
rect 20622 3068 20628 3080
rect 20680 3108 20686 3120
rect 22005 3111 22063 3117
rect 22005 3108 22017 3111
rect 20680 3080 22017 3108
rect 20680 3068 20686 3080
rect 22005 3077 22017 3080
rect 22051 3077 22063 3111
rect 22005 3071 22063 3077
rect 22097 3111 22155 3117
rect 22097 3077 22109 3111
rect 22143 3077 22155 3111
rect 22097 3071 22155 3077
rect 19613 3043 19671 3049
rect 19613 3009 19625 3043
rect 19659 3009 19671 3043
rect 19613 3003 19671 3009
rect 19705 3043 19763 3049
rect 19705 3009 19717 3043
rect 19751 3040 19763 3043
rect 20070 3040 20076 3052
rect 19751 3012 20076 3040
rect 19751 3009 19763 3012
rect 19705 3003 19763 3009
rect 17000 2944 19104 2972
rect 19628 2972 19656 3003
rect 20070 3000 20076 3012
rect 20128 3000 20134 3052
rect 20254 3000 20260 3052
rect 20312 3040 20318 3052
rect 20349 3043 20407 3049
rect 20349 3040 20361 3043
rect 20312 3012 20361 3040
rect 20312 3000 20318 3012
rect 20349 3009 20361 3012
rect 20395 3009 20407 3043
rect 20349 3003 20407 3009
rect 20533 3043 20591 3049
rect 20533 3009 20545 3043
rect 20579 3040 20591 3043
rect 20990 3040 20996 3052
rect 20579 3012 20996 3040
rect 20579 3009 20591 3012
rect 20533 3003 20591 3009
rect 20364 2972 20392 3003
rect 20990 3000 20996 3012
rect 21048 3000 21054 3052
rect 21726 3000 21732 3052
rect 21784 3040 21790 3052
rect 21821 3043 21879 3049
rect 21821 3040 21833 3043
rect 21784 3012 21833 3040
rect 21784 3000 21790 3012
rect 21821 3009 21833 3012
rect 21867 3009 21879 3043
rect 21821 3003 21879 3009
rect 21910 2972 21916 2984
rect 19628 2944 21916 2972
rect 17000 2932 17006 2944
rect 21910 2932 21916 2944
rect 21968 2932 21974 2984
rect 22112 2972 22140 3071
rect 22646 3068 22652 3120
rect 22704 3108 22710 3120
rect 23474 3108 23480 3120
rect 22704 3080 23480 3108
rect 22704 3068 22710 3080
rect 23474 3068 23480 3080
rect 23532 3068 23538 3120
rect 23658 3068 23664 3120
rect 23716 3108 23722 3120
rect 27341 3111 27399 3117
rect 23716 3080 26464 3108
rect 23716 3068 23722 3080
rect 22186 3000 22192 3052
rect 22244 3040 22250 3052
rect 22244 3012 22289 3040
rect 22244 3000 22250 3012
rect 22922 3000 22928 3052
rect 22980 3040 22986 3052
rect 23017 3043 23075 3049
rect 23017 3040 23029 3043
rect 22980 3012 23029 3040
rect 22980 3000 22986 3012
rect 23017 3009 23029 3012
rect 23063 3009 23075 3043
rect 23017 3003 23075 3009
rect 24305 3043 24363 3049
rect 24305 3009 24317 3043
rect 24351 3040 24363 3043
rect 25958 3040 25964 3052
rect 24351 3012 25964 3040
rect 24351 3009 24363 3012
rect 24305 3003 24363 3009
rect 25958 3000 25964 3012
rect 26016 3000 26022 3052
rect 26436 3049 26464 3080
rect 27341 3077 27353 3111
rect 27387 3108 27399 3111
rect 27982 3108 27988 3120
rect 27387 3080 27988 3108
rect 27387 3077 27399 3080
rect 27341 3071 27399 3077
rect 27982 3068 27988 3080
rect 28040 3068 28046 3120
rect 28445 3111 28503 3117
rect 28445 3077 28457 3111
rect 28491 3108 28503 3111
rect 28534 3108 28540 3120
rect 28491 3080 28540 3108
rect 28491 3077 28503 3080
rect 28445 3071 28503 3077
rect 28534 3068 28540 3080
rect 28592 3068 28598 3120
rect 28810 3068 28816 3120
rect 28868 3108 28874 3120
rect 29273 3111 29331 3117
rect 29273 3108 29285 3111
rect 28868 3080 29285 3108
rect 28868 3068 28874 3080
rect 29273 3077 29285 3080
rect 29319 3077 29331 3111
rect 29273 3071 29331 3077
rect 30368 3111 30426 3117
rect 30368 3077 30380 3111
rect 30414 3108 30426 3111
rect 31018 3108 31024 3120
rect 30414 3080 31024 3108
rect 30414 3077 30426 3080
rect 30368 3071 30426 3077
rect 31018 3068 31024 3080
rect 31076 3068 31082 3120
rect 31726 3108 31754 3148
rect 33870 3136 33876 3188
rect 33928 3176 33934 3188
rect 33981 3179 34039 3185
rect 33981 3176 33993 3179
rect 33928 3148 33993 3176
rect 33928 3136 33934 3148
rect 33980 3145 33993 3148
rect 34027 3145 34039 3179
rect 34146 3176 34152 3188
rect 34107 3148 34152 3176
rect 33980 3139 34039 3145
rect 33781 3111 33839 3117
rect 33781 3108 33793 3111
rect 31726 3080 33793 3108
rect 33781 3077 33793 3080
rect 33827 3077 33839 3111
rect 33980 3108 34008 3139
rect 34146 3136 34152 3148
rect 34204 3136 34210 3188
rect 35545 3179 35603 3185
rect 35545 3176 35557 3179
rect 35176 3148 35557 3176
rect 35176 3108 35204 3148
rect 35545 3145 35557 3148
rect 35591 3176 35603 3179
rect 35713 3179 35771 3185
rect 35591 3148 35664 3176
rect 35591 3145 35603 3148
rect 35545 3139 35603 3145
rect 35342 3108 35348 3120
rect 33980 3080 35204 3108
rect 35303 3080 35348 3108
rect 33781 3071 33839 3077
rect 35342 3068 35348 3080
rect 35400 3068 35406 3120
rect 26421 3043 26479 3049
rect 26421 3009 26433 3043
rect 26467 3009 26479 3043
rect 26421 3003 26479 3009
rect 26878 3000 26884 3052
rect 26936 3040 26942 3052
rect 29638 3040 29644 3052
rect 26936 3012 29644 3040
rect 26936 3000 26942 3012
rect 29638 3000 29644 3012
rect 29696 3000 29702 3052
rect 29730 3000 29736 3052
rect 29788 3040 29794 3052
rect 30101 3043 30159 3049
rect 30101 3040 30113 3043
rect 29788 3012 30113 3040
rect 29788 3000 29794 3012
rect 30101 3009 30113 3012
rect 30147 3009 30159 3043
rect 30101 3003 30159 3009
rect 30834 3000 30840 3052
rect 30892 3040 30898 3052
rect 30892 3012 31248 3040
rect 30892 3000 30898 3012
rect 22112 2944 22232 2972
rect 10226 2904 10232 2916
rect 9646 2876 10232 2904
rect 10226 2864 10232 2876
rect 10284 2904 10290 2916
rect 10594 2904 10600 2916
rect 10284 2876 10600 2904
rect 10284 2864 10290 2876
rect 10594 2864 10600 2876
rect 10652 2864 10658 2916
rect 13722 2904 13728 2916
rect 12820 2876 13728 2904
rect 7064 2808 7696 2836
rect 7064 2796 7070 2808
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 9122 2836 9128 2848
rect 8352 2808 9128 2836
rect 8352 2796 8358 2808
rect 9122 2796 9128 2808
rect 9180 2796 9186 2848
rect 9306 2796 9312 2848
rect 9364 2836 9370 2848
rect 9490 2836 9496 2848
rect 9364 2808 9496 2836
rect 9364 2796 9370 2808
rect 9490 2796 9496 2808
rect 9548 2796 9554 2848
rect 10134 2796 10140 2848
rect 10192 2836 10198 2848
rect 10689 2839 10747 2845
rect 10689 2836 10701 2839
rect 10192 2808 10701 2836
rect 10192 2796 10198 2808
rect 10689 2805 10701 2808
rect 10735 2805 10747 2839
rect 10689 2799 10747 2805
rect 10778 2796 10784 2848
rect 10836 2836 10842 2848
rect 12820 2836 12848 2876
rect 13722 2864 13728 2876
rect 13780 2864 13786 2916
rect 21266 2904 21272 2916
rect 21100 2876 21272 2904
rect 21100 2848 21128 2876
rect 21266 2864 21272 2876
rect 21324 2864 21330 2916
rect 10836 2808 12848 2836
rect 12897 2839 12955 2845
rect 10836 2796 10842 2808
rect 12897 2805 12909 2839
rect 12943 2836 12955 2839
rect 12986 2836 12992 2848
rect 12943 2808 12992 2836
rect 12943 2805 12955 2808
rect 12897 2799 12955 2805
rect 12986 2796 12992 2808
rect 13044 2796 13050 2848
rect 13906 2836 13912 2848
rect 13867 2808 13912 2836
rect 13906 2796 13912 2808
rect 13964 2796 13970 2848
rect 14550 2796 14556 2848
rect 14608 2836 14614 2848
rect 16666 2836 16672 2848
rect 14608 2808 16672 2836
rect 14608 2796 14614 2808
rect 16666 2796 16672 2808
rect 16724 2836 16730 2848
rect 18046 2836 18052 2848
rect 16724 2808 18052 2836
rect 16724 2796 16730 2808
rect 18046 2796 18052 2808
rect 18104 2796 18110 2848
rect 21082 2796 21088 2848
rect 21140 2796 21146 2848
rect 21174 2796 21180 2848
rect 21232 2836 21238 2848
rect 22094 2836 22100 2848
rect 21232 2808 22100 2836
rect 21232 2796 21238 2808
rect 22094 2796 22100 2808
rect 22152 2796 22158 2848
rect 22204 2836 22232 2944
rect 22278 2932 22284 2984
rect 22336 2972 22342 2984
rect 22833 2975 22891 2981
rect 22833 2972 22845 2975
rect 22336 2944 22845 2972
rect 22336 2932 22342 2944
rect 22833 2941 22845 2944
rect 22879 2972 22891 2975
rect 24121 2975 24179 2981
rect 24121 2972 24133 2975
rect 22879 2944 24133 2972
rect 22879 2941 22891 2944
rect 22833 2935 22891 2941
rect 24121 2941 24133 2944
rect 24167 2972 24179 2975
rect 24394 2972 24400 2984
rect 24167 2944 24400 2972
rect 24167 2941 24179 2944
rect 24121 2935 24179 2941
rect 24394 2932 24400 2944
rect 24452 2932 24458 2984
rect 25130 2932 25136 2984
rect 25188 2972 25194 2984
rect 25317 2975 25375 2981
rect 25317 2972 25329 2975
rect 25188 2944 25329 2972
rect 25188 2932 25194 2944
rect 25317 2941 25329 2944
rect 25363 2941 25375 2975
rect 29178 2972 29184 2984
rect 25317 2935 25375 2941
rect 25424 2944 29184 2972
rect 22370 2904 22376 2916
rect 22331 2876 22376 2904
rect 22370 2864 22376 2876
rect 22428 2864 22434 2916
rect 22922 2864 22928 2916
rect 22980 2904 22986 2916
rect 23290 2904 23296 2916
rect 22980 2876 23296 2904
rect 22980 2864 22986 2876
rect 23290 2864 23296 2876
rect 23348 2864 23354 2916
rect 23842 2864 23848 2916
rect 23900 2904 23906 2916
rect 25424 2904 25452 2944
rect 29178 2932 29184 2944
rect 29236 2932 29242 2984
rect 31220 2972 31248 3012
rect 31294 3000 31300 3052
rect 31352 3040 31358 3052
rect 31754 3040 31760 3052
rect 31352 3012 31760 3040
rect 31352 3000 31358 3012
rect 31754 3000 31760 3012
rect 31812 3000 31818 3052
rect 32125 3043 32183 3049
rect 32125 3009 32137 3043
rect 32171 3040 32183 3043
rect 32858 3040 32864 3052
rect 32171 3012 32720 3040
rect 32819 3012 32864 3040
rect 32171 3009 32183 3012
rect 32125 3003 32183 3009
rect 32306 2972 32312 2984
rect 31220 2944 32312 2972
rect 32306 2932 32312 2944
rect 32364 2932 32370 2984
rect 32692 2972 32720 3012
rect 32858 3000 32864 3012
rect 32916 3000 32922 3052
rect 34609 3043 34667 3049
rect 34609 3009 34621 3043
rect 34655 3040 34667 3043
rect 34655 3012 35388 3040
rect 34655 3009 34667 3012
rect 34609 3003 34667 3009
rect 33318 2972 33324 2984
rect 32692 2944 33324 2972
rect 33318 2932 33324 2944
rect 33376 2932 33382 2984
rect 23900 2876 25452 2904
rect 23900 2864 23906 2876
rect 25498 2864 25504 2916
rect 25556 2904 25562 2916
rect 25685 2907 25743 2913
rect 25685 2904 25697 2907
rect 25556 2876 25697 2904
rect 25556 2864 25562 2876
rect 25685 2873 25697 2876
rect 25731 2904 25743 2907
rect 26050 2904 26056 2916
rect 25731 2876 26056 2904
rect 25731 2873 25743 2876
rect 25685 2867 25743 2873
rect 26050 2864 26056 2876
rect 26108 2864 26114 2916
rect 27709 2907 27767 2913
rect 27709 2873 27721 2907
rect 27755 2904 27767 2907
rect 28074 2904 28080 2916
rect 27755 2876 28080 2904
rect 27755 2873 27767 2876
rect 27709 2867 27767 2873
rect 28074 2864 28080 2876
rect 28132 2864 28138 2916
rect 28534 2864 28540 2916
rect 28592 2904 28598 2916
rect 33045 2907 33103 2913
rect 33045 2904 33057 2907
rect 28592 2876 29776 2904
rect 28592 2864 28598 2876
rect 23106 2836 23112 2848
rect 22204 2808 23112 2836
rect 23106 2796 23112 2808
rect 23164 2796 23170 2848
rect 23201 2839 23259 2845
rect 23201 2805 23213 2839
rect 23247 2836 23259 2839
rect 24302 2836 24308 2848
rect 23247 2808 24308 2836
rect 23247 2805 23259 2808
rect 23201 2799 23259 2805
rect 24302 2796 24308 2808
rect 24360 2796 24366 2848
rect 24762 2796 24768 2848
rect 24820 2836 24826 2848
rect 26237 2839 26295 2845
rect 26237 2836 26249 2839
rect 24820 2808 26249 2836
rect 24820 2796 24826 2808
rect 26237 2805 26249 2808
rect 26283 2805 26295 2839
rect 28626 2836 28632 2848
rect 28587 2808 28632 2836
rect 26237 2799 26295 2805
rect 28626 2796 28632 2808
rect 28684 2796 28690 2848
rect 28718 2796 28724 2848
rect 28776 2836 28782 2848
rect 28813 2839 28871 2845
rect 28813 2836 28825 2839
rect 28776 2808 28825 2836
rect 28776 2796 28782 2808
rect 28813 2805 28825 2808
rect 28859 2805 28871 2839
rect 28813 2799 28871 2805
rect 28902 2796 28908 2848
rect 28960 2836 28966 2848
rect 29454 2836 29460 2848
rect 28960 2808 29460 2836
rect 28960 2796 28966 2808
rect 29454 2796 29460 2808
rect 29512 2796 29518 2848
rect 29748 2836 29776 2876
rect 32232 2876 33057 2904
rect 30742 2836 30748 2848
rect 29748 2808 30748 2836
rect 30742 2796 30748 2808
rect 30800 2796 30806 2848
rect 31570 2796 31576 2848
rect 31628 2836 31634 2848
rect 32232 2836 32260 2876
rect 33045 2873 33057 2876
rect 33091 2873 33103 2907
rect 33045 2867 33103 2873
rect 33778 2864 33784 2916
rect 33836 2904 33842 2916
rect 34793 2907 34851 2913
rect 34793 2904 34805 2907
rect 33836 2876 34805 2904
rect 33836 2864 33842 2876
rect 34793 2873 34805 2876
rect 34839 2873 34851 2907
rect 35360 2904 35388 3012
rect 35636 2972 35664 3148
rect 35713 3145 35725 3179
rect 35759 3176 35771 3179
rect 36262 3176 36268 3188
rect 35759 3148 36268 3176
rect 35759 3145 35771 3148
rect 35713 3139 35771 3145
rect 36262 3136 36268 3148
rect 36320 3136 36326 3188
rect 36541 3179 36599 3185
rect 36541 3145 36553 3179
rect 36587 3176 36599 3179
rect 37090 3176 37096 3188
rect 36587 3148 37096 3176
rect 36587 3145 36599 3148
rect 36541 3139 36599 3145
rect 37090 3136 37096 3148
rect 37148 3136 37154 3188
rect 35802 3068 35808 3120
rect 35860 3108 35866 3120
rect 36173 3111 36231 3117
rect 36173 3108 36185 3111
rect 35860 3080 36185 3108
rect 35860 3068 35866 3080
rect 36173 3077 36185 3080
rect 36219 3077 36231 3111
rect 36354 3108 36360 3120
rect 36412 3117 36418 3120
rect 36412 3111 36431 3117
rect 36173 3071 36231 3077
rect 36280 3080 36360 3108
rect 36280 2972 36308 3080
rect 36354 3068 36360 3080
rect 36419 3108 36431 3111
rect 36419 3080 36505 3108
rect 36419 3077 36431 3080
rect 36412 3071 36431 3077
rect 36412 3068 36418 3071
rect 37277 3043 37335 3049
rect 37277 3009 37289 3043
rect 37323 3040 37335 3043
rect 37366 3040 37372 3052
rect 37323 3012 37372 3040
rect 37323 3009 37335 3012
rect 37277 3003 37335 3009
rect 37366 3000 37372 3012
rect 37424 3000 37430 3052
rect 35636 2944 36308 2972
rect 36170 2904 36176 2916
rect 35360 2876 36176 2904
rect 34793 2867 34851 2873
rect 36170 2864 36176 2876
rect 36228 2864 36234 2916
rect 31628 2808 32260 2836
rect 31628 2796 31634 2808
rect 32306 2796 32312 2848
rect 32364 2836 32370 2848
rect 33965 2839 34023 2845
rect 32364 2808 32409 2836
rect 32364 2796 32370 2808
rect 33965 2805 33977 2839
rect 34011 2836 34023 2839
rect 35529 2839 35587 2845
rect 35529 2836 35541 2839
rect 34011 2808 35541 2836
rect 34011 2805 34023 2808
rect 33965 2799 34023 2805
rect 35529 2805 35541 2808
rect 35575 2836 35587 2839
rect 36357 2839 36415 2845
rect 36357 2836 36369 2839
rect 35575 2808 36369 2836
rect 35575 2805 35587 2808
rect 35529 2799 35587 2805
rect 36357 2805 36369 2808
rect 36403 2836 36415 2839
rect 36446 2836 36452 2848
rect 36403 2808 36452 2836
rect 36403 2805 36415 2808
rect 36357 2799 36415 2805
rect 36446 2796 36452 2808
rect 36504 2796 36510 2848
rect 36814 2796 36820 2848
rect 36872 2836 36878 2848
rect 37461 2839 37519 2845
rect 37461 2836 37473 2839
rect 36872 2808 37473 2836
rect 36872 2796 36878 2808
rect 37461 2805 37473 2808
rect 37507 2805 37519 2839
rect 37461 2799 37519 2805
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 3234 2632 3240 2644
rect 2608 2604 3240 2632
rect 566 2388 572 2440
rect 624 2428 630 2440
rect 2608 2437 2636 2604
rect 3234 2592 3240 2604
rect 3292 2592 3298 2644
rect 3326 2592 3332 2644
rect 3384 2632 3390 2644
rect 5350 2632 5356 2644
rect 3384 2604 5356 2632
rect 3384 2592 3390 2604
rect 5350 2592 5356 2604
rect 5408 2592 5414 2644
rect 6454 2592 6460 2644
rect 6512 2632 6518 2644
rect 6733 2635 6791 2641
rect 6733 2632 6745 2635
rect 6512 2604 6745 2632
rect 6512 2592 6518 2604
rect 6733 2601 6745 2604
rect 6779 2601 6791 2635
rect 7374 2632 7380 2644
rect 7335 2604 7380 2632
rect 6733 2595 6791 2601
rect 7374 2592 7380 2604
rect 7432 2592 7438 2644
rect 8110 2592 8116 2644
rect 8168 2632 8174 2644
rect 9214 2632 9220 2644
rect 8168 2604 9220 2632
rect 8168 2592 8174 2604
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 10318 2632 10324 2644
rect 10279 2604 10324 2632
rect 10318 2592 10324 2604
rect 10376 2592 10382 2644
rect 10781 2635 10839 2641
rect 10781 2601 10793 2635
rect 10827 2632 10839 2635
rect 11238 2632 11244 2644
rect 10827 2604 11244 2632
rect 10827 2601 10839 2604
rect 10781 2595 10839 2601
rect 11238 2592 11244 2604
rect 11296 2592 11302 2644
rect 11790 2592 11796 2644
rect 11848 2632 11854 2644
rect 11885 2635 11943 2641
rect 11885 2632 11897 2635
rect 11848 2604 11897 2632
rect 11848 2592 11854 2604
rect 11885 2601 11897 2604
rect 11931 2601 11943 2635
rect 11885 2595 11943 2601
rect 15838 2592 15844 2644
rect 15896 2632 15902 2644
rect 15933 2635 15991 2641
rect 15933 2632 15945 2635
rect 15896 2604 15945 2632
rect 15896 2592 15902 2604
rect 15933 2601 15945 2604
rect 15979 2601 15991 2635
rect 15933 2595 15991 2601
rect 16574 2592 16580 2644
rect 16632 2632 16638 2644
rect 19429 2635 19487 2641
rect 19429 2632 19441 2635
rect 16632 2604 19441 2632
rect 16632 2592 16638 2604
rect 19429 2601 19441 2604
rect 19475 2601 19487 2635
rect 19429 2595 19487 2601
rect 21269 2635 21327 2641
rect 21269 2601 21281 2635
rect 21315 2632 21327 2635
rect 21542 2632 21548 2644
rect 21315 2604 21548 2632
rect 21315 2601 21327 2604
rect 21269 2595 21327 2601
rect 21542 2592 21548 2604
rect 21600 2592 21606 2644
rect 22741 2635 22799 2641
rect 22741 2601 22753 2635
rect 22787 2632 22799 2635
rect 23014 2632 23020 2644
rect 22787 2604 23020 2632
rect 22787 2601 22799 2604
rect 22741 2595 22799 2601
rect 23014 2592 23020 2604
rect 23072 2592 23078 2644
rect 24946 2592 24952 2644
rect 25004 2632 25010 2644
rect 26237 2635 26295 2641
rect 26237 2632 26249 2635
rect 25004 2604 26249 2632
rect 25004 2592 25010 2604
rect 26237 2601 26249 2604
rect 26283 2601 26295 2635
rect 26237 2595 26295 2601
rect 27709 2635 27767 2641
rect 27709 2601 27721 2635
rect 27755 2632 27767 2635
rect 27890 2632 27896 2644
rect 27755 2604 27896 2632
rect 27755 2601 27767 2604
rect 27709 2595 27767 2601
rect 27890 2592 27896 2604
rect 27948 2592 27954 2644
rect 28537 2635 28595 2641
rect 28537 2601 28549 2635
rect 28583 2632 28595 2635
rect 28626 2632 28632 2644
rect 28583 2604 28632 2632
rect 28583 2601 28595 2604
rect 28537 2595 28595 2601
rect 28626 2592 28632 2604
rect 28684 2632 28690 2644
rect 28902 2632 28908 2644
rect 28684 2604 28908 2632
rect 28684 2592 28690 2604
rect 28902 2592 28908 2604
rect 28960 2592 28966 2644
rect 30742 2592 30748 2644
rect 30800 2632 30806 2644
rect 31205 2635 31263 2641
rect 31205 2632 31217 2635
rect 30800 2604 31217 2632
rect 30800 2592 30806 2604
rect 31205 2601 31217 2604
rect 31251 2601 31263 2635
rect 31205 2595 31263 2601
rect 6086 2524 6092 2576
rect 6144 2564 6150 2576
rect 6914 2564 6920 2576
rect 6144 2536 6920 2564
rect 6144 2524 6150 2536
rect 6914 2524 6920 2536
rect 6972 2524 6978 2576
rect 8018 2524 8024 2576
rect 8076 2564 8082 2576
rect 13262 2564 13268 2576
rect 8076 2536 8984 2564
rect 8076 2524 8082 2536
rect 3237 2499 3295 2505
rect 3237 2465 3249 2499
rect 3283 2496 3295 2499
rect 3878 2496 3884 2508
rect 3283 2468 3884 2496
rect 3283 2465 3295 2468
rect 3237 2459 3295 2465
rect 3878 2456 3884 2468
rect 3936 2456 3942 2508
rect 3970 2456 3976 2508
rect 4028 2496 4034 2508
rect 7374 2496 7380 2508
rect 4028 2468 7380 2496
rect 4028 2456 4034 2468
rect 7374 2456 7380 2468
rect 7432 2456 7438 2508
rect 8389 2499 8447 2505
rect 8389 2496 8401 2499
rect 7576 2468 8401 2496
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 624 2400 1409 2428
rect 624 2388 630 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2397 2651 2431
rect 2593 2391 2651 2397
rect 3602 2388 3608 2440
rect 3660 2428 3666 2440
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3660 2400 3801 2428
rect 3660 2388 3666 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 4614 2388 4620 2440
rect 4672 2428 4678 2440
rect 4709 2431 4767 2437
rect 4709 2428 4721 2431
rect 4672 2400 4721 2428
rect 4672 2388 4678 2400
rect 4709 2397 4721 2400
rect 4755 2397 4767 2431
rect 4982 2428 4988 2440
rect 4943 2400 4988 2428
rect 4709 2391 4767 2397
rect 4982 2388 4988 2400
rect 5040 2388 5046 2440
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2428 6975 2431
rect 7466 2428 7472 2440
rect 6963 2400 7472 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 7466 2388 7472 2400
rect 7524 2388 7530 2440
rect 7576 2437 7604 2468
rect 8389 2465 8401 2468
rect 8435 2465 8447 2499
rect 8389 2459 8447 2465
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2397 7619 2431
rect 8110 2428 8116 2440
rect 8071 2400 8116 2428
rect 7561 2391 7619 2397
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 8202 2388 8208 2440
rect 8260 2428 8266 2440
rect 8956 2437 8984 2536
rect 10980 2536 13268 2564
rect 9214 2456 9220 2508
rect 9272 2496 9278 2508
rect 9953 2499 10011 2505
rect 9953 2496 9965 2499
rect 9272 2468 9965 2496
rect 9272 2456 9278 2468
rect 9953 2465 9965 2468
rect 9999 2465 10011 2499
rect 9953 2459 10011 2465
rect 8941 2431 8999 2437
rect 8260 2400 8305 2428
rect 8260 2388 8266 2400
rect 8941 2397 8953 2431
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9309 2431 9367 2437
rect 9088 2400 9168 2428
rect 9088 2388 9094 2400
rect 7834 2360 7840 2372
rect 2424 2332 7840 2360
rect 1578 2292 1584 2304
rect 1539 2264 1584 2292
rect 1578 2252 1584 2264
rect 1636 2252 1642 2304
rect 2424 2301 2452 2332
rect 7834 2320 7840 2332
rect 7892 2320 7898 2372
rect 9140 2369 9168 2400
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 9398 2428 9404 2440
rect 9355 2400 9404 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 9398 2388 9404 2400
rect 9456 2388 9462 2440
rect 10134 2428 10140 2440
rect 10095 2400 10140 2428
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 10980 2437 11008 2536
rect 13262 2524 13268 2536
rect 13320 2524 13326 2576
rect 16298 2564 16304 2576
rect 14108 2536 16304 2564
rect 12618 2496 12624 2508
rect 12579 2468 12624 2496
rect 12618 2456 12624 2468
rect 12676 2456 12682 2508
rect 14108 2505 14136 2536
rect 16298 2524 16304 2536
rect 16356 2524 16362 2576
rect 17313 2567 17371 2573
rect 17313 2533 17325 2567
rect 17359 2533 17371 2567
rect 17313 2527 17371 2533
rect 14093 2499 14151 2505
rect 14093 2465 14105 2499
rect 14139 2465 14151 2499
rect 14093 2459 14151 2465
rect 14369 2499 14427 2505
rect 14369 2465 14381 2499
rect 14415 2496 14427 2499
rect 14826 2496 14832 2508
rect 14415 2468 14832 2496
rect 14415 2465 14427 2468
rect 14369 2459 14427 2465
rect 10965 2431 11023 2437
rect 10965 2397 10977 2431
rect 11011 2397 11023 2431
rect 10965 2391 11023 2397
rect 12069 2431 12127 2437
rect 12069 2397 12081 2431
rect 12115 2428 12127 2431
rect 12805 2431 12863 2437
rect 12115 2400 12434 2428
rect 12115 2397 12127 2400
rect 12069 2391 12127 2397
rect 9125 2363 9183 2369
rect 9125 2329 9137 2363
rect 9171 2329 9183 2363
rect 9125 2323 9183 2329
rect 9217 2363 9275 2369
rect 9217 2329 9229 2363
rect 9263 2329 9275 2363
rect 12406 2360 12434 2400
rect 12805 2397 12817 2431
rect 12851 2428 12863 2431
rect 13906 2428 13912 2440
rect 12851 2400 13912 2428
rect 12851 2397 12863 2400
rect 12805 2391 12863 2397
rect 13906 2388 13912 2400
rect 13964 2388 13970 2440
rect 12989 2363 13047 2369
rect 12989 2360 13001 2363
rect 12406 2332 13001 2360
rect 9217 2323 9275 2329
rect 12989 2329 13001 2332
rect 13035 2329 13047 2363
rect 12989 2323 13047 2329
rect 2409 2295 2467 2301
rect 2409 2261 2421 2295
rect 2455 2261 2467 2295
rect 2409 2255 2467 2261
rect 3142 2252 3148 2304
rect 3200 2292 3206 2304
rect 3973 2295 4031 2301
rect 3973 2292 3985 2295
rect 3200 2264 3985 2292
rect 3200 2252 3206 2264
rect 3973 2261 3985 2264
rect 4019 2261 4031 2295
rect 3973 2255 4031 2261
rect 4706 2252 4712 2304
rect 4764 2292 4770 2304
rect 7282 2292 7288 2304
rect 4764 2264 7288 2292
rect 4764 2252 4770 2264
rect 7282 2252 7288 2264
rect 7340 2252 7346 2304
rect 7374 2252 7380 2304
rect 7432 2292 7438 2304
rect 9232 2292 9260 2323
rect 7432 2264 9260 2292
rect 7432 2252 7438 2264
rect 9306 2252 9312 2304
rect 9364 2292 9370 2304
rect 9493 2295 9551 2301
rect 9493 2292 9505 2295
rect 9364 2264 9505 2292
rect 9364 2252 9370 2264
rect 9493 2261 9505 2264
rect 9539 2261 9551 2295
rect 9493 2255 9551 2261
rect 12342 2252 12348 2304
rect 12400 2292 12406 2304
rect 14108 2292 14136 2459
rect 14826 2456 14832 2468
rect 14884 2496 14890 2508
rect 17328 2496 17356 2527
rect 17402 2524 17408 2576
rect 17460 2564 17466 2576
rect 20165 2567 20223 2573
rect 20165 2564 20177 2567
rect 17460 2536 20177 2564
rect 17460 2524 17466 2536
rect 20165 2533 20177 2536
rect 20211 2533 20223 2567
rect 20165 2527 20223 2533
rect 23753 2567 23811 2573
rect 23753 2533 23765 2567
rect 23799 2564 23811 2567
rect 24854 2564 24860 2576
rect 23799 2536 24860 2564
rect 23799 2533 23811 2536
rect 23753 2527 23811 2533
rect 24854 2524 24860 2536
rect 24912 2524 24918 2576
rect 25590 2524 25596 2576
rect 25648 2564 25654 2576
rect 27157 2567 27215 2573
rect 27157 2564 27169 2567
rect 25648 2536 27169 2564
rect 25648 2524 25654 2536
rect 27157 2533 27169 2536
rect 27203 2533 27215 2567
rect 27157 2527 27215 2533
rect 27798 2524 27804 2576
rect 27856 2564 27862 2576
rect 30469 2567 30527 2573
rect 30469 2564 30481 2567
rect 27856 2536 30481 2564
rect 27856 2524 27862 2536
rect 30469 2533 30481 2536
rect 30515 2533 30527 2567
rect 30469 2527 30527 2533
rect 32306 2524 32312 2576
rect 32364 2564 32370 2576
rect 33781 2567 33839 2573
rect 33781 2564 33793 2567
rect 32364 2536 33793 2564
rect 32364 2524 32370 2536
rect 33781 2533 33793 2536
rect 33827 2533 33839 2567
rect 33781 2527 33839 2533
rect 34606 2524 34612 2576
rect 34664 2564 34670 2576
rect 35621 2567 35679 2573
rect 35621 2564 35633 2567
rect 34664 2536 35633 2564
rect 34664 2524 34670 2536
rect 35621 2533 35633 2536
rect 35667 2533 35679 2567
rect 35621 2527 35679 2533
rect 36078 2524 36084 2576
rect 36136 2564 36142 2576
rect 37461 2567 37519 2573
rect 37461 2564 37473 2567
rect 36136 2536 37473 2564
rect 36136 2524 36142 2536
rect 37461 2533 37473 2536
rect 37507 2533 37519 2567
rect 37461 2527 37519 2533
rect 17586 2496 17592 2508
rect 14884 2468 15608 2496
rect 17328 2468 17592 2496
rect 14884 2456 14890 2468
rect 15580 2437 15608 2468
rect 17586 2456 17592 2468
rect 17644 2456 17650 2508
rect 18322 2496 18328 2508
rect 17696 2468 18328 2496
rect 15381 2431 15439 2437
rect 15381 2397 15393 2431
rect 15427 2397 15439 2431
rect 15381 2391 15439 2397
rect 15565 2431 15623 2437
rect 15565 2397 15577 2431
rect 15611 2397 15623 2431
rect 15746 2428 15752 2440
rect 15707 2400 15752 2428
rect 15565 2391 15623 2397
rect 12400 2264 14136 2292
rect 15396 2292 15424 2391
rect 15746 2388 15752 2400
rect 15804 2388 15810 2440
rect 16758 2428 16764 2440
rect 16719 2400 16764 2428
rect 16758 2388 16764 2400
rect 16816 2388 16822 2440
rect 16942 2428 16948 2440
rect 16903 2400 16948 2428
rect 16942 2388 16948 2400
rect 17000 2388 17006 2440
rect 17126 2388 17132 2440
rect 17184 2437 17190 2440
rect 17184 2431 17233 2437
rect 17184 2397 17187 2431
rect 17221 2428 17233 2431
rect 17696 2428 17724 2468
rect 18322 2456 18328 2468
rect 18380 2456 18386 2508
rect 19334 2496 19340 2508
rect 18524 2468 19340 2496
rect 17862 2428 17868 2440
rect 17221 2400 17724 2428
rect 17823 2400 17868 2428
rect 17221 2397 17233 2400
rect 17184 2391 17233 2397
rect 17184 2388 17190 2391
rect 17862 2388 17868 2400
rect 17920 2388 17926 2440
rect 17957 2431 18015 2437
rect 17957 2397 17969 2431
rect 18003 2397 18015 2431
rect 17957 2391 18015 2397
rect 15654 2360 15660 2372
rect 15615 2332 15660 2360
rect 15654 2320 15660 2332
rect 15712 2320 15718 2372
rect 16022 2320 16028 2372
rect 16080 2360 16086 2372
rect 17034 2360 17040 2372
rect 16080 2332 16896 2360
rect 16995 2332 17040 2360
rect 16080 2320 16086 2332
rect 16482 2292 16488 2304
rect 15396 2264 16488 2292
rect 12400 2252 12406 2264
rect 16482 2252 16488 2264
rect 16540 2252 16546 2304
rect 16868 2292 16896 2332
rect 17034 2320 17040 2332
rect 17092 2320 17098 2372
rect 17586 2320 17592 2372
rect 17644 2360 17650 2372
rect 17975 2360 18003 2391
rect 18046 2388 18052 2440
rect 18104 2428 18110 2440
rect 18524 2428 18552 2468
rect 19334 2456 19340 2468
rect 19392 2496 19398 2508
rect 20901 2499 20959 2505
rect 20901 2496 20913 2499
rect 19392 2468 20913 2496
rect 19392 2456 19398 2468
rect 20901 2465 20913 2468
rect 20947 2465 20959 2499
rect 22370 2496 22376 2508
rect 22331 2468 22376 2496
rect 20901 2459 20959 2465
rect 22370 2456 22376 2468
rect 22428 2456 22434 2508
rect 24210 2456 24216 2508
rect 24268 2496 24274 2508
rect 25777 2499 25835 2505
rect 24268 2468 25636 2496
rect 24268 2456 24274 2468
rect 18104 2400 18552 2428
rect 18104 2388 18110 2400
rect 18598 2388 18604 2440
rect 18656 2428 18662 2440
rect 19245 2431 19303 2437
rect 19245 2428 19257 2431
rect 18656 2400 19257 2428
rect 18656 2388 18662 2400
rect 19245 2397 19257 2400
rect 19291 2397 19303 2431
rect 19245 2391 19303 2397
rect 19981 2431 20039 2437
rect 19981 2397 19993 2431
rect 20027 2428 20039 2431
rect 20806 2428 20812 2440
rect 20027 2400 20812 2428
rect 20027 2397 20039 2400
rect 19981 2391 20039 2397
rect 20806 2388 20812 2400
rect 20864 2388 20870 2440
rect 21082 2428 21088 2440
rect 21043 2400 21088 2428
rect 21082 2388 21088 2400
rect 21140 2388 21146 2440
rect 22554 2428 22560 2440
rect 22515 2400 22560 2428
rect 22554 2388 22560 2400
rect 22612 2388 22618 2440
rect 23569 2431 23627 2437
rect 23569 2397 23581 2431
rect 23615 2428 23627 2431
rect 24026 2428 24032 2440
rect 23615 2400 24032 2428
rect 23615 2397 23627 2400
rect 23569 2391 23627 2397
rect 24026 2388 24032 2400
rect 24084 2388 24090 2440
rect 24397 2431 24455 2437
rect 24397 2397 24409 2431
rect 24443 2428 24455 2431
rect 25222 2428 25228 2440
rect 24443 2400 25228 2428
rect 24443 2397 24455 2400
rect 24397 2391 24455 2397
rect 25222 2388 25228 2400
rect 25280 2388 25286 2440
rect 25498 2428 25504 2440
rect 25459 2400 25504 2428
rect 25498 2388 25504 2400
rect 25556 2388 25562 2440
rect 25608 2437 25636 2468
rect 25777 2465 25789 2499
rect 25823 2496 25835 2499
rect 29270 2496 29276 2508
rect 25823 2468 29276 2496
rect 25823 2465 25835 2468
rect 25777 2459 25835 2465
rect 29270 2456 29276 2468
rect 29328 2456 29334 2508
rect 29914 2456 29920 2508
rect 29972 2496 29978 2508
rect 29972 2468 31064 2496
rect 29972 2456 29978 2468
rect 25593 2431 25651 2437
rect 25593 2397 25605 2431
rect 25639 2397 25651 2431
rect 25593 2391 25651 2397
rect 26234 2388 26240 2440
rect 26292 2428 26298 2440
rect 26421 2431 26479 2437
rect 26421 2428 26433 2431
rect 26292 2400 26433 2428
rect 26292 2388 26298 2400
rect 26421 2397 26433 2400
rect 26467 2397 26479 2431
rect 26421 2391 26479 2397
rect 26510 2388 26516 2440
rect 26568 2428 26574 2440
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26568 2400 26985 2428
rect 26568 2388 26574 2400
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 27893 2431 27951 2437
rect 27893 2397 27905 2431
rect 27939 2397 27951 2431
rect 27893 2391 27951 2397
rect 17644 2332 18003 2360
rect 17644 2320 17650 2332
rect 24302 2320 24308 2372
rect 24360 2360 24366 2372
rect 27908 2360 27936 2391
rect 28074 2388 28080 2440
rect 28132 2428 28138 2440
rect 29546 2428 29552 2440
rect 28132 2400 28580 2428
rect 29507 2400 29552 2428
rect 28132 2388 28138 2400
rect 28350 2360 28356 2372
rect 24360 2332 27936 2360
rect 28311 2332 28356 2360
rect 24360 2320 24366 2332
rect 28350 2320 28356 2332
rect 28408 2320 28414 2372
rect 28552 2369 28580 2400
rect 29546 2388 29552 2400
rect 29604 2388 29610 2440
rect 30285 2431 30343 2437
rect 30285 2397 30297 2431
rect 30331 2428 30343 2431
rect 30374 2428 30380 2440
rect 30331 2400 30380 2428
rect 30331 2397 30343 2400
rect 30285 2391 30343 2397
rect 30374 2388 30380 2400
rect 30432 2388 30438 2440
rect 31036 2437 31064 2468
rect 35526 2456 35532 2508
rect 35584 2496 35590 2508
rect 35584 2468 36216 2496
rect 35584 2456 35590 2468
rect 31021 2431 31079 2437
rect 31021 2397 31033 2431
rect 31067 2397 31079 2431
rect 31021 2391 31079 2397
rect 32030 2388 32036 2440
rect 32088 2428 32094 2440
rect 32125 2431 32183 2437
rect 32125 2428 32137 2431
rect 32088 2400 32137 2428
rect 32088 2388 32094 2400
rect 32125 2397 32137 2400
rect 32171 2397 32183 2431
rect 32125 2391 32183 2397
rect 32861 2431 32919 2437
rect 32861 2397 32873 2431
rect 32907 2428 32919 2431
rect 33226 2428 33232 2440
rect 32907 2400 33232 2428
rect 32907 2397 32919 2400
rect 32861 2391 32919 2397
rect 33226 2388 33232 2400
rect 33284 2388 33290 2440
rect 33410 2388 33416 2440
rect 33468 2428 33474 2440
rect 33597 2431 33655 2437
rect 33597 2428 33609 2431
rect 33468 2400 33609 2428
rect 33468 2388 33474 2400
rect 33597 2397 33609 2400
rect 33643 2397 33655 2431
rect 34698 2428 34704 2440
rect 34659 2400 34704 2428
rect 33597 2391 33655 2397
rect 34698 2388 34704 2400
rect 34756 2388 34762 2440
rect 35437 2431 35495 2437
rect 35437 2397 35449 2431
rect 35483 2428 35495 2431
rect 35894 2428 35900 2440
rect 35483 2400 35900 2428
rect 35483 2397 35495 2400
rect 35437 2391 35495 2397
rect 35894 2388 35900 2400
rect 35952 2388 35958 2440
rect 36188 2437 36216 2468
rect 36173 2431 36231 2437
rect 36173 2397 36185 2431
rect 36219 2397 36231 2431
rect 37274 2428 37280 2440
rect 37235 2400 37280 2428
rect 36173 2391 36231 2397
rect 37274 2388 37280 2400
rect 37332 2388 37338 2440
rect 28552 2363 28627 2369
rect 28552 2332 28581 2363
rect 28569 2329 28581 2332
rect 28615 2329 28627 2363
rect 29822 2360 29828 2372
rect 28569 2323 28627 2329
rect 28736 2332 29828 2360
rect 18141 2295 18199 2301
rect 18141 2292 18153 2295
rect 16868 2264 18153 2292
rect 18141 2261 18153 2264
rect 18187 2261 18199 2295
rect 18141 2255 18199 2261
rect 24118 2252 24124 2304
rect 24176 2292 24182 2304
rect 28736 2301 28764 2332
rect 29822 2320 29828 2332
rect 29880 2320 29886 2372
rect 30098 2320 30104 2372
rect 30156 2360 30162 2372
rect 30156 2332 33088 2360
rect 30156 2320 30162 2332
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 24176 2264 24593 2292
rect 24176 2252 24182 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 28721 2295 28779 2301
rect 28721 2261 28733 2295
rect 28767 2261 28779 2295
rect 28721 2255 28779 2261
rect 28810 2252 28816 2304
rect 28868 2292 28874 2304
rect 29733 2295 29791 2301
rect 29733 2292 29745 2295
rect 28868 2264 29745 2292
rect 28868 2252 28874 2264
rect 29733 2261 29745 2264
rect 29779 2261 29791 2295
rect 29733 2255 29791 2261
rect 31754 2252 31760 2304
rect 31812 2292 31818 2304
rect 33060 2301 33088 2332
rect 35342 2320 35348 2372
rect 35400 2360 35406 2372
rect 35400 2332 35894 2360
rect 35400 2320 35406 2332
rect 32309 2295 32367 2301
rect 32309 2292 32321 2295
rect 31812 2264 32321 2292
rect 31812 2252 31818 2264
rect 32309 2261 32321 2264
rect 32355 2261 32367 2295
rect 32309 2255 32367 2261
rect 33045 2295 33103 2301
rect 33045 2261 33057 2295
rect 33091 2261 33103 2295
rect 33045 2255 33103 2261
rect 33134 2252 33140 2304
rect 33192 2292 33198 2304
rect 34885 2295 34943 2301
rect 34885 2292 34897 2295
rect 33192 2264 34897 2292
rect 33192 2252 33198 2264
rect 34885 2261 34897 2264
rect 34931 2261 34943 2295
rect 35866 2292 35894 2332
rect 36357 2295 36415 2301
rect 36357 2292 36369 2295
rect 35866 2264 36369 2292
rect 34885 2255 34943 2261
rect 36357 2261 36369 2264
rect 36403 2261 36415 2295
rect 36357 2255 36415 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 3234 2048 3240 2100
rect 3292 2088 3298 2100
rect 8386 2088 8392 2100
rect 3292 2060 8392 2088
rect 3292 2048 3298 2060
rect 8386 2048 8392 2060
rect 8444 2048 8450 2100
rect 8846 2048 8852 2100
rect 8904 2088 8910 2100
rect 12342 2088 12348 2100
rect 8904 2060 12348 2088
rect 8904 2048 8910 2060
rect 12342 2048 12348 2060
rect 12400 2048 12406 2100
rect 7466 1980 7472 2032
rect 7524 2020 7530 2032
rect 13998 2020 14004 2032
rect 7524 1992 14004 2020
rect 7524 1980 7530 1992
rect 13998 1980 14004 1992
rect 14056 1980 14062 2032
rect 1946 1912 1952 1964
rect 2004 1952 2010 1964
rect 11330 1952 11336 1964
rect 2004 1924 11336 1952
rect 2004 1912 2010 1924
rect 11330 1912 11336 1924
rect 11388 1912 11394 1964
rect 1578 1844 1584 1896
rect 1636 1884 1642 1896
rect 1636 1856 2774 1884
rect 1636 1844 1642 1856
rect 2746 1748 2774 1856
rect 4982 1844 4988 1896
rect 5040 1884 5046 1896
rect 11146 1884 11152 1896
rect 5040 1856 11152 1884
rect 5040 1844 5046 1856
rect 11146 1844 11152 1856
rect 11204 1844 11210 1896
rect 3050 1776 3056 1828
rect 3108 1816 3114 1828
rect 17034 1816 17040 1828
rect 3108 1788 17040 1816
rect 3108 1776 3114 1788
rect 17034 1776 17040 1788
rect 17092 1776 17098 1828
rect 18966 1748 18972 1760
rect 2746 1720 18972 1748
rect 18966 1708 18972 1720
rect 19024 1708 19030 1760
rect 2774 1640 2780 1692
rect 2832 1680 2838 1692
rect 13262 1680 13268 1692
rect 2832 1652 13268 1680
rect 2832 1640 2838 1652
rect 13262 1640 13268 1652
rect 13320 1640 13326 1692
rect 1762 1572 1768 1624
rect 1820 1612 1826 1624
rect 4982 1612 4988 1624
rect 1820 1584 4988 1612
rect 1820 1572 1826 1584
rect 4982 1572 4988 1584
rect 5040 1572 5046 1624
rect 5166 1572 5172 1624
rect 5224 1612 5230 1624
rect 15654 1612 15660 1624
rect 5224 1584 15660 1612
rect 5224 1572 5230 1584
rect 15654 1572 15660 1584
rect 15712 1572 15718 1624
rect 3786 1368 3792 1420
rect 3844 1408 3850 1420
rect 8018 1408 8024 1420
rect 3844 1380 8024 1408
rect 3844 1368 3850 1380
rect 8018 1368 8024 1380
rect 8076 1368 8082 1420
rect 27062 1368 27068 1420
rect 27120 1408 27126 1420
rect 28810 1408 28816 1420
rect 27120 1380 28816 1408
rect 27120 1368 27126 1380
rect 28810 1368 28816 1380
rect 28868 1368 28874 1420
<< via1 >>
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 12256 47243 12308 47252
rect 12256 47209 12265 47243
rect 12265 47209 12299 47243
rect 12299 47209 12308 47243
rect 12256 47200 12308 47209
rect 20260 47243 20312 47252
rect 20260 47209 20269 47243
rect 20269 47209 20303 47243
rect 20303 47209 20312 47243
rect 20260 47200 20312 47209
rect 28264 47243 28316 47252
rect 28264 47209 28273 47243
rect 28273 47209 28307 47243
rect 28307 47209 28316 47243
rect 28264 47200 28316 47209
rect 4160 46996 4212 47048
rect 12440 46996 12492 47048
rect 20352 46996 20404 47048
rect 28080 47039 28132 47048
rect 28080 47005 28089 47039
rect 28089 47005 28123 47039
rect 28123 47005 28132 47039
rect 28080 46996 28132 47005
rect 36176 47039 36228 47048
rect 36176 47005 36185 47039
rect 36185 47005 36219 47039
rect 36219 47005 36228 47039
rect 36176 46996 36228 47005
rect 4620 46971 4672 46980
rect 4620 46937 4629 46971
rect 4629 46937 4663 46971
rect 4663 46937 4672 46971
rect 4620 46928 4672 46937
rect 36268 46903 36320 46912
rect 36268 46869 36277 46903
rect 36277 46869 36311 46903
rect 36311 46869 36320 46903
rect 36268 46860 36320 46869
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 12440 46699 12492 46708
rect 12440 46665 12449 46699
rect 12449 46665 12483 46699
rect 12483 46665 12492 46699
rect 12440 46656 12492 46665
rect 12624 46563 12676 46572
rect 12624 46529 12633 46563
rect 12633 46529 12667 46563
rect 12667 46529 12676 46563
rect 12624 46520 12676 46529
rect 15384 46520 15436 46572
rect 28080 46316 28132 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 22008 34595 22060 34604
rect 22008 34561 22017 34595
rect 22017 34561 22051 34595
rect 22051 34561 22060 34595
rect 22008 34552 22060 34561
rect 21824 34391 21876 34400
rect 21824 34357 21833 34391
rect 21833 34357 21867 34391
rect 21867 34357 21876 34391
rect 21824 34348 21876 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 17960 33940 18012 33992
rect 21180 33940 21232 33992
rect 22468 33983 22520 33992
rect 22468 33949 22477 33983
rect 22477 33949 22511 33983
rect 22511 33949 22520 33983
rect 22468 33940 22520 33949
rect 22652 33983 22704 33992
rect 22652 33949 22661 33983
rect 22661 33949 22695 33983
rect 22695 33949 22704 33983
rect 22652 33940 22704 33949
rect 20260 33872 20312 33924
rect 19432 33804 19484 33856
rect 21916 33847 21968 33856
rect 21916 33813 21925 33847
rect 21925 33813 21959 33847
rect 21959 33813 21968 33847
rect 21916 33804 21968 33813
rect 23296 33847 23348 33856
rect 23296 33813 23305 33847
rect 23305 33813 23339 33847
rect 23339 33813 23348 33847
rect 23296 33804 23348 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 20260 33643 20312 33652
rect 20260 33609 20269 33643
rect 20269 33609 20303 33643
rect 20303 33609 20312 33643
rect 20260 33600 20312 33609
rect 22008 33600 22060 33652
rect 18420 33464 18472 33516
rect 20812 33464 20864 33516
rect 22468 33532 22520 33584
rect 23296 33532 23348 33584
rect 21088 33507 21140 33516
rect 21088 33473 21097 33507
rect 21097 33473 21131 33507
rect 21131 33473 21140 33507
rect 21088 33464 21140 33473
rect 24400 33507 24452 33516
rect 24400 33473 24409 33507
rect 24409 33473 24443 33507
rect 24443 33473 24452 33507
rect 24400 33464 24452 33473
rect 16948 33396 17000 33448
rect 21180 33396 21232 33448
rect 19984 33260 20036 33312
rect 22376 33260 22428 33312
rect 24216 33303 24268 33312
rect 24216 33269 24225 33303
rect 24225 33269 24259 33303
rect 24259 33269 24268 33303
rect 24216 33260 24268 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 17960 33056 18012 33108
rect 18420 33056 18472 33108
rect 20812 33056 20864 33108
rect 24400 33056 24452 33108
rect 17408 32920 17460 32972
rect 22468 32920 22520 32972
rect 24768 32920 24820 32972
rect 17040 32895 17092 32904
rect 17040 32861 17049 32895
rect 17049 32861 17083 32895
rect 17083 32861 17092 32895
rect 17040 32852 17092 32861
rect 17684 32895 17736 32904
rect 17684 32861 17693 32895
rect 17693 32861 17727 32895
rect 17727 32861 17736 32895
rect 17684 32852 17736 32861
rect 18512 32895 18564 32904
rect 18512 32861 18521 32895
rect 18521 32861 18555 32895
rect 18555 32861 18564 32895
rect 18512 32852 18564 32861
rect 16856 32759 16908 32768
rect 16856 32725 16865 32759
rect 16865 32725 16899 32759
rect 16899 32725 16908 32759
rect 16856 32716 16908 32725
rect 19432 32784 19484 32836
rect 21180 32852 21232 32904
rect 21824 32852 21876 32904
rect 24584 32895 24636 32904
rect 21456 32784 21508 32836
rect 24584 32861 24593 32895
rect 24593 32861 24627 32895
rect 24627 32861 24636 32895
rect 24584 32852 24636 32861
rect 20628 32759 20680 32768
rect 20628 32725 20637 32759
rect 20637 32725 20671 32759
rect 20671 32725 20680 32759
rect 20628 32716 20680 32725
rect 20996 32716 21048 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 17684 32512 17736 32564
rect 21088 32512 21140 32564
rect 22652 32555 22704 32564
rect 16856 32444 16908 32496
rect 20536 32444 20588 32496
rect 22376 32487 22428 32496
rect 16672 32376 16724 32428
rect 16948 32419 17000 32428
rect 16948 32385 16957 32419
rect 16957 32385 16991 32419
rect 16991 32385 17000 32419
rect 16948 32376 17000 32385
rect 19340 32419 19392 32428
rect 19340 32385 19349 32419
rect 19349 32385 19383 32419
rect 19383 32385 19392 32419
rect 19340 32376 19392 32385
rect 19248 32308 19300 32360
rect 19616 32376 19668 32428
rect 20720 32419 20772 32428
rect 20720 32385 20729 32419
rect 20729 32385 20763 32419
rect 20763 32385 20772 32419
rect 20720 32376 20772 32385
rect 20996 32419 21048 32428
rect 20996 32385 21005 32419
rect 21005 32385 21039 32419
rect 21039 32385 21048 32419
rect 20996 32376 21048 32385
rect 22376 32453 22385 32487
rect 22385 32453 22419 32487
rect 22419 32453 22428 32487
rect 22376 32444 22428 32453
rect 22008 32376 22060 32428
rect 22284 32419 22336 32428
rect 22284 32385 22293 32419
rect 22293 32385 22327 32419
rect 22327 32385 22336 32419
rect 22284 32376 22336 32385
rect 22652 32521 22661 32555
rect 22661 32521 22695 32555
rect 22695 32521 22704 32555
rect 22652 32512 22704 32521
rect 24216 32444 24268 32496
rect 22560 32376 22612 32428
rect 23480 32376 23532 32428
rect 25412 32419 25464 32428
rect 25412 32385 25421 32419
rect 25421 32385 25455 32419
rect 25455 32385 25464 32419
rect 25412 32376 25464 32385
rect 20628 32308 20680 32360
rect 18420 32172 18472 32224
rect 18880 32172 18932 32224
rect 23572 32172 23624 32224
rect 25228 32215 25280 32224
rect 25228 32181 25237 32215
rect 25237 32181 25271 32215
rect 25271 32181 25280 32215
rect 25228 32172 25280 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 17040 31968 17092 32020
rect 18512 31968 18564 32020
rect 21456 32011 21508 32020
rect 21456 31977 21465 32011
rect 21465 31977 21499 32011
rect 21499 31977 21508 32011
rect 21456 31968 21508 31977
rect 22284 31968 22336 32020
rect 24584 31968 24636 32020
rect 23480 31900 23532 31952
rect 17408 31807 17460 31816
rect 17408 31773 17417 31807
rect 17417 31773 17451 31807
rect 17451 31773 17460 31807
rect 17408 31764 17460 31773
rect 18512 31807 18564 31816
rect 17960 31628 18012 31680
rect 18512 31773 18521 31807
rect 18521 31773 18555 31807
rect 18555 31773 18564 31807
rect 20720 31832 20772 31884
rect 19248 31807 19300 31816
rect 18512 31764 18564 31773
rect 19248 31773 19257 31807
rect 19257 31773 19291 31807
rect 19291 31773 19300 31807
rect 19248 31764 19300 31773
rect 19432 31807 19484 31816
rect 19432 31773 19441 31807
rect 19441 31773 19475 31807
rect 19475 31773 19484 31807
rect 19432 31764 19484 31773
rect 19616 31807 19668 31816
rect 19616 31773 19625 31807
rect 19625 31773 19659 31807
rect 19659 31773 19668 31807
rect 19616 31764 19668 31773
rect 18328 31739 18380 31748
rect 18328 31705 18337 31739
rect 18337 31705 18371 31739
rect 18371 31705 18380 31739
rect 18328 31696 18380 31705
rect 18420 31739 18472 31748
rect 18420 31705 18429 31739
rect 18429 31705 18463 31739
rect 18463 31705 18472 31739
rect 18420 31696 18472 31705
rect 19984 31764 20036 31816
rect 20444 31764 20496 31816
rect 22008 31832 22060 31884
rect 22468 31875 22520 31884
rect 22468 31841 22477 31875
rect 22477 31841 22511 31875
rect 22511 31841 22520 31875
rect 22468 31832 22520 31841
rect 21088 31739 21140 31748
rect 21088 31705 21097 31739
rect 21097 31705 21131 31739
rect 21131 31705 21140 31739
rect 21088 31696 21140 31705
rect 19248 31628 19300 31680
rect 22560 31764 22612 31816
rect 23388 31832 23440 31884
rect 24400 31875 24452 31884
rect 24400 31841 24409 31875
rect 24409 31841 24443 31875
rect 24443 31841 24452 31875
rect 24400 31832 24452 31841
rect 21548 31696 21600 31748
rect 22008 31696 22060 31748
rect 23204 31764 23256 31816
rect 25228 31764 25280 31816
rect 21824 31628 21876 31680
rect 22284 31671 22336 31680
rect 22284 31637 22293 31671
rect 22293 31637 22327 31671
rect 22327 31637 22336 31671
rect 22284 31628 22336 31637
rect 22376 31671 22428 31680
rect 22376 31637 22385 31671
rect 22385 31637 22419 31671
rect 22419 31637 22428 31671
rect 23572 31696 23624 31748
rect 24584 31696 24636 31748
rect 22376 31628 22428 31637
rect 24216 31628 24268 31680
rect 25044 31628 25096 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 18328 31424 18380 31476
rect 19340 31424 19392 31476
rect 21088 31424 21140 31476
rect 18052 31356 18104 31408
rect 16856 31331 16908 31340
rect 16856 31297 16865 31331
rect 16865 31297 16899 31331
rect 16899 31297 16908 31331
rect 16856 31288 16908 31297
rect 17960 31331 18012 31340
rect 17960 31297 17969 31331
rect 17969 31297 18003 31331
rect 18003 31297 18012 31331
rect 17960 31288 18012 31297
rect 18144 31331 18196 31340
rect 18144 31297 18153 31331
rect 18153 31297 18187 31331
rect 18187 31297 18196 31331
rect 18144 31288 18196 31297
rect 18512 31288 18564 31340
rect 18788 31288 18840 31340
rect 18880 31288 18932 31340
rect 20260 31288 20312 31340
rect 20628 31331 20680 31340
rect 20628 31297 20637 31331
rect 20637 31297 20671 31331
rect 20671 31297 20680 31331
rect 20628 31288 20680 31297
rect 21824 31288 21876 31340
rect 22376 31356 22428 31408
rect 25412 31424 25464 31476
rect 24216 31331 24268 31340
rect 24216 31297 24225 31331
rect 24225 31297 24259 31331
rect 24259 31297 24268 31331
rect 24216 31288 24268 31297
rect 25044 31356 25096 31408
rect 24584 31331 24636 31340
rect 24584 31297 24593 31331
rect 24593 31297 24627 31331
rect 24627 31297 24636 31331
rect 24584 31288 24636 31297
rect 24768 31288 24820 31340
rect 26240 31331 26292 31340
rect 20720 31220 20772 31272
rect 20904 31263 20956 31272
rect 20904 31229 20913 31263
rect 20913 31229 20947 31263
rect 20947 31229 20956 31263
rect 20904 31220 20956 31229
rect 22376 31263 22428 31272
rect 22376 31229 22385 31263
rect 22385 31229 22419 31263
rect 22419 31229 22428 31263
rect 22376 31220 22428 31229
rect 23296 31220 23348 31272
rect 23020 31152 23072 31204
rect 24032 31220 24084 31272
rect 26240 31297 26249 31331
rect 26249 31297 26283 31331
rect 26283 31297 26292 31331
rect 26240 31288 26292 31297
rect 16580 31084 16632 31136
rect 16764 31084 16816 31136
rect 26056 31127 26108 31136
rect 26056 31093 26065 31127
rect 26065 31093 26099 31127
rect 26099 31093 26108 31127
rect 26056 31084 26108 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 23296 30880 23348 30932
rect 17408 30812 17460 30864
rect 16948 30540 17000 30592
rect 18236 30676 18288 30728
rect 18788 30676 18840 30728
rect 19156 30676 19208 30728
rect 21548 30787 21600 30796
rect 18328 30651 18380 30660
rect 18328 30617 18337 30651
rect 18337 30617 18371 30651
rect 18371 30617 18380 30651
rect 18328 30608 18380 30617
rect 19248 30540 19300 30592
rect 20076 30540 20128 30592
rect 20628 30540 20680 30592
rect 21548 30753 21557 30787
rect 21557 30753 21591 30787
rect 21591 30753 21600 30787
rect 21548 30744 21600 30753
rect 23388 30744 23440 30796
rect 24400 30744 24452 30796
rect 22100 30676 22152 30728
rect 24584 30719 24636 30728
rect 24584 30685 24593 30719
rect 24593 30685 24627 30719
rect 24627 30685 24636 30719
rect 24584 30676 24636 30685
rect 26424 30676 26476 30728
rect 26056 30608 26108 30660
rect 23480 30540 23532 30592
rect 26608 30540 26660 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 16764 30336 16816 30388
rect 16856 30336 16908 30388
rect 20260 30379 20312 30388
rect 20260 30345 20269 30379
rect 20269 30345 20303 30379
rect 20303 30345 20312 30379
rect 20260 30336 20312 30345
rect 23296 30379 23348 30388
rect 23296 30345 23305 30379
rect 23305 30345 23339 30379
rect 23339 30345 23348 30379
rect 23296 30336 23348 30345
rect 24032 30379 24084 30388
rect 24032 30345 24041 30379
rect 24041 30345 24075 30379
rect 24075 30345 24084 30379
rect 24032 30336 24084 30345
rect 26240 30336 26292 30388
rect 20444 30268 20496 30320
rect 16764 30200 16816 30252
rect 18788 30243 18840 30252
rect 18788 30209 18797 30243
rect 18797 30209 18831 30243
rect 18831 30209 18840 30243
rect 18788 30200 18840 30209
rect 22560 30268 22612 30320
rect 26608 30268 26660 30320
rect 22192 30200 22244 30252
rect 23296 30200 23348 30252
rect 24032 30200 24084 30252
rect 24860 30200 24912 30252
rect 25136 30243 25188 30252
rect 25136 30209 25145 30243
rect 25145 30209 25179 30243
rect 25179 30209 25188 30243
rect 25136 30200 25188 30209
rect 25320 30243 25372 30252
rect 25320 30209 25329 30243
rect 25329 30209 25363 30243
rect 25363 30209 25372 30243
rect 25320 30200 25372 30209
rect 16672 30175 16724 30184
rect 14740 29996 14792 30048
rect 16672 30141 16681 30175
rect 16681 30141 16715 30175
rect 16715 30141 16724 30175
rect 16672 30132 16724 30141
rect 18512 30175 18564 30184
rect 18512 30141 18521 30175
rect 18521 30141 18555 30175
rect 18555 30141 18564 30175
rect 18512 30132 18564 30141
rect 19432 30064 19484 30116
rect 23388 30175 23440 30184
rect 23388 30141 23397 30175
rect 23397 30141 23431 30175
rect 23431 30141 23440 30175
rect 23388 30132 23440 30141
rect 22100 30064 22152 30116
rect 23204 30064 23256 30116
rect 27528 30200 27580 30252
rect 17408 29996 17460 30048
rect 18236 29996 18288 30048
rect 23664 29996 23716 30048
rect 26976 30175 27028 30184
rect 26976 30141 26985 30175
rect 26985 30141 27019 30175
rect 27019 30141 27028 30175
rect 26976 30132 27028 30141
rect 28448 29996 28500 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 14740 29835 14792 29844
rect 14740 29801 14749 29835
rect 14749 29801 14783 29835
rect 14783 29801 14792 29835
rect 14740 29792 14792 29801
rect 15568 29724 15620 29776
rect 14648 29656 14700 29708
rect 16672 29792 16724 29844
rect 18328 29792 18380 29844
rect 20536 29835 20588 29844
rect 20536 29801 20545 29835
rect 20545 29801 20579 29835
rect 20579 29801 20588 29835
rect 20536 29792 20588 29801
rect 22376 29792 22428 29844
rect 23388 29835 23440 29844
rect 23388 29801 23397 29835
rect 23397 29801 23431 29835
rect 23431 29801 23440 29835
rect 23388 29792 23440 29801
rect 25136 29792 25188 29844
rect 22836 29724 22888 29776
rect 20628 29656 20680 29708
rect 20996 29656 21048 29708
rect 25228 29699 25280 29708
rect 25228 29665 25237 29699
rect 25237 29665 25271 29699
rect 25271 29665 25280 29699
rect 25228 29656 25280 29665
rect 26424 29699 26476 29708
rect 26424 29665 26433 29699
rect 26433 29665 26467 29699
rect 26467 29665 26476 29699
rect 26424 29656 26476 29665
rect 14740 29588 14792 29640
rect 16672 29631 16724 29640
rect 16672 29597 16706 29631
rect 16706 29597 16724 29631
rect 15292 29520 15344 29572
rect 16672 29588 16724 29597
rect 20260 29588 20312 29640
rect 23296 29588 23348 29640
rect 28448 29631 28500 29640
rect 16580 29520 16632 29572
rect 23112 29520 23164 29572
rect 28448 29597 28457 29631
rect 28457 29597 28491 29631
rect 28491 29597 28500 29631
rect 28448 29588 28500 29597
rect 14924 29452 14976 29504
rect 18052 29452 18104 29504
rect 18236 29452 18288 29504
rect 20444 29452 20496 29504
rect 21088 29452 21140 29504
rect 21640 29452 21692 29504
rect 21916 29495 21968 29504
rect 21916 29461 21941 29495
rect 21941 29461 21968 29495
rect 21916 29452 21968 29461
rect 22100 29452 22152 29504
rect 22744 29495 22796 29504
rect 22744 29461 22769 29495
rect 22769 29461 22796 29495
rect 22744 29452 22796 29461
rect 24952 29452 25004 29504
rect 25872 29452 25924 29504
rect 26608 29452 26660 29504
rect 27252 29452 27304 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4620 29248 4672 29300
rect 16764 29291 16816 29300
rect 13084 29155 13136 29164
rect 13084 29121 13093 29155
rect 13093 29121 13127 29155
rect 13127 29121 13136 29155
rect 13084 29112 13136 29121
rect 14648 29180 14700 29232
rect 16764 29257 16773 29291
rect 16773 29257 16807 29291
rect 16807 29257 16816 29291
rect 16764 29248 16816 29257
rect 18144 29248 18196 29300
rect 20260 29248 20312 29300
rect 20904 29248 20956 29300
rect 14464 29155 14516 29164
rect 14464 29121 14498 29155
rect 14498 29121 14516 29155
rect 16948 29155 17000 29164
rect 12624 29044 12676 29096
rect 14464 29112 14516 29121
rect 16948 29121 16957 29155
rect 16957 29121 16991 29155
rect 16991 29121 17000 29155
rect 16948 29112 17000 29121
rect 18052 29112 18104 29164
rect 20904 29112 20956 29164
rect 22192 29248 22244 29300
rect 23020 29291 23072 29300
rect 22284 29180 22336 29232
rect 23020 29257 23029 29291
rect 23029 29257 23063 29291
rect 23063 29257 23072 29291
rect 23020 29248 23072 29257
rect 23664 29291 23716 29300
rect 23664 29257 23673 29291
rect 23673 29257 23707 29291
rect 23707 29257 23716 29291
rect 23664 29248 23716 29257
rect 27528 29291 27580 29300
rect 22192 29112 22244 29164
rect 23112 29180 23164 29232
rect 24584 29180 24636 29232
rect 24952 29180 25004 29232
rect 24032 29112 24084 29164
rect 25964 29155 26016 29164
rect 25964 29121 25973 29155
rect 25973 29121 26007 29155
rect 26007 29121 26016 29155
rect 25964 29112 26016 29121
rect 12440 28908 12492 28960
rect 16672 28976 16724 29028
rect 23480 28976 23532 29028
rect 24860 29044 24912 29096
rect 26056 29087 26108 29096
rect 26056 29053 26065 29087
rect 26065 29053 26099 29087
rect 26099 29053 26108 29087
rect 26332 29180 26384 29232
rect 26700 29180 26752 29232
rect 27528 29257 27537 29291
rect 27537 29257 27571 29291
rect 27571 29257 27580 29291
rect 27528 29248 27580 29257
rect 26056 29044 26108 29053
rect 24400 28976 24452 29028
rect 25688 28976 25740 29028
rect 27252 29155 27304 29164
rect 27252 29121 27261 29155
rect 27261 29121 27295 29155
rect 27295 29121 27304 29155
rect 27252 29112 27304 29121
rect 15660 28908 15712 28960
rect 22836 28951 22888 28960
rect 22836 28917 22845 28951
rect 22845 28917 22879 28951
rect 22879 28917 22888 28951
rect 22836 28908 22888 28917
rect 26148 28908 26200 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 16580 28704 16632 28756
rect 20720 28704 20772 28756
rect 22468 28704 22520 28756
rect 25228 28704 25280 28756
rect 26332 28704 26384 28756
rect 15844 28568 15896 28620
rect 19248 28568 19300 28620
rect 9956 28500 10008 28552
rect 11060 28543 11112 28552
rect 11060 28509 11069 28543
rect 11069 28509 11103 28543
rect 11103 28509 11112 28543
rect 11060 28500 11112 28509
rect 8392 28432 8444 28484
rect 9588 28432 9640 28484
rect 11244 28543 11296 28552
rect 11244 28509 11253 28543
rect 11253 28509 11287 28543
rect 11287 28509 11296 28543
rect 11244 28500 11296 28509
rect 12440 28543 12492 28552
rect 12440 28509 12474 28543
rect 12474 28509 12492 28543
rect 14648 28543 14700 28552
rect 9772 28364 9824 28416
rect 10784 28407 10836 28416
rect 10784 28373 10793 28407
rect 10793 28373 10827 28407
rect 10827 28373 10836 28407
rect 10784 28364 10836 28373
rect 11336 28432 11388 28484
rect 12440 28500 12492 28509
rect 14648 28509 14657 28543
rect 14657 28509 14691 28543
rect 14691 28509 14700 28543
rect 14648 28500 14700 28509
rect 15108 28432 15160 28484
rect 16580 28543 16632 28552
rect 16580 28509 16589 28543
rect 16589 28509 16623 28543
rect 16623 28509 16632 28543
rect 20812 28636 20864 28688
rect 21916 28636 21968 28688
rect 22008 28636 22060 28688
rect 21456 28568 21508 28620
rect 22652 28568 22704 28620
rect 24768 28568 24820 28620
rect 16580 28500 16632 28509
rect 17500 28432 17552 28484
rect 22100 28500 22152 28552
rect 19984 28432 20036 28484
rect 21088 28432 21140 28484
rect 22744 28500 22796 28552
rect 23296 28500 23348 28552
rect 23664 28500 23716 28552
rect 23848 28500 23900 28552
rect 25320 28500 25372 28552
rect 26424 28500 26476 28552
rect 26884 28500 26936 28552
rect 13544 28407 13596 28416
rect 13544 28373 13553 28407
rect 13553 28373 13587 28407
rect 13587 28373 13596 28407
rect 13544 28364 13596 28373
rect 16028 28407 16080 28416
rect 16028 28373 16037 28407
rect 16037 28373 16071 28407
rect 16071 28373 16080 28407
rect 16028 28364 16080 28373
rect 20168 28364 20220 28416
rect 20260 28364 20312 28416
rect 21456 28364 21508 28416
rect 21916 28407 21968 28416
rect 21916 28373 21925 28407
rect 21925 28373 21959 28407
rect 21959 28373 21968 28407
rect 21916 28364 21968 28373
rect 22652 28364 22704 28416
rect 23940 28432 23992 28484
rect 25872 28432 25924 28484
rect 23020 28364 23072 28416
rect 26056 28364 26108 28416
rect 26332 28407 26384 28416
rect 26332 28373 26341 28407
rect 26341 28373 26375 28407
rect 26375 28373 26384 28407
rect 26332 28364 26384 28373
rect 27804 28432 27856 28484
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 15108 28203 15160 28212
rect 9680 28092 9732 28144
rect 12716 28092 12768 28144
rect 15108 28169 15117 28203
rect 15117 28169 15151 28203
rect 15151 28169 15160 28203
rect 15108 28160 15160 28169
rect 18512 28160 18564 28212
rect 20628 28203 20680 28212
rect 20628 28169 20637 28203
rect 20637 28169 20671 28203
rect 20671 28169 20680 28203
rect 20628 28160 20680 28169
rect 25320 28160 25372 28212
rect 26148 28160 26200 28212
rect 27804 28203 27856 28212
rect 27804 28169 27813 28203
rect 27813 28169 27847 28203
rect 27847 28169 27856 28203
rect 27804 28160 27856 28169
rect 14188 28092 14240 28144
rect 8576 28067 8628 28076
rect 8576 28033 8585 28067
rect 8585 28033 8619 28067
rect 8619 28033 8628 28067
rect 8576 28024 8628 28033
rect 8760 28067 8812 28076
rect 8760 28033 8769 28067
rect 8769 28033 8803 28067
rect 8803 28033 8812 28067
rect 8760 28024 8812 28033
rect 11980 28067 12032 28076
rect 11980 28033 12014 28067
rect 12014 28033 12032 28067
rect 11980 28024 12032 28033
rect 15292 28067 15344 28076
rect 9128 27820 9180 27872
rect 13544 27956 13596 28008
rect 15292 28033 15301 28067
rect 15301 28033 15335 28067
rect 15335 28033 15344 28067
rect 15292 28024 15344 28033
rect 16028 28092 16080 28144
rect 23664 28092 23716 28144
rect 26056 28135 26108 28144
rect 26056 28101 26065 28135
rect 26065 28101 26099 28135
rect 26099 28101 26108 28135
rect 26056 28092 26108 28101
rect 15568 28067 15620 28076
rect 15568 28033 15577 28067
rect 15577 28033 15611 28067
rect 15611 28033 15620 28067
rect 15568 28024 15620 28033
rect 15660 28067 15712 28076
rect 15660 28033 15669 28067
rect 15669 28033 15703 28067
rect 15703 28033 15712 28067
rect 15660 28024 15712 28033
rect 15936 28024 15988 28076
rect 16856 28067 16908 28076
rect 16856 28033 16865 28067
rect 16865 28033 16899 28067
rect 16899 28033 16908 28067
rect 16856 28024 16908 28033
rect 17132 28024 17184 28076
rect 18604 28067 18656 28076
rect 18604 28033 18613 28067
rect 18613 28033 18647 28067
rect 18647 28033 18656 28067
rect 18604 28024 18656 28033
rect 19340 28067 19392 28076
rect 17776 27999 17828 28008
rect 17776 27965 17785 27999
rect 17785 27965 17819 27999
rect 17819 27965 17828 27999
rect 17776 27956 17828 27965
rect 19340 28033 19349 28067
rect 19349 28033 19383 28067
rect 19383 28033 19392 28067
rect 19340 28024 19392 28033
rect 20168 28067 20220 28076
rect 20168 28033 20177 28067
rect 20177 28033 20211 28067
rect 20211 28033 20220 28067
rect 20168 28024 20220 28033
rect 15568 27888 15620 27940
rect 19248 27956 19300 28008
rect 21088 28024 21140 28076
rect 21272 28067 21324 28076
rect 21272 28033 21281 28067
rect 21281 28033 21315 28067
rect 21315 28033 21324 28067
rect 21272 28024 21324 28033
rect 22284 28024 22336 28076
rect 23756 28067 23808 28076
rect 23756 28033 23765 28067
rect 23765 28033 23799 28067
rect 23799 28033 23808 28067
rect 23756 28024 23808 28033
rect 24584 28067 24636 28076
rect 24584 28033 24593 28067
rect 24593 28033 24627 28067
rect 24627 28033 24636 28067
rect 24584 28024 24636 28033
rect 25688 28024 25740 28076
rect 26976 28067 27028 28076
rect 9956 27820 10008 27872
rect 10508 27820 10560 27872
rect 10600 27863 10652 27872
rect 10600 27829 10609 27863
rect 10609 27829 10643 27863
rect 10643 27829 10652 27863
rect 10600 27820 10652 27829
rect 14004 27820 14056 27872
rect 14556 27820 14608 27872
rect 17960 27820 18012 27872
rect 20076 27820 20128 27872
rect 20628 27956 20680 28008
rect 21732 27956 21784 28008
rect 21916 27956 21968 28008
rect 23940 27999 23992 28008
rect 23940 27965 23949 27999
rect 23949 27965 23983 27999
rect 23983 27965 23992 27999
rect 23940 27956 23992 27965
rect 25780 27956 25832 28008
rect 26976 28033 26985 28067
rect 26985 28033 27019 28067
rect 27019 28033 27028 28067
rect 26976 28024 27028 28033
rect 26332 27956 26384 28008
rect 20720 27820 20772 27872
rect 21088 27863 21140 27872
rect 21088 27829 21097 27863
rect 21097 27829 21131 27863
rect 21131 27829 21140 27863
rect 21088 27820 21140 27829
rect 24584 27820 24636 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 8392 27659 8444 27668
rect 8392 27625 8401 27659
rect 8401 27625 8435 27659
rect 8435 27625 8444 27659
rect 8392 27616 8444 27625
rect 15844 27659 15896 27668
rect 15844 27625 15853 27659
rect 15853 27625 15887 27659
rect 15887 27625 15896 27659
rect 15844 27616 15896 27625
rect 9680 27591 9732 27600
rect 9680 27557 9689 27591
rect 9689 27557 9723 27591
rect 9723 27557 9732 27591
rect 9680 27548 9732 27557
rect 17960 27616 18012 27668
rect 20076 27616 20128 27668
rect 21732 27616 21784 27668
rect 22192 27616 22244 27668
rect 23296 27659 23348 27668
rect 23296 27625 23305 27659
rect 23305 27625 23339 27659
rect 23339 27625 23348 27659
rect 23296 27616 23348 27625
rect 8116 27480 8168 27532
rect 8024 27455 8076 27464
rect 8024 27421 8033 27455
rect 8033 27421 8067 27455
rect 8067 27421 8076 27455
rect 8024 27412 8076 27421
rect 8944 27455 8996 27464
rect 8944 27421 8953 27455
rect 8953 27421 8987 27455
rect 8987 27421 8996 27455
rect 8944 27412 8996 27421
rect 9128 27455 9180 27464
rect 9128 27421 9137 27455
rect 9137 27421 9171 27455
rect 9171 27421 9180 27455
rect 9128 27412 9180 27421
rect 9220 27455 9272 27464
rect 9220 27421 9229 27455
rect 9229 27421 9263 27455
rect 9263 27421 9272 27455
rect 10324 27480 10376 27532
rect 10600 27480 10652 27532
rect 12716 27523 12768 27532
rect 12716 27489 12725 27523
rect 12725 27489 12759 27523
rect 12759 27489 12768 27523
rect 12716 27480 12768 27489
rect 13544 27480 13596 27532
rect 15292 27480 15344 27532
rect 19432 27548 19484 27600
rect 20996 27591 21048 27600
rect 20996 27557 21005 27591
rect 21005 27557 21039 27591
rect 21039 27557 21048 27591
rect 20996 27548 21048 27557
rect 21088 27548 21140 27600
rect 23848 27548 23900 27600
rect 9220 27412 9272 27421
rect 10508 27412 10560 27464
rect 10784 27412 10836 27464
rect 12992 27455 13044 27464
rect 12992 27421 13001 27455
rect 13001 27421 13035 27455
rect 13035 27421 13044 27455
rect 12992 27412 13044 27421
rect 16488 27455 16540 27464
rect 9864 27344 9916 27396
rect 12256 27344 12308 27396
rect 16488 27421 16497 27455
rect 16497 27421 16531 27455
rect 16531 27421 16540 27455
rect 16488 27412 16540 27421
rect 17316 27412 17368 27464
rect 17776 27412 17828 27464
rect 19156 27480 19208 27532
rect 19984 27480 20036 27532
rect 22008 27480 22060 27532
rect 18972 27412 19024 27464
rect 20720 27455 20772 27464
rect 20720 27421 20729 27455
rect 20729 27421 20763 27455
rect 20763 27421 20772 27455
rect 20720 27412 20772 27421
rect 21088 27412 21140 27464
rect 21272 27412 21324 27464
rect 22192 27455 22244 27464
rect 22192 27421 22201 27455
rect 22201 27421 22235 27455
rect 22235 27421 22244 27455
rect 22192 27412 22244 27421
rect 22744 27412 22796 27464
rect 22928 27455 22980 27464
rect 22928 27421 22937 27455
rect 22937 27421 22971 27455
rect 22971 27421 22980 27455
rect 22928 27412 22980 27421
rect 24400 27455 24452 27464
rect 24400 27421 24409 27455
rect 24409 27421 24443 27455
rect 24443 27421 24452 27455
rect 24400 27412 24452 27421
rect 24584 27455 24636 27464
rect 24584 27421 24593 27455
rect 24593 27421 24627 27455
rect 24627 27421 24636 27455
rect 24584 27412 24636 27421
rect 24768 27455 24820 27464
rect 24768 27421 24777 27455
rect 24777 27421 24811 27455
rect 24811 27421 24820 27455
rect 24768 27412 24820 27421
rect 25688 27455 25740 27464
rect 25688 27421 25697 27455
rect 25697 27421 25731 27455
rect 25731 27421 25740 27455
rect 25688 27412 25740 27421
rect 25780 27412 25832 27464
rect 28172 27548 28224 27600
rect 26976 27480 27028 27532
rect 26148 27412 26200 27464
rect 16120 27344 16172 27396
rect 16856 27344 16908 27396
rect 20628 27344 20680 27396
rect 22652 27344 22704 27396
rect 23756 27344 23808 27396
rect 25228 27344 25280 27396
rect 25504 27344 25556 27396
rect 28356 27412 28408 27464
rect 8760 27276 8812 27328
rect 11060 27276 11112 27328
rect 11612 27276 11664 27328
rect 14096 27276 14148 27328
rect 14832 27276 14884 27328
rect 16396 27276 16448 27328
rect 17960 27276 18012 27328
rect 24952 27319 25004 27328
rect 24952 27285 24961 27319
rect 24961 27285 24995 27319
rect 24995 27285 25004 27319
rect 24952 27276 25004 27285
rect 27068 27319 27120 27328
rect 27068 27285 27077 27319
rect 27077 27285 27111 27319
rect 27111 27285 27120 27319
rect 27068 27276 27120 27285
rect 27528 27319 27580 27328
rect 27528 27285 27537 27319
rect 27537 27285 27571 27319
rect 27571 27285 27580 27319
rect 27528 27276 27580 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 8024 27115 8076 27124
rect 8024 27081 8033 27115
rect 8033 27081 8067 27115
rect 8067 27081 8076 27115
rect 8024 27072 8076 27081
rect 9220 27072 9272 27124
rect 9864 27115 9916 27124
rect 9864 27081 9873 27115
rect 9873 27081 9907 27115
rect 9907 27081 9916 27115
rect 9864 27072 9916 27081
rect 11244 27072 11296 27124
rect 13084 27072 13136 27124
rect 8944 27004 8996 27056
rect 8392 26936 8444 26988
rect 8760 26936 8812 26988
rect 9772 26936 9824 26988
rect 8300 26868 8352 26920
rect 8576 26868 8628 26920
rect 8944 26911 8996 26920
rect 8944 26877 8953 26911
rect 8953 26877 8987 26911
rect 8987 26877 8996 26911
rect 8944 26868 8996 26877
rect 10600 26936 10652 26988
rect 10692 26911 10744 26920
rect 8852 26800 8904 26852
rect 10692 26877 10701 26911
rect 10701 26877 10735 26911
rect 10735 26877 10744 26911
rect 10692 26868 10744 26877
rect 11152 26868 11204 26920
rect 12164 26911 12216 26920
rect 12164 26877 12173 26911
rect 12173 26877 12207 26911
rect 12207 26877 12216 26911
rect 12164 26868 12216 26877
rect 12808 27004 12860 27056
rect 14464 27072 14516 27124
rect 13268 26936 13320 26988
rect 14096 26979 14148 26988
rect 14096 26945 14105 26979
rect 14105 26945 14139 26979
rect 14139 26945 14148 26979
rect 14096 26936 14148 26945
rect 15200 27072 15252 27124
rect 15844 27072 15896 27124
rect 18604 27072 18656 27124
rect 20076 27115 20128 27124
rect 20076 27081 20085 27115
rect 20085 27081 20119 27115
rect 20119 27081 20128 27115
rect 20076 27072 20128 27081
rect 22192 27072 22244 27124
rect 22744 27072 22796 27124
rect 25504 27115 25556 27124
rect 15016 27004 15068 27056
rect 14924 26979 14976 26988
rect 14924 26945 14933 26979
rect 14933 26945 14967 26979
rect 14967 26945 14976 26979
rect 15108 26979 15160 27012
rect 15108 26960 15117 26979
rect 15117 26960 15151 26979
rect 15151 26960 15160 26979
rect 14924 26936 14976 26945
rect 15200 26936 15252 26988
rect 15476 26936 15528 26988
rect 15936 26979 15988 26988
rect 15936 26945 15945 26979
rect 15945 26945 15979 26979
rect 15979 26945 15988 26979
rect 15936 26936 15988 26945
rect 16212 26936 16264 26988
rect 17960 27004 18012 27056
rect 17224 26936 17276 26988
rect 17868 26979 17920 26988
rect 17868 26945 17877 26979
rect 17877 26945 17911 26979
rect 17911 26945 17920 26979
rect 17868 26936 17920 26945
rect 15568 26868 15620 26920
rect 16028 26868 16080 26920
rect 13268 26800 13320 26852
rect 8024 26732 8076 26784
rect 10416 26732 10468 26784
rect 15200 26800 15252 26852
rect 16488 26800 16540 26852
rect 16856 26800 16908 26852
rect 19340 27004 19392 27056
rect 25504 27081 25513 27115
rect 25513 27081 25547 27115
rect 25547 27081 25556 27115
rect 25504 27072 25556 27081
rect 25780 27072 25832 27124
rect 26056 27072 26108 27124
rect 28356 27115 28408 27124
rect 28356 27081 28365 27115
rect 28365 27081 28399 27115
rect 28399 27081 28408 27115
rect 28356 27072 28408 27081
rect 19984 26936 20036 26988
rect 22744 26936 22796 26988
rect 22928 26936 22980 26988
rect 23112 26936 23164 26988
rect 26884 27004 26936 27056
rect 28448 27004 28500 27056
rect 14280 26732 14332 26784
rect 14924 26732 14976 26784
rect 16948 26732 17000 26784
rect 18972 26868 19024 26920
rect 22008 26911 22060 26920
rect 22008 26877 22017 26911
rect 22017 26877 22051 26911
rect 22051 26877 22060 26911
rect 22008 26868 22060 26877
rect 19432 26800 19484 26852
rect 20628 26800 20680 26852
rect 23112 26800 23164 26852
rect 19524 26732 19576 26784
rect 19984 26732 20036 26784
rect 22100 26775 22152 26784
rect 22100 26741 22109 26775
rect 22109 26741 22143 26775
rect 22143 26741 22152 26775
rect 22100 26732 22152 26741
rect 22560 26732 22612 26784
rect 22928 26775 22980 26784
rect 22928 26741 22937 26775
rect 22937 26741 22971 26775
rect 22971 26741 22980 26775
rect 25780 26936 25832 26988
rect 25688 26868 25740 26920
rect 27160 26979 27212 26988
rect 27160 26945 27169 26979
rect 27169 26945 27203 26979
rect 27203 26945 27212 26979
rect 27160 26936 27212 26945
rect 24676 26800 24728 26852
rect 26148 26868 26200 26920
rect 22928 26732 22980 26741
rect 25228 26732 25280 26784
rect 26976 26732 27028 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 8024 26571 8076 26580
rect 8024 26537 8033 26571
rect 8033 26537 8067 26571
rect 8067 26537 8076 26571
rect 8024 26528 8076 26537
rect 8760 26528 8812 26580
rect 8668 26460 8720 26512
rect 10692 26528 10744 26580
rect 11152 26571 11204 26580
rect 11152 26537 11161 26571
rect 11161 26537 11195 26571
rect 11195 26537 11204 26571
rect 11152 26528 11204 26537
rect 11980 26528 12032 26580
rect 15844 26528 15896 26580
rect 9036 26460 9088 26512
rect 8300 26392 8352 26444
rect 9312 26392 9364 26444
rect 11336 26460 11388 26512
rect 10416 26435 10468 26444
rect 10416 26401 10425 26435
rect 10425 26401 10459 26435
rect 10459 26401 10468 26435
rect 10416 26392 10468 26401
rect 10784 26392 10836 26444
rect 14096 26460 14148 26512
rect 14648 26460 14700 26512
rect 15200 26460 15252 26512
rect 17408 26528 17460 26580
rect 17868 26528 17920 26580
rect 19340 26571 19392 26580
rect 19340 26537 19349 26571
rect 19349 26537 19383 26571
rect 19383 26537 19392 26571
rect 19340 26528 19392 26537
rect 20260 26528 20312 26580
rect 20812 26571 20864 26580
rect 20812 26537 20821 26571
rect 20821 26537 20855 26571
rect 20855 26537 20864 26571
rect 20812 26528 20864 26537
rect 20904 26528 20956 26580
rect 22836 26528 22888 26580
rect 27160 26528 27212 26580
rect 8944 26367 8996 26376
rect 8944 26333 8953 26367
rect 8953 26333 8987 26367
rect 8987 26333 8996 26367
rect 8944 26324 8996 26333
rect 9128 26367 9180 26376
rect 9128 26333 9137 26367
rect 9137 26333 9171 26367
rect 9171 26333 9180 26367
rect 9128 26324 9180 26333
rect 10324 26367 10376 26376
rect 8300 26256 8352 26308
rect 10324 26333 10333 26367
rect 10333 26333 10367 26367
rect 10367 26333 10376 26367
rect 10324 26324 10376 26333
rect 11336 26367 11388 26376
rect 11336 26333 11345 26367
rect 11345 26333 11379 26367
rect 11379 26333 11388 26367
rect 11336 26324 11388 26333
rect 11520 26367 11572 26376
rect 11520 26333 11529 26367
rect 11529 26333 11563 26367
rect 11563 26333 11572 26367
rect 11520 26324 11572 26333
rect 11612 26367 11664 26376
rect 11612 26333 11621 26367
rect 11621 26333 11655 26367
rect 11655 26333 11664 26367
rect 11612 26324 11664 26333
rect 12440 26324 12492 26376
rect 14924 26392 14976 26444
rect 12992 26324 13044 26376
rect 13268 26367 13320 26376
rect 13268 26333 13277 26367
rect 13277 26333 13311 26367
rect 13311 26333 13320 26367
rect 13268 26324 13320 26333
rect 14648 26324 14700 26376
rect 15292 26392 15344 26444
rect 22100 26460 22152 26512
rect 23020 26460 23072 26512
rect 28172 26460 28224 26512
rect 15844 26324 15896 26376
rect 15292 26256 15344 26308
rect 7748 26188 7800 26240
rect 12348 26188 12400 26240
rect 12532 26188 12584 26240
rect 13728 26188 13780 26240
rect 16120 26324 16172 26376
rect 16948 26392 17000 26444
rect 16396 26367 16448 26376
rect 16396 26333 16405 26367
rect 16405 26333 16439 26367
rect 16439 26333 16448 26367
rect 16396 26324 16448 26333
rect 16672 26324 16724 26376
rect 17224 26367 17276 26376
rect 17224 26333 17233 26367
rect 17233 26333 17267 26367
rect 17267 26333 17276 26367
rect 17224 26324 17276 26333
rect 19248 26367 19300 26376
rect 16856 26256 16908 26308
rect 17040 26256 17092 26308
rect 19248 26333 19257 26367
rect 19257 26333 19291 26367
rect 19291 26333 19300 26367
rect 19248 26324 19300 26333
rect 19340 26324 19392 26376
rect 20720 26324 20772 26376
rect 20996 26392 21048 26444
rect 21088 26324 21140 26376
rect 21548 26324 21600 26376
rect 22008 26392 22060 26444
rect 22100 26367 22152 26376
rect 22100 26333 22109 26367
rect 22109 26333 22143 26367
rect 22143 26333 22152 26367
rect 22652 26367 22704 26376
rect 22100 26324 22152 26333
rect 22652 26333 22661 26367
rect 22661 26333 22695 26367
rect 22695 26333 22704 26367
rect 22652 26324 22704 26333
rect 23664 26392 23716 26444
rect 26884 26435 26936 26444
rect 26884 26401 26893 26435
rect 26893 26401 26927 26435
rect 26927 26401 26936 26435
rect 26884 26392 26936 26401
rect 23296 26324 23348 26376
rect 24400 26367 24452 26376
rect 17960 26299 18012 26308
rect 17960 26265 17969 26299
rect 17969 26265 18003 26299
rect 18003 26265 18012 26299
rect 17960 26256 18012 26265
rect 19524 26256 19576 26308
rect 24400 26333 24409 26367
rect 24409 26333 24443 26367
rect 24443 26333 24452 26367
rect 24400 26324 24452 26333
rect 24952 26324 25004 26376
rect 25872 26324 25924 26376
rect 26148 26256 26200 26308
rect 28448 26324 28500 26376
rect 17224 26188 17276 26240
rect 17592 26188 17644 26240
rect 18328 26231 18380 26240
rect 18328 26197 18337 26231
rect 18337 26197 18371 26231
rect 18371 26197 18380 26231
rect 18328 26188 18380 26197
rect 20260 26188 20312 26240
rect 20444 26188 20496 26240
rect 20904 26188 20956 26240
rect 23480 26188 23532 26240
rect 26976 26256 27028 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 9036 25984 9088 26036
rect 9128 25984 9180 26036
rect 11336 25984 11388 26036
rect 12256 25984 12308 26036
rect 12440 25984 12492 26036
rect 15844 25984 15896 26036
rect 16028 26027 16080 26036
rect 16028 25993 16037 26027
rect 16037 25993 16071 26027
rect 16071 25993 16080 26027
rect 16028 25984 16080 25993
rect 9772 25916 9824 25968
rect 11520 25916 11572 25968
rect 14188 25916 14240 25968
rect 20996 25984 21048 26036
rect 22284 25984 22336 26036
rect 23664 25984 23716 26036
rect 26240 25984 26292 26036
rect 26884 25984 26936 26036
rect 16304 25916 16356 25968
rect 7748 25891 7800 25900
rect 7748 25857 7757 25891
rect 7757 25857 7791 25891
rect 7791 25857 7800 25891
rect 7748 25848 7800 25857
rect 7932 25891 7984 25900
rect 7932 25857 7941 25891
rect 7941 25857 7975 25891
rect 7975 25857 7984 25891
rect 7932 25848 7984 25857
rect 8116 25891 8168 25900
rect 8116 25857 8125 25891
rect 8125 25857 8159 25891
rect 8159 25857 8168 25891
rect 8116 25848 8168 25857
rect 8392 25848 8444 25900
rect 9404 25848 9456 25900
rect 10784 25891 10836 25900
rect 8024 25823 8076 25832
rect 8024 25789 8033 25823
rect 8033 25789 8067 25823
rect 8067 25789 8076 25823
rect 9680 25823 9732 25832
rect 8024 25780 8076 25789
rect 9680 25789 9689 25823
rect 9689 25789 9723 25823
rect 9723 25789 9732 25823
rect 9680 25780 9732 25789
rect 10784 25857 10793 25891
rect 10793 25857 10827 25891
rect 10827 25857 10836 25891
rect 10784 25848 10836 25857
rect 13268 25848 13320 25900
rect 14096 25891 14148 25900
rect 14096 25857 14105 25891
rect 14105 25857 14139 25891
rect 14139 25857 14148 25891
rect 14096 25848 14148 25857
rect 12992 25823 13044 25832
rect 12992 25789 13001 25823
rect 13001 25789 13035 25823
rect 13035 25789 13044 25823
rect 12992 25780 13044 25789
rect 10784 25712 10836 25764
rect 12348 25712 12400 25764
rect 13176 25823 13228 25832
rect 13176 25789 13185 25823
rect 13185 25789 13219 25823
rect 13219 25789 13228 25823
rect 13176 25780 13228 25789
rect 13728 25780 13780 25832
rect 16120 25780 16172 25832
rect 13360 25712 13412 25764
rect 15200 25712 15252 25764
rect 17960 25848 18012 25900
rect 16764 25780 16816 25832
rect 17500 25780 17552 25832
rect 19432 25848 19484 25900
rect 18788 25823 18840 25832
rect 18788 25789 18797 25823
rect 18797 25789 18831 25823
rect 18831 25789 18840 25823
rect 18788 25780 18840 25789
rect 20812 25848 20864 25900
rect 17408 25755 17460 25764
rect 17408 25721 17417 25755
rect 17417 25721 17451 25755
rect 17451 25721 17460 25755
rect 17408 25712 17460 25721
rect 17684 25712 17736 25764
rect 20628 25780 20680 25832
rect 21456 25780 21508 25832
rect 21916 25780 21968 25832
rect 21272 25712 21324 25764
rect 22100 25891 22152 25900
rect 22100 25857 22109 25891
rect 22109 25857 22143 25891
rect 22143 25857 22152 25891
rect 22284 25891 22336 25900
rect 22100 25848 22152 25857
rect 22284 25857 22293 25891
rect 22293 25857 22327 25891
rect 22327 25857 22336 25891
rect 22284 25848 22336 25857
rect 22560 25848 22612 25900
rect 23388 25916 23440 25968
rect 26792 25916 26844 25968
rect 23480 25891 23532 25900
rect 23480 25857 23489 25891
rect 23489 25857 23523 25891
rect 23523 25857 23532 25891
rect 23480 25848 23532 25857
rect 23664 25891 23716 25900
rect 23664 25857 23685 25891
rect 23685 25857 23716 25891
rect 23664 25848 23716 25857
rect 24032 25848 24084 25900
rect 26148 25848 26200 25900
rect 27528 25916 27580 25968
rect 24676 25780 24728 25832
rect 25504 25712 25556 25764
rect 25780 25712 25832 25764
rect 8484 25687 8536 25696
rect 8484 25653 8493 25687
rect 8493 25653 8527 25687
rect 8527 25653 8536 25687
rect 8484 25644 8536 25653
rect 9036 25644 9088 25696
rect 10048 25644 10100 25696
rect 13268 25644 13320 25696
rect 19340 25644 19392 25696
rect 20444 25644 20496 25696
rect 21916 25644 21968 25696
rect 24032 25644 24084 25696
rect 24400 25644 24452 25696
rect 28448 25644 28500 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 8024 25440 8076 25492
rect 9680 25440 9732 25492
rect 10324 25440 10376 25492
rect 10692 25483 10744 25492
rect 10692 25449 10701 25483
rect 10701 25449 10735 25483
rect 10735 25449 10744 25483
rect 10692 25440 10744 25449
rect 8392 25415 8444 25424
rect 8392 25381 8401 25415
rect 8401 25381 8435 25415
rect 8435 25381 8444 25415
rect 8392 25372 8444 25381
rect 9128 25372 9180 25424
rect 12164 25440 12216 25492
rect 14924 25440 14976 25492
rect 15108 25483 15160 25492
rect 15108 25449 15117 25483
rect 15117 25449 15151 25483
rect 15151 25449 15160 25483
rect 15108 25440 15160 25449
rect 15568 25440 15620 25492
rect 16028 25440 16080 25492
rect 17408 25483 17460 25492
rect 17408 25449 17417 25483
rect 17417 25449 17451 25483
rect 17451 25449 17460 25483
rect 17408 25440 17460 25449
rect 17592 25483 17644 25492
rect 17592 25449 17601 25483
rect 17601 25449 17635 25483
rect 17635 25449 17644 25483
rect 17592 25440 17644 25449
rect 19248 25440 19300 25492
rect 22284 25440 22336 25492
rect 26976 25440 27028 25492
rect 8668 25304 8720 25356
rect 9772 25304 9824 25356
rect 10416 25304 10468 25356
rect 14004 25372 14056 25424
rect 15016 25372 15068 25424
rect 7012 25279 7064 25288
rect 7012 25245 7021 25279
rect 7021 25245 7055 25279
rect 7055 25245 7064 25279
rect 7012 25236 7064 25245
rect 8484 25236 8536 25288
rect 8392 25168 8444 25220
rect 9956 25236 10008 25288
rect 12900 25304 12952 25356
rect 10140 25168 10192 25220
rect 11796 25279 11848 25288
rect 11796 25245 11805 25279
rect 11805 25245 11839 25279
rect 11839 25245 11848 25279
rect 11796 25236 11848 25245
rect 12348 25236 12400 25288
rect 14556 25304 14608 25356
rect 15108 25304 15160 25356
rect 11612 25168 11664 25220
rect 12256 25168 12308 25220
rect 15200 25236 15252 25288
rect 16120 25372 16172 25424
rect 16580 25236 16632 25288
rect 17776 25304 17828 25356
rect 20996 25304 21048 25356
rect 8852 25100 8904 25152
rect 11980 25100 12032 25152
rect 13268 25100 13320 25152
rect 13360 25100 13412 25152
rect 14924 25100 14976 25152
rect 15476 25168 15528 25220
rect 15752 25211 15804 25220
rect 15752 25177 15761 25211
rect 15761 25177 15795 25211
rect 15795 25177 15804 25211
rect 17224 25211 17276 25220
rect 15752 25168 15804 25177
rect 16212 25100 16264 25152
rect 17224 25177 17233 25211
rect 17233 25177 17267 25211
rect 17267 25177 17276 25211
rect 17224 25168 17276 25177
rect 18420 25168 18472 25220
rect 19340 25168 19392 25220
rect 20720 25236 20772 25288
rect 20904 25236 20956 25288
rect 21364 25279 21416 25288
rect 21364 25245 21373 25279
rect 21373 25245 21407 25279
rect 21407 25245 21416 25279
rect 21364 25236 21416 25245
rect 22100 25304 22152 25356
rect 22928 25372 22980 25424
rect 22744 25279 22796 25288
rect 20076 25211 20128 25220
rect 20076 25177 20085 25211
rect 20085 25177 20119 25211
rect 20119 25177 20128 25211
rect 20076 25168 20128 25177
rect 20444 25211 20496 25220
rect 20444 25177 20462 25211
rect 20462 25177 20496 25211
rect 22744 25245 22753 25279
rect 22753 25245 22787 25279
rect 22787 25245 22796 25279
rect 22744 25236 22796 25245
rect 20444 25168 20496 25177
rect 22192 25168 22244 25220
rect 23112 25279 23164 25288
rect 23112 25245 23121 25279
rect 23121 25245 23155 25279
rect 23155 25245 23164 25279
rect 23112 25236 23164 25245
rect 24400 25279 24452 25288
rect 24400 25245 24409 25279
rect 24409 25245 24443 25279
rect 24443 25245 24452 25279
rect 24400 25236 24452 25245
rect 24584 25279 24636 25288
rect 24584 25245 24593 25279
rect 24593 25245 24627 25279
rect 24627 25245 24636 25279
rect 24584 25236 24636 25245
rect 26884 25236 26936 25288
rect 27068 25279 27120 25288
rect 27068 25245 27077 25279
rect 27077 25245 27111 25279
rect 27111 25245 27120 25279
rect 27068 25236 27120 25245
rect 25688 25168 25740 25220
rect 26148 25168 26200 25220
rect 18972 25100 19024 25152
rect 20812 25100 20864 25152
rect 23664 25143 23716 25152
rect 23664 25109 23673 25143
rect 23673 25109 23707 25143
rect 23707 25109 23716 25143
rect 23664 25100 23716 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 7932 24896 7984 24948
rect 8668 24896 8720 24948
rect 9128 24939 9180 24948
rect 9128 24905 9137 24939
rect 9137 24905 9171 24939
rect 9171 24905 9180 24939
rect 9128 24896 9180 24905
rect 14464 24896 14516 24948
rect 17960 24896 18012 24948
rect 22560 24896 22612 24948
rect 25504 24939 25556 24948
rect 25504 24905 25513 24939
rect 25513 24905 25547 24939
rect 25547 24905 25556 24939
rect 25504 24896 25556 24905
rect 8392 24760 8444 24812
rect 9956 24828 10008 24880
rect 10416 24871 10468 24880
rect 10416 24837 10425 24871
rect 10425 24837 10459 24871
rect 10459 24837 10468 24871
rect 10416 24828 10468 24837
rect 10140 24803 10192 24812
rect 10140 24769 10149 24803
rect 10149 24769 10183 24803
rect 10183 24769 10192 24803
rect 10140 24760 10192 24769
rect 10600 24760 10652 24812
rect 10692 24760 10744 24812
rect 14832 24828 14884 24880
rect 15752 24828 15804 24880
rect 9220 24735 9272 24744
rect 9220 24701 9229 24735
rect 9229 24701 9263 24735
rect 9263 24701 9272 24735
rect 9220 24692 9272 24701
rect 9404 24735 9456 24744
rect 9404 24701 9413 24735
rect 9413 24701 9447 24735
rect 9447 24701 9456 24735
rect 9404 24692 9456 24701
rect 10048 24692 10100 24744
rect 13452 24760 13504 24812
rect 14556 24760 14608 24812
rect 15200 24760 15252 24812
rect 15844 24760 15896 24812
rect 13728 24692 13780 24744
rect 14004 24735 14056 24744
rect 14004 24701 14013 24735
rect 14013 24701 14047 24735
rect 14047 24701 14056 24735
rect 14004 24692 14056 24701
rect 14648 24692 14700 24744
rect 16212 24760 16264 24812
rect 16948 24803 17000 24812
rect 16948 24769 16957 24803
rect 16957 24769 16991 24803
rect 16991 24769 17000 24803
rect 16948 24760 17000 24769
rect 17684 24760 17736 24812
rect 18788 24803 18840 24812
rect 15108 24624 15160 24676
rect 17776 24692 17828 24744
rect 18788 24769 18797 24803
rect 18797 24769 18831 24803
rect 18831 24769 18840 24803
rect 18788 24760 18840 24769
rect 18972 24803 19024 24812
rect 18972 24769 18981 24803
rect 18981 24769 19015 24803
rect 19015 24769 19024 24803
rect 18972 24760 19024 24769
rect 20904 24803 20956 24812
rect 20904 24769 20913 24803
rect 20913 24769 20947 24803
rect 20947 24769 20956 24803
rect 20904 24760 20956 24769
rect 21272 24828 21324 24880
rect 21456 24760 21508 24812
rect 22468 24803 22520 24812
rect 22468 24769 22477 24803
rect 22477 24769 22511 24803
rect 22511 24769 22520 24803
rect 22468 24760 22520 24769
rect 23664 24828 23716 24880
rect 26516 24828 26568 24880
rect 22744 24760 22796 24812
rect 19432 24692 19484 24744
rect 18420 24624 18472 24676
rect 11520 24556 11572 24608
rect 11612 24556 11664 24608
rect 12808 24556 12860 24608
rect 14556 24556 14608 24608
rect 17132 24556 17184 24608
rect 22192 24735 22244 24744
rect 22192 24701 22201 24735
rect 22201 24701 22235 24735
rect 22235 24701 22244 24735
rect 22192 24692 22244 24701
rect 22284 24692 22336 24744
rect 28356 24760 28408 24812
rect 25964 24735 26016 24744
rect 22652 24624 22704 24676
rect 21548 24556 21600 24608
rect 25964 24701 25973 24735
rect 25973 24701 26007 24735
rect 26007 24701 26016 24735
rect 25964 24692 26016 24701
rect 26148 24735 26200 24744
rect 26148 24701 26157 24735
rect 26157 24701 26191 24735
rect 26191 24701 26200 24735
rect 26148 24692 26200 24701
rect 26240 24624 26292 24676
rect 27436 24624 27488 24676
rect 24676 24556 24728 24608
rect 25044 24599 25096 24608
rect 25044 24565 25053 24599
rect 25053 24565 25087 24599
rect 25087 24565 25096 24599
rect 25044 24556 25096 24565
rect 26976 24556 27028 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 9220 24352 9272 24404
rect 10600 24352 10652 24404
rect 10968 24352 11020 24404
rect 10232 24284 10284 24336
rect 11796 24284 11848 24336
rect 14280 24395 14332 24404
rect 14280 24361 14289 24395
rect 14289 24361 14323 24395
rect 14323 24361 14332 24395
rect 14280 24352 14332 24361
rect 13176 24284 13228 24336
rect 13636 24284 13688 24336
rect 15108 24327 15160 24336
rect 15108 24293 15117 24327
rect 15117 24293 15151 24327
rect 15151 24293 15160 24327
rect 15108 24284 15160 24293
rect 15384 24352 15436 24404
rect 16120 24352 16172 24404
rect 16304 24352 16356 24404
rect 16948 24395 17000 24404
rect 16948 24361 16957 24395
rect 16957 24361 16991 24395
rect 16991 24361 17000 24395
rect 16948 24352 17000 24361
rect 18052 24352 18104 24404
rect 18512 24352 18564 24404
rect 18696 24352 18748 24404
rect 19248 24352 19300 24404
rect 21088 24352 21140 24404
rect 21272 24352 21324 24404
rect 22284 24352 22336 24404
rect 22560 24352 22612 24404
rect 10416 24216 10468 24268
rect 11520 24259 11572 24268
rect 9680 24148 9732 24200
rect 10048 24148 10100 24200
rect 10600 24191 10652 24200
rect 10600 24157 10609 24191
rect 10609 24157 10643 24191
rect 10643 24157 10652 24191
rect 11520 24225 11529 24259
rect 11529 24225 11563 24259
rect 11563 24225 11572 24259
rect 11520 24216 11572 24225
rect 11612 24259 11664 24268
rect 11612 24225 11621 24259
rect 11621 24225 11655 24259
rect 11655 24225 11664 24259
rect 11612 24216 11664 24225
rect 14004 24216 14056 24268
rect 10600 24148 10652 24157
rect 11704 24191 11756 24200
rect 11704 24157 11713 24191
rect 11713 24157 11747 24191
rect 11747 24157 11756 24191
rect 11704 24148 11756 24157
rect 12256 24191 12308 24200
rect 12256 24157 12265 24191
rect 12265 24157 12299 24191
rect 12299 24157 12308 24191
rect 12256 24148 12308 24157
rect 12900 24191 12952 24200
rect 12900 24157 12909 24191
rect 12909 24157 12943 24191
rect 12943 24157 12952 24191
rect 12900 24148 12952 24157
rect 14188 24123 14240 24132
rect 14188 24089 14197 24123
rect 14197 24089 14231 24123
rect 14231 24089 14240 24123
rect 14188 24080 14240 24089
rect 14832 24123 14884 24132
rect 14832 24089 14841 24123
rect 14841 24089 14875 24123
rect 14875 24089 14884 24123
rect 14832 24080 14884 24089
rect 14924 24080 14976 24132
rect 15384 24080 15436 24132
rect 10600 24012 10652 24064
rect 11888 24012 11940 24064
rect 12348 24055 12400 24064
rect 12348 24021 12357 24055
rect 12357 24021 12391 24055
rect 12391 24021 12400 24055
rect 12348 24012 12400 24021
rect 13360 24055 13412 24064
rect 13360 24021 13369 24055
rect 13369 24021 13403 24055
rect 13403 24021 13412 24055
rect 13360 24012 13412 24021
rect 15752 24191 15804 24200
rect 15752 24157 15761 24191
rect 15761 24157 15795 24191
rect 15795 24157 15804 24191
rect 17040 24216 17092 24268
rect 17224 24216 17276 24268
rect 17776 24259 17828 24268
rect 17776 24225 17785 24259
rect 17785 24225 17819 24259
rect 17819 24225 17828 24259
rect 17776 24216 17828 24225
rect 15752 24148 15804 24157
rect 16120 24191 16172 24200
rect 16120 24157 16129 24191
rect 16129 24157 16163 24191
rect 16163 24157 16172 24191
rect 16120 24148 16172 24157
rect 16948 24148 17000 24200
rect 16028 24123 16080 24132
rect 16028 24089 16037 24123
rect 16037 24089 16071 24123
rect 16071 24089 16080 24123
rect 16028 24080 16080 24089
rect 20076 24216 20128 24268
rect 18788 24148 18840 24200
rect 19432 24080 19484 24132
rect 22284 24191 22336 24200
rect 16396 24012 16448 24064
rect 16856 24012 16908 24064
rect 17132 24012 17184 24064
rect 19984 24012 20036 24064
rect 20628 24012 20680 24064
rect 22284 24157 22293 24191
rect 22293 24157 22327 24191
rect 22327 24157 22336 24191
rect 22284 24148 22336 24157
rect 22468 24148 22520 24200
rect 24492 24352 24544 24404
rect 26516 24395 26568 24404
rect 26516 24361 26525 24395
rect 26525 24361 26559 24395
rect 26559 24361 26568 24395
rect 26516 24352 26568 24361
rect 28356 24352 28408 24404
rect 24676 24259 24728 24268
rect 22652 24191 22704 24200
rect 22652 24157 22661 24191
rect 22661 24157 22695 24191
rect 22695 24157 22704 24191
rect 22652 24148 22704 24157
rect 23112 24148 23164 24200
rect 24676 24225 24685 24259
rect 24685 24225 24719 24259
rect 24719 24225 24728 24259
rect 24676 24216 24728 24225
rect 26976 24259 27028 24268
rect 26976 24225 26985 24259
rect 26985 24225 27019 24259
rect 27019 24225 27028 24259
rect 26976 24216 27028 24225
rect 27160 24259 27212 24268
rect 27160 24225 27169 24259
rect 27169 24225 27203 24259
rect 27203 24225 27212 24259
rect 27160 24216 27212 24225
rect 28540 24148 28592 24200
rect 22744 24080 22796 24132
rect 24952 24123 25004 24132
rect 24952 24089 24986 24123
rect 24986 24089 25004 24123
rect 24952 24080 25004 24089
rect 27344 24080 27396 24132
rect 21456 24055 21508 24064
rect 21456 24021 21481 24055
rect 21481 24021 21508 24055
rect 21456 24012 21508 24021
rect 22284 24012 22336 24064
rect 23112 24012 23164 24064
rect 23480 24055 23532 24064
rect 23480 24021 23489 24055
rect 23489 24021 23523 24055
rect 23523 24021 23532 24055
rect 23480 24012 23532 24021
rect 26056 24012 26108 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 7012 23672 7064 23724
rect 10508 23740 10560 23792
rect 8944 23672 8996 23724
rect 10140 23672 10192 23724
rect 11888 23808 11940 23860
rect 11520 23715 11572 23724
rect 9496 23604 9548 23656
rect 9680 23536 9732 23588
rect 11520 23681 11529 23715
rect 11529 23681 11563 23715
rect 11563 23681 11572 23715
rect 11520 23672 11572 23681
rect 11704 23715 11756 23724
rect 11704 23681 11713 23715
rect 11713 23681 11747 23715
rect 11747 23681 11756 23715
rect 11704 23672 11756 23681
rect 12532 23808 12584 23860
rect 13176 23808 13228 23860
rect 13452 23783 13504 23792
rect 13452 23749 13461 23783
rect 13461 23749 13495 23783
rect 13495 23749 13504 23783
rect 13452 23740 13504 23749
rect 15108 23808 15160 23860
rect 16856 23808 16908 23860
rect 15200 23740 15252 23792
rect 15476 23740 15528 23792
rect 15568 23740 15620 23792
rect 15844 23740 15896 23792
rect 18328 23808 18380 23860
rect 18788 23808 18840 23860
rect 21180 23851 21232 23860
rect 21180 23817 21189 23851
rect 21189 23817 21223 23851
rect 21223 23817 21232 23851
rect 21180 23808 21232 23817
rect 21364 23808 21416 23860
rect 24584 23808 24636 23860
rect 25688 23851 25740 23860
rect 25688 23817 25697 23851
rect 25697 23817 25731 23851
rect 25731 23817 25740 23851
rect 25688 23808 25740 23817
rect 25964 23808 26016 23860
rect 28540 23851 28592 23860
rect 28540 23817 28549 23851
rect 28549 23817 28583 23851
rect 28583 23817 28592 23851
rect 28540 23808 28592 23817
rect 17684 23740 17736 23792
rect 24308 23740 24360 23792
rect 11336 23604 11388 23656
rect 8668 23511 8720 23520
rect 8668 23477 8677 23511
rect 8677 23477 8711 23511
rect 8711 23477 8720 23511
rect 8668 23468 8720 23477
rect 9772 23511 9824 23520
rect 9772 23477 9781 23511
rect 9781 23477 9815 23511
rect 9815 23477 9824 23511
rect 9772 23468 9824 23477
rect 9956 23468 10008 23520
rect 10416 23511 10468 23520
rect 10416 23477 10425 23511
rect 10425 23477 10459 23511
rect 10459 23477 10468 23511
rect 10416 23468 10468 23477
rect 11612 23468 11664 23520
rect 12440 23468 12492 23520
rect 12992 23672 13044 23724
rect 13084 23672 13136 23724
rect 13544 23715 13596 23724
rect 13544 23681 13553 23715
rect 13553 23681 13587 23715
rect 13587 23681 13596 23715
rect 13544 23672 13596 23681
rect 14188 23715 14240 23724
rect 14188 23681 14197 23715
rect 14197 23681 14231 23715
rect 14231 23681 14240 23715
rect 14188 23672 14240 23681
rect 12716 23536 12768 23588
rect 13268 23536 13320 23588
rect 13820 23536 13872 23588
rect 14924 23672 14976 23724
rect 16120 23672 16172 23724
rect 16488 23672 16540 23724
rect 21548 23672 21600 23724
rect 22192 23715 22244 23724
rect 22192 23681 22201 23715
rect 22201 23681 22235 23715
rect 22235 23681 22244 23715
rect 22192 23672 22244 23681
rect 22468 23672 22520 23724
rect 23572 23715 23624 23724
rect 15016 23647 15068 23656
rect 15016 23613 15025 23647
rect 15025 23613 15059 23647
rect 15059 23613 15068 23647
rect 15016 23604 15068 23613
rect 13544 23468 13596 23520
rect 14280 23468 14332 23520
rect 15384 23604 15436 23656
rect 15752 23604 15804 23656
rect 17132 23604 17184 23656
rect 17776 23604 17828 23656
rect 22284 23647 22336 23656
rect 22284 23613 22293 23647
rect 22293 23613 22327 23647
rect 22327 23613 22336 23647
rect 22284 23604 22336 23613
rect 22652 23604 22704 23656
rect 23572 23681 23581 23715
rect 23581 23681 23615 23715
rect 23615 23681 23624 23715
rect 23572 23672 23624 23681
rect 23756 23715 23808 23724
rect 23756 23681 23765 23715
rect 23765 23681 23799 23715
rect 23799 23681 23808 23715
rect 23756 23672 23808 23681
rect 25044 23740 25096 23792
rect 26700 23740 26752 23792
rect 27528 23740 27580 23792
rect 24952 23672 25004 23724
rect 27068 23672 27120 23724
rect 27252 23672 27304 23724
rect 28356 23715 28408 23724
rect 28356 23681 28365 23715
rect 28365 23681 28399 23715
rect 28399 23681 28408 23715
rect 28356 23672 28408 23681
rect 29184 23715 29236 23724
rect 29184 23681 29193 23715
rect 29193 23681 29227 23715
rect 29227 23681 29236 23715
rect 29184 23672 29236 23681
rect 29920 23672 29972 23724
rect 23940 23604 23992 23656
rect 24400 23647 24452 23656
rect 24400 23613 24409 23647
rect 24409 23613 24443 23647
rect 24443 23613 24452 23647
rect 24400 23604 24452 23613
rect 27160 23604 27212 23656
rect 26424 23536 26476 23588
rect 27344 23536 27396 23588
rect 28264 23604 28316 23656
rect 15476 23468 15528 23520
rect 16948 23468 17000 23520
rect 24032 23468 24084 23520
rect 29000 23511 29052 23520
rect 29000 23477 29009 23511
rect 29009 23477 29043 23511
rect 29043 23477 29052 23511
rect 29000 23468 29052 23477
rect 29644 23511 29696 23520
rect 29644 23477 29653 23511
rect 29653 23477 29687 23511
rect 29687 23477 29696 23511
rect 29644 23468 29696 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 8116 23264 8168 23316
rect 8944 23307 8996 23316
rect 8944 23273 8953 23307
rect 8953 23273 8987 23307
rect 8987 23273 8996 23307
rect 8944 23264 8996 23273
rect 9404 23264 9456 23316
rect 11152 23264 11204 23316
rect 11336 23307 11388 23316
rect 11336 23273 11345 23307
rect 11345 23273 11379 23307
rect 11379 23273 11388 23307
rect 11336 23264 11388 23273
rect 12532 23264 12584 23316
rect 14832 23264 14884 23316
rect 9220 23196 9272 23248
rect 11520 23196 11572 23248
rect 8944 23128 8996 23180
rect 9128 23128 9180 23180
rect 8668 23060 8720 23112
rect 9496 23128 9548 23180
rect 9404 23103 9456 23112
rect 9404 23069 9413 23103
rect 9413 23069 9447 23103
rect 9447 23069 9456 23103
rect 9404 23060 9456 23069
rect 9588 23103 9640 23112
rect 9588 23069 9597 23103
rect 9597 23069 9631 23103
rect 9631 23069 9640 23103
rect 9588 23060 9640 23069
rect 9772 23060 9824 23112
rect 11612 23103 11664 23112
rect 8852 22992 8904 23044
rect 9036 22992 9088 23044
rect 11612 23069 11621 23103
rect 11621 23069 11655 23103
rect 11655 23069 11664 23103
rect 11612 23060 11664 23069
rect 8668 22924 8720 22976
rect 9312 22924 9364 22976
rect 9588 22924 9640 22976
rect 9772 22924 9824 22976
rect 11888 23060 11940 23112
rect 12256 23196 12308 23248
rect 12624 23196 12676 23248
rect 13912 23196 13964 23248
rect 15660 23264 15712 23316
rect 16304 23264 16356 23316
rect 17224 23264 17276 23316
rect 12440 23128 12492 23180
rect 15568 23128 15620 23180
rect 16120 23171 16172 23180
rect 16120 23137 16129 23171
rect 16129 23137 16163 23171
rect 16163 23137 16172 23171
rect 16120 23128 16172 23137
rect 20076 23264 20128 23316
rect 22192 23264 22244 23316
rect 23296 23264 23348 23316
rect 24768 23196 24820 23248
rect 23112 23171 23164 23180
rect 12624 23103 12676 23112
rect 12624 23069 12633 23103
rect 12633 23069 12667 23103
rect 12667 23069 12676 23103
rect 12624 23060 12676 23069
rect 12900 23060 12952 23112
rect 13176 23060 13228 23112
rect 12532 22992 12584 23044
rect 13268 22992 13320 23044
rect 15108 23060 15160 23112
rect 16396 23103 16448 23112
rect 16396 23069 16430 23103
rect 16430 23069 16448 23103
rect 16396 23060 16448 23069
rect 16856 23060 16908 23112
rect 17776 23060 17828 23112
rect 23112 23137 23121 23171
rect 23121 23137 23155 23171
rect 23155 23137 23164 23171
rect 23112 23128 23164 23137
rect 23756 23128 23808 23180
rect 24952 23307 25004 23316
rect 24952 23273 24961 23307
rect 24961 23273 24995 23307
rect 24995 23273 25004 23307
rect 24952 23264 25004 23273
rect 28356 23264 28408 23316
rect 29184 23264 29236 23316
rect 18328 23103 18380 23112
rect 18328 23069 18337 23103
rect 18337 23069 18371 23103
rect 18371 23069 18380 23103
rect 18328 23060 18380 23069
rect 21180 23060 21232 23112
rect 24032 23060 24084 23112
rect 24492 23060 24544 23112
rect 26424 23128 26476 23180
rect 25596 23103 25648 23112
rect 25596 23069 25605 23103
rect 25605 23069 25639 23103
rect 25639 23069 25648 23103
rect 25596 23060 25648 23069
rect 26240 23060 26292 23112
rect 26976 23128 27028 23180
rect 27436 23128 27488 23180
rect 28080 23060 28132 23112
rect 28264 23103 28316 23112
rect 28264 23069 28273 23103
rect 28273 23069 28307 23103
rect 28307 23069 28316 23103
rect 28264 23060 28316 23069
rect 28448 23103 28500 23112
rect 28448 23069 28457 23103
rect 28457 23069 28491 23103
rect 28491 23069 28500 23103
rect 28448 23060 28500 23069
rect 29000 23060 29052 23112
rect 11796 22924 11848 22976
rect 12348 22924 12400 22976
rect 12808 22924 12860 22976
rect 14004 22924 14056 22976
rect 14832 22924 14884 22976
rect 15016 22924 15068 22976
rect 15476 22924 15528 22976
rect 15568 22924 15620 22976
rect 17132 22924 17184 22976
rect 17868 22924 17920 22976
rect 20720 22992 20772 23044
rect 21088 22992 21140 23044
rect 21916 22992 21968 23044
rect 23572 22992 23624 23044
rect 21364 22924 21416 22976
rect 22100 22924 22152 22976
rect 22560 22924 22612 22976
rect 22928 22967 22980 22976
rect 22928 22933 22937 22967
rect 22937 22933 22971 22967
rect 22971 22933 22980 22967
rect 24676 23035 24728 23044
rect 24676 23001 24685 23035
rect 24685 23001 24719 23035
rect 24719 23001 24728 23035
rect 24676 22992 24728 23001
rect 25412 22967 25464 22976
rect 22928 22924 22980 22933
rect 25412 22933 25421 22967
rect 25421 22933 25455 22967
rect 25455 22933 25464 22967
rect 25412 22924 25464 22933
rect 26424 22924 26476 22976
rect 27620 22992 27672 23044
rect 27528 22924 27580 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 9404 22720 9456 22772
rect 10232 22763 10284 22772
rect 10232 22729 10241 22763
rect 10241 22729 10275 22763
rect 10275 22729 10284 22763
rect 10232 22720 10284 22729
rect 10508 22720 10560 22772
rect 11152 22720 11204 22772
rect 12624 22720 12676 22772
rect 12716 22763 12768 22772
rect 12716 22729 12725 22763
rect 12725 22729 12759 22763
rect 12759 22729 12768 22763
rect 12716 22720 12768 22729
rect 6920 22627 6972 22636
rect 6920 22593 6929 22627
rect 6929 22593 6963 22627
rect 6963 22593 6972 22627
rect 6920 22584 6972 22593
rect 8116 22652 8168 22704
rect 8208 22627 8260 22636
rect 8208 22593 8217 22627
rect 8217 22593 8251 22627
rect 8251 22593 8260 22627
rect 8208 22584 8260 22593
rect 8576 22652 8628 22704
rect 13084 22652 13136 22704
rect 9128 22627 9180 22636
rect 9128 22593 9137 22627
rect 9137 22593 9171 22627
rect 9171 22593 9180 22627
rect 9128 22584 9180 22593
rect 9220 22584 9272 22636
rect 10508 22584 10560 22636
rect 11336 22584 11388 22636
rect 11980 22584 12032 22636
rect 12808 22584 12860 22636
rect 14280 22720 14332 22772
rect 15108 22720 15160 22772
rect 15292 22720 15344 22772
rect 16948 22763 17000 22772
rect 16948 22729 16957 22763
rect 16957 22729 16991 22763
rect 16991 22729 17000 22763
rect 16948 22720 17000 22729
rect 22284 22720 22336 22772
rect 22928 22720 22980 22772
rect 9312 22448 9364 22500
rect 9496 22516 9548 22568
rect 10416 22516 10468 22568
rect 14096 22652 14148 22704
rect 13176 22516 13228 22568
rect 15108 22584 15160 22636
rect 15384 22584 15436 22636
rect 15568 22584 15620 22636
rect 16856 22584 16908 22636
rect 18328 22652 18380 22704
rect 22100 22652 22152 22704
rect 17040 22584 17092 22636
rect 17592 22627 17644 22636
rect 17592 22593 17601 22627
rect 17601 22593 17635 22627
rect 17635 22593 17644 22627
rect 17592 22584 17644 22593
rect 17776 22584 17828 22636
rect 22192 22627 22244 22636
rect 11060 22448 11112 22500
rect 8300 22423 8352 22432
rect 8300 22389 8309 22423
rect 8309 22389 8343 22423
rect 8343 22389 8352 22423
rect 8300 22380 8352 22389
rect 8392 22380 8444 22432
rect 8944 22380 8996 22432
rect 9220 22380 9272 22432
rect 9404 22423 9456 22432
rect 9404 22389 9413 22423
rect 9413 22389 9447 22423
rect 9447 22389 9456 22423
rect 9404 22380 9456 22389
rect 9496 22380 9548 22432
rect 13176 22380 13228 22432
rect 13452 22380 13504 22432
rect 14004 22516 14056 22568
rect 17868 22559 17920 22568
rect 17868 22525 17877 22559
rect 17877 22525 17911 22559
rect 17911 22525 17920 22559
rect 17868 22516 17920 22525
rect 18144 22516 18196 22568
rect 18328 22559 18380 22568
rect 18328 22525 18337 22559
rect 18337 22525 18371 22559
rect 18371 22525 18380 22559
rect 18328 22516 18380 22525
rect 22192 22593 22201 22627
rect 22201 22593 22235 22627
rect 22235 22593 22244 22627
rect 22192 22584 22244 22593
rect 22928 22584 22980 22636
rect 27436 22720 27488 22772
rect 23572 22695 23624 22704
rect 23572 22661 23581 22695
rect 23581 22661 23615 22695
rect 23615 22661 23624 22695
rect 23572 22652 23624 22661
rect 25412 22652 25464 22704
rect 26424 22652 26476 22704
rect 13912 22380 13964 22432
rect 14832 22448 14884 22500
rect 15384 22448 15436 22500
rect 18236 22448 18288 22500
rect 17316 22380 17368 22432
rect 17500 22380 17552 22432
rect 18604 22380 18656 22432
rect 18696 22423 18748 22432
rect 18696 22389 18705 22423
rect 18705 22389 18739 22423
rect 18739 22389 18748 22423
rect 18696 22380 18748 22389
rect 19432 22380 19484 22432
rect 21456 22516 21508 22568
rect 23296 22516 23348 22568
rect 20904 22448 20956 22500
rect 23756 22627 23808 22636
rect 23756 22593 23765 22627
rect 23765 22593 23799 22627
rect 23799 22593 23808 22627
rect 27528 22627 27580 22636
rect 23756 22584 23808 22593
rect 27528 22593 27537 22627
rect 27537 22593 27571 22627
rect 27571 22593 27580 22627
rect 27528 22584 27580 22593
rect 27804 22695 27856 22704
rect 27804 22661 27813 22695
rect 27813 22661 27847 22695
rect 27847 22661 27856 22695
rect 27804 22652 27856 22661
rect 24492 22559 24544 22568
rect 24492 22525 24501 22559
rect 24501 22525 24535 22559
rect 24535 22525 24544 22559
rect 24492 22516 24544 22525
rect 28448 22720 28500 22772
rect 29644 22652 29696 22704
rect 28080 22448 28132 22500
rect 21088 22380 21140 22432
rect 24124 22380 24176 22432
rect 26700 22380 26752 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 6920 22176 6972 22228
rect 9128 22176 9180 22228
rect 12808 22176 12860 22228
rect 13544 22176 13596 22228
rect 8208 22108 8260 22160
rect 11060 22108 11112 22160
rect 8300 22040 8352 22092
rect 7932 21904 7984 21956
rect 8576 21904 8628 21956
rect 8208 21836 8260 21888
rect 9312 22040 9364 22092
rect 9496 22040 9548 22092
rect 9680 22040 9732 22092
rect 9128 21972 9180 22024
rect 10508 21972 10560 22024
rect 11060 22015 11112 22024
rect 11060 21981 11069 22015
rect 11069 21981 11103 22015
rect 11103 21981 11112 22015
rect 11060 21972 11112 21981
rect 14832 22176 14884 22228
rect 15384 22176 15436 22228
rect 15936 22176 15988 22228
rect 13912 22108 13964 22160
rect 14188 22108 14240 22160
rect 12900 22040 12952 22092
rect 13544 22083 13596 22092
rect 13544 22049 13553 22083
rect 13553 22049 13587 22083
rect 13587 22049 13596 22083
rect 13544 22040 13596 22049
rect 11428 21972 11480 22024
rect 11520 21972 11572 22024
rect 11888 21972 11940 22024
rect 12348 21972 12400 22024
rect 12532 22015 12584 22024
rect 12532 21981 12541 22015
rect 12541 21981 12575 22015
rect 12575 21981 12584 22015
rect 12716 22015 12768 22024
rect 12532 21972 12584 21981
rect 12716 21981 12725 22015
rect 12725 21981 12759 22015
rect 12759 21981 12768 22015
rect 12716 21972 12768 21981
rect 12808 22015 12860 22024
rect 12808 21981 12817 22015
rect 12817 21981 12851 22015
rect 12851 21981 12860 22015
rect 12808 21972 12860 21981
rect 13360 21972 13412 22024
rect 14924 22015 14976 22024
rect 9588 21904 9640 21956
rect 9496 21836 9548 21888
rect 10784 21836 10836 21888
rect 12072 21904 12124 21956
rect 12624 21836 12676 21888
rect 13452 21836 13504 21888
rect 14924 21981 14933 22015
rect 14933 21981 14967 22015
rect 14967 21981 14976 22015
rect 14924 21972 14976 21981
rect 18236 22108 18288 22160
rect 21456 22176 21508 22228
rect 28264 22176 28316 22228
rect 28632 22176 28684 22228
rect 20720 22108 20772 22160
rect 18604 22040 18656 22092
rect 22468 22108 22520 22160
rect 21548 22083 21600 22092
rect 21548 22049 21557 22083
rect 21557 22049 21591 22083
rect 21591 22049 21600 22083
rect 21548 22040 21600 22049
rect 17224 22015 17276 22024
rect 17224 21981 17233 22015
rect 17233 21981 17267 22015
rect 17267 21981 17276 22015
rect 17224 21972 17276 21981
rect 17500 22015 17552 22024
rect 17500 21981 17534 22015
rect 17534 21981 17552 22015
rect 17500 21972 17552 21981
rect 20168 21972 20220 22024
rect 20352 21972 20404 22024
rect 20812 22015 20864 22024
rect 20812 21981 20821 22015
rect 20821 21981 20855 22015
rect 20855 21981 20864 22015
rect 20812 21972 20864 21981
rect 17316 21904 17368 21956
rect 21824 21972 21876 22024
rect 22100 22015 22152 22024
rect 22100 21981 22110 22015
rect 22110 21981 22144 22015
rect 22144 21981 22152 22015
rect 22100 21972 22152 21981
rect 22468 22015 22520 22024
rect 22468 21981 22482 22015
rect 22482 21981 22516 22015
rect 22516 21981 22520 22015
rect 22468 21972 22520 21981
rect 22928 21972 22980 22024
rect 21364 21947 21416 21956
rect 21364 21913 21373 21947
rect 21373 21913 21407 21947
rect 21407 21913 21416 21947
rect 21364 21904 21416 21913
rect 22284 21947 22336 21956
rect 22284 21913 22293 21947
rect 22293 21913 22327 21947
rect 22327 21913 22336 21947
rect 22284 21904 22336 21913
rect 14188 21879 14240 21888
rect 14188 21845 14197 21879
rect 14197 21845 14231 21879
rect 14231 21845 14240 21879
rect 14188 21836 14240 21845
rect 15384 21836 15436 21888
rect 22100 21836 22152 21888
rect 22652 21879 22704 21888
rect 22652 21845 22661 21879
rect 22661 21845 22695 21879
rect 22695 21845 22704 21879
rect 22652 21836 22704 21845
rect 22836 21904 22888 21956
rect 23756 21972 23808 22024
rect 24676 22015 24728 22024
rect 24676 21981 24685 22015
rect 24685 21981 24719 22015
rect 24719 21981 24728 22015
rect 24676 21972 24728 21981
rect 26700 21972 26752 22024
rect 28080 22040 28132 22092
rect 28632 22040 28684 22092
rect 29920 22083 29972 22092
rect 29920 22049 29929 22083
rect 29929 22049 29963 22083
rect 29963 22049 29972 22083
rect 29920 22040 29972 22049
rect 28724 22015 28776 22024
rect 28724 21981 28733 22015
rect 28733 21981 28767 22015
rect 28767 21981 28776 22015
rect 28724 21972 28776 21981
rect 24400 21904 24452 21956
rect 26240 21904 26292 21956
rect 23020 21836 23072 21888
rect 23664 21879 23716 21888
rect 23664 21845 23673 21879
rect 23673 21845 23707 21879
rect 23707 21845 23716 21879
rect 23664 21836 23716 21845
rect 27896 21836 27948 21888
rect 27988 21836 28040 21888
rect 28356 21836 28408 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 9220 21632 9272 21684
rect 9496 21632 9548 21684
rect 11704 21675 11756 21684
rect 11704 21641 11713 21675
rect 11713 21641 11747 21675
rect 11747 21641 11756 21675
rect 11704 21632 11756 21641
rect 7748 21539 7800 21548
rect 7748 21505 7757 21539
rect 7757 21505 7791 21539
rect 7791 21505 7800 21539
rect 7748 21496 7800 21505
rect 7932 21539 7984 21548
rect 7932 21505 7941 21539
rect 7941 21505 7975 21539
rect 7975 21505 7984 21539
rect 7932 21496 7984 21505
rect 8484 21496 8536 21548
rect 12348 21564 12400 21616
rect 13912 21632 13964 21684
rect 14832 21632 14884 21684
rect 15200 21632 15252 21684
rect 15384 21632 15436 21684
rect 16488 21632 16540 21684
rect 17316 21675 17368 21684
rect 17316 21641 17325 21675
rect 17325 21641 17359 21675
rect 17359 21641 17368 21675
rect 17316 21632 17368 21641
rect 17592 21632 17644 21684
rect 20812 21632 20864 21684
rect 25596 21632 25648 21684
rect 26884 21632 26936 21684
rect 8024 21471 8076 21480
rect 8024 21437 8033 21471
rect 8033 21437 8067 21471
rect 8067 21437 8076 21471
rect 8024 21428 8076 21437
rect 9404 21539 9456 21548
rect 9404 21505 9413 21539
rect 9413 21505 9447 21539
rect 9447 21505 9456 21539
rect 9404 21496 9456 21505
rect 9588 21539 9640 21548
rect 9588 21505 9597 21539
rect 9597 21505 9631 21539
rect 9631 21505 9640 21539
rect 9588 21496 9640 21505
rect 11060 21496 11112 21548
rect 11888 21496 11940 21548
rect 12072 21496 12124 21548
rect 13268 21539 13320 21548
rect 13268 21505 13277 21539
rect 13277 21505 13311 21539
rect 13311 21505 13320 21539
rect 13268 21496 13320 21505
rect 13544 21496 13596 21548
rect 10692 21471 10744 21480
rect 10692 21437 10701 21471
rect 10701 21437 10735 21471
rect 10735 21437 10744 21471
rect 10692 21428 10744 21437
rect 11336 21428 11388 21480
rect 12164 21471 12216 21480
rect 12164 21437 12173 21471
rect 12173 21437 12207 21471
rect 12207 21437 12216 21471
rect 12164 21428 12216 21437
rect 10416 21360 10468 21412
rect 11980 21360 12032 21412
rect 12348 21360 12400 21412
rect 13820 21496 13872 21548
rect 14832 21496 14884 21548
rect 15292 21564 15344 21616
rect 16028 21564 16080 21616
rect 18696 21564 18748 21616
rect 21548 21564 21600 21616
rect 21640 21564 21692 21616
rect 22928 21564 22980 21616
rect 23756 21564 23808 21616
rect 15844 21496 15896 21548
rect 16856 21496 16908 21548
rect 17316 21496 17368 21548
rect 19340 21539 19392 21548
rect 19340 21505 19374 21539
rect 19374 21505 19392 21539
rect 21824 21539 21876 21548
rect 19340 21496 19392 21505
rect 21824 21505 21833 21539
rect 21833 21505 21867 21539
rect 21867 21505 21876 21539
rect 21824 21496 21876 21505
rect 15384 21428 15436 21480
rect 22100 21539 22152 21548
rect 22100 21505 22109 21539
rect 22109 21505 22143 21539
rect 22143 21505 22152 21539
rect 22100 21496 22152 21505
rect 22468 21496 22520 21548
rect 23664 21496 23716 21548
rect 23940 21539 23992 21548
rect 23940 21505 23949 21539
rect 23949 21505 23983 21539
rect 23983 21505 23992 21539
rect 23940 21496 23992 21505
rect 24124 21539 24176 21548
rect 24124 21505 24133 21539
rect 24133 21505 24167 21539
rect 24167 21505 24176 21539
rect 24124 21496 24176 21505
rect 24676 21564 24728 21616
rect 26240 21607 26292 21616
rect 26240 21573 26249 21607
rect 26249 21573 26283 21607
rect 26283 21573 26292 21607
rect 26240 21564 26292 21573
rect 27160 21496 27212 21548
rect 27712 21496 27764 21548
rect 28356 21539 28408 21548
rect 15568 21360 15620 21412
rect 16580 21360 16632 21412
rect 8300 21292 8352 21344
rect 8944 21335 8996 21344
rect 8944 21301 8953 21335
rect 8953 21301 8987 21335
rect 8987 21301 8996 21335
rect 8944 21292 8996 21301
rect 9036 21292 9088 21344
rect 9588 21292 9640 21344
rect 10140 21292 10192 21344
rect 10784 21292 10836 21344
rect 12164 21292 12216 21344
rect 12900 21292 12952 21344
rect 14924 21292 14976 21344
rect 22560 21428 22612 21480
rect 22836 21428 22888 21480
rect 23664 21360 23716 21412
rect 27344 21360 27396 21412
rect 19984 21292 20036 21344
rect 20536 21292 20588 21344
rect 22008 21292 22060 21344
rect 22468 21335 22520 21344
rect 22468 21301 22477 21335
rect 22477 21301 22511 21335
rect 22511 21301 22520 21335
rect 22468 21292 22520 21301
rect 24400 21292 24452 21344
rect 26884 21292 26936 21344
rect 28356 21505 28365 21539
rect 28365 21505 28399 21539
rect 28399 21505 28408 21539
rect 28356 21496 28408 21505
rect 28816 21471 28868 21480
rect 28816 21437 28825 21471
rect 28825 21437 28859 21471
rect 28859 21437 28868 21471
rect 28816 21428 28868 21437
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 8024 21088 8076 21140
rect 8484 21088 8536 21140
rect 8668 20952 8720 21004
rect 9128 20952 9180 21004
rect 11060 21088 11112 21140
rect 19340 21088 19392 21140
rect 22192 21088 22244 21140
rect 25872 21088 25924 21140
rect 27068 21131 27120 21140
rect 27068 21097 27077 21131
rect 27077 21097 27111 21131
rect 27111 21097 27120 21131
rect 27068 21088 27120 21097
rect 28724 21088 28776 21140
rect 10416 20952 10468 21004
rect 12348 20952 12400 21004
rect 8392 20884 8444 20936
rect 10508 20927 10560 20936
rect 10508 20893 10517 20927
rect 10517 20893 10551 20927
rect 10551 20893 10560 20927
rect 10508 20884 10560 20893
rect 11152 20884 11204 20936
rect 13728 20952 13780 21004
rect 19340 20952 19392 21004
rect 23664 21020 23716 21072
rect 12900 20927 12952 20936
rect 12900 20893 12909 20927
rect 12909 20893 12943 20927
rect 12943 20893 12952 20927
rect 13360 20927 13412 20936
rect 12900 20884 12952 20893
rect 13360 20893 13369 20927
rect 13369 20893 13403 20927
rect 13403 20893 13412 20927
rect 13360 20884 13412 20893
rect 16580 20884 16632 20936
rect 19432 20927 19484 20936
rect 19432 20893 19441 20927
rect 19441 20893 19475 20927
rect 19475 20893 19484 20927
rect 19432 20884 19484 20893
rect 11980 20816 12032 20868
rect 8576 20748 8628 20800
rect 12624 20859 12676 20868
rect 12624 20825 12633 20859
rect 12633 20825 12667 20859
rect 12667 20825 12676 20859
rect 12624 20816 12676 20825
rect 14188 20816 14240 20868
rect 14832 20859 14884 20868
rect 14832 20825 14866 20859
rect 14866 20825 14884 20859
rect 17132 20859 17184 20868
rect 14832 20816 14884 20825
rect 17132 20825 17166 20859
rect 17166 20825 17184 20859
rect 17132 20816 17184 20825
rect 17224 20816 17276 20868
rect 16304 20748 16356 20800
rect 17408 20748 17460 20800
rect 19984 20884 20036 20936
rect 20812 20884 20864 20936
rect 21824 20884 21876 20936
rect 22008 20927 22060 20936
rect 22008 20893 22017 20927
rect 22017 20893 22051 20927
rect 22051 20893 22060 20927
rect 22008 20884 22060 20893
rect 22928 20884 22980 20936
rect 23204 20927 23256 20936
rect 23204 20893 23213 20927
rect 23213 20893 23247 20927
rect 23247 20893 23256 20927
rect 23204 20884 23256 20893
rect 23388 20927 23440 20936
rect 23388 20893 23395 20927
rect 23395 20893 23440 20927
rect 23388 20884 23440 20893
rect 20536 20748 20588 20800
rect 20720 20748 20772 20800
rect 22284 20859 22336 20868
rect 22284 20825 22293 20859
rect 22293 20825 22327 20859
rect 22327 20825 22336 20859
rect 23756 20884 23808 20936
rect 24400 20927 24452 20936
rect 24400 20893 24409 20927
rect 24409 20893 24443 20927
rect 24443 20893 24452 20927
rect 24400 20884 24452 20893
rect 27988 20952 28040 21004
rect 28356 20952 28408 21004
rect 25136 20884 25188 20936
rect 27712 20927 27764 20936
rect 27712 20893 27721 20927
rect 27721 20893 27755 20927
rect 27755 20893 27764 20927
rect 27712 20884 27764 20893
rect 27896 20927 27948 20936
rect 27896 20893 27905 20927
rect 27905 20893 27939 20927
rect 27939 20893 27948 20927
rect 27896 20884 27948 20893
rect 28080 20927 28132 20936
rect 28080 20893 28089 20927
rect 28089 20893 28123 20927
rect 28123 20893 28132 20927
rect 28080 20884 28132 20893
rect 22284 20816 22336 20825
rect 23572 20859 23624 20868
rect 23572 20825 23581 20859
rect 23581 20825 23615 20859
rect 23615 20825 23624 20859
rect 23572 20816 23624 20825
rect 26240 20816 26292 20868
rect 26792 20816 26844 20868
rect 27528 20816 27580 20868
rect 27988 20859 28040 20868
rect 27988 20825 27997 20859
rect 27997 20825 28031 20859
rect 28031 20825 28040 20859
rect 27988 20816 28040 20825
rect 23940 20748 23992 20800
rect 27436 20748 27488 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 9128 20544 9180 20596
rect 10508 20544 10560 20596
rect 10600 20544 10652 20596
rect 8944 20476 8996 20528
rect 9404 20476 9456 20528
rect 12256 20544 12308 20596
rect 12348 20587 12400 20596
rect 12348 20553 12357 20587
rect 12357 20553 12391 20587
rect 12391 20553 12400 20587
rect 13084 20587 13136 20596
rect 12348 20544 12400 20553
rect 13084 20553 13093 20587
rect 13093 20553 13127 20587
rect 13127 20553 13136 20587
rect 13084 20544 13136 20553
rect 15568 20587 15620 20596
rect 15568 20553 15577 20587
rect 15577 20553 15611 20587
rect 15611 20553 15620 20587
rect 15568 20544 15620 20553
rect 17132 20587 17184 20596
rect 17132 20553 17141 20587
rect 17141 20553 17175 20587
rect 17175 20553 17184 20587
rect 17132 20544 17184 20553
rect 11796 20519 11848 20528
rect 11796 20485 11805 20519
rect 11805 20485 11839 20519
rect 11839 20485 11848 20519
rect 11796 20476 11848 20485
rect 8300 20408 8352 20460
rect 8484 20451 8536 20460
rect 8484 20417 8493 20451
rect 8493 20417 8527 20451
rect 8527 20417 8536 20451
rect 8484 20408 8536 20417
rect 10232 20408 10284 20460
rect 10784 20451 10836 20460
rect 10784 20417 10793 20451
rect 10793 20417 10827 20451
rect 10827 20417 10836 20451
rect 10784 20408 10836 20417
rect 10876 20451 10928 20460
rect 10876 20417 10885 20451
rect 10885 20417 10919 20451
rect 10919 20417 10928 20451
rect 10876 20408 10928 20417
rect 11888 20408 11940 20460
rect 12716 20476 12768 20528
rect 15476 20476 15528 20528
rect 12992 20451 13044 20460
rect 12992 20417 13001 20451
rect 13001 20417 13035 20451
rect 13035 20417 13044 20451
rect 12992 20408 13044 20417
rect 9496 20340 9548 20392
rect 16764 20408 16816 20460
rect 17040 20408 17092 20460
rect 17408 20451 17460 20460
rect 17408 20417 17417 20451
rect 17417 20417 17451 20451
rect 17451 20417 17460 20451
rect 17408 20408 17460 20417
rect 14096 20340 14148 20392
rect 17592 20451 17644 20460
rect 17592 20417 17601 20451
rect 17601 20417 17635 20451
rect 17635 20417 17644 20451
rect 17592 20408 17644 20417
rect 18696 20408 18748 20460
rect 20812 20544 20864 20596
rect 22192 20544 22244 20596
rect 23204 20544 23256 20596
rect 23480 20544 23532 20596
rect 25136 20544 25188 20596
rect 19984 20476 20036 20528
rect 22468 20476 22520 20528
rect 26884 20544 26936 20596
rect 11060 20272 11112 20324
rect 11980 20247 12032 20256
rect 11980 20213 11989 20247
rect 11989 20213 12023 20247
rect 12023 20213 12032 20247
rect 11980 20204 12032 20213
rect 17500 20272 17552 20324
rect 12348 20204 12400 20256
rect 13452 20204 13504 20256
rect 15476 20204 15528 20256
rect 19156 20340 19208 20392
rect 21180 20408 21232 20460
rect 21548 20408 21600 20460
rect 23664 20451 23716 20460
rect 23664 20417 23673 20451
rect 23673 20417 23707 20451
rect 23707 20417 23716 20451
rect 23664 20408 23716 20417
rect 23940 20451 23992 20460
rect 23940 20417 23974 20451
rect 23974 20417 23992 20451
rect 23940 20408 23992 20417
rect 25688 20451 25740 20460
rect 25688 20417 25695 20451
rect 25695 20417 25740 20451
rect 25688 20408 25740 20417
rect 26884 20408 26936 20460
rect 27344 20544 27396 20596
rect 27528 20476 27580 20528
rect 22836 20272 22888 20324
rect 25872 20272 25924 20324
rect 25964 20272 26016 20324
rect 27436 20451 27488 20460
rect 27436 20417 27450 20451
rect 27450 20417 27484 20451
rect 27484 20417 27488 20451
rect 27436 20408 27488 20417
rect 28356 20340 28408 20392
rect 27252 20272 27304 20324
rect 27528 20272 27580 20324
rect 18144 20204 18196 20256
rect 19248 20204 19300 20256
rect 20536 20204 20588 20256
rect 20812 20204 20864 20256
rect 26148 20247 26200 20256
rect 26148 20213 26157 20247
rect 26157 20213 26191 20247
rect 26191 20213 26200 20247
rect 26148 20204 26200 20213
rect 27620 20247 27672 20256
rect 27620 20213 27629 20247
rect 27629 20213 27663 20247
rect 27663 20213 27672 20247
rect 27620 20204 27672 20213
rect 28816 20272 28868 20324
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 9496 20000 9548 20052
rect 10692 20000 10744 20052
rect 10784 20000 10836 20052
rect 9956 19932 10008 19984
rect 11704 20000 11756 20052
rect 13176 20043 13228 20052
rect 13176 20009 13185 20043
rect 13185 20009 13219 20043
rect 13219 20009 13228 20043
rect 13176 20000 13228 20009
rect 14832 20000 14884 20052
rect 9496 19839 9548 19848
rect 9496 19805 9505 19839
rect 9505 19805 9539 19839
rect 9539 19805 9548 19839
rect 9496 19796 9548 19805
rect 10140 19839 10192 19848
rect 10140 19805 10149 19839
rect 10149 19805 10183 19839
rect 10183 19805 10192 19839
rect 10140 19796 10192 19805
rect 10600 19796 10652 19848
rect 11060 19796 11112 19848
rect 10692 19728 10744 19780
rect 11796 19796 11848 19848
rect 13360 19932 13412 19984
rect 13728 19932 13780 19984
rect 13452 19796 13504 19848
rect 12256 19728 12308 19780
rect 17408 20000 17460 20052
rect 17592 20000 17644 20052
rect 18696 20043 18748 20052
rect 18696 20009 18705 20043
rect 18705 20009 18739 20043
rect 18739 20009 18748 20043
rect 18696 20000 18748 20009
rect 19432 20000 19484 20052
rect 20536 20000 20588 20052
rect 22744 20000 22796 20052
rect 25688 20000 25740 20052
rect 26056 20000 26108 20052
rect 26792 20043 26844 20052
rect 26792 20009 26801 20043
rect 26801 20009 26835 20043
rect 26835 20009 26844 20043
rect 26792 20000 26844 20009
rect 27252 20000 27304 20052
rect 15016 19932 15068 19984
rect 16304 19932 16356 19984
rect 18972 19932 19024 19984
rect 9588 19660 9640 19712
rect 12716 19660 12768 19712
rect 15476 19796 15528 19848
rect 16396 19796 16448 19848
rect 18144 19839 18196 19848
rect 17592 19728 17644 19780
rect 17868 19728 17920 19780
rect 18144 19805 18153 19839
rect 18153 19805 18187 19839
rect 18187 19805 18196 19839
rect 18144 19796 18196 19805
rect 19616 19932 19668 19984
rect 19708 19864 19760 19916
rect 18512 19839 18564 19848
rect 18512 19805 18521 19839
rect 18521 19805 18555 19839
rect 18555 19805 18564 19839
rect 18512 19796 18564 19805
rect 19340 19796 19392 19848
rect 19616 19839 19668 19848
rect 19616 19805 19625 19839
rect 19625 19805 19659 19839
rect 19659 19805 19668 19839
rect 20260 19932 20312 19984
rect 21548 19907 21600 19916
rect 21548 19873 21557 19907
rect 21557 19873 21591 19907
rect 21591 19873 21600 19907
rect 21548 19864 21600 19873
rect 24492 19864 24544 19916
rect 19616 19796 19668 19805
rect 20628 19839 20680 19848
rect 20628 19805 20637 19839
rect 20637 19805 20671 19839
rect 20671 19805 20680 19839
rect 20628 19796 20680 19805
rect 20904 19839 20956 19848
rect 20904 19805 20913 19839
rect 20913 19805 20947 19839
rect 20947 19805 20956 19839
rect 20904 19796 20956 19805
rect 21180 19796 21232 19848
rect 22652 19796 22704 19848
rect 26148 19796 26200 19848
rect 26976 19796 27028 19848
rect 27528 19796 27580 19848
rect 26700 19771 26752 19780
rect 26700 19737 26709 19771
rect 26709 19737 26743 19771
rect 26743 19737 26752 19771
rect 26700 19728 26752 19737
rect 27620 19728 27672 19780
rect 15752 19660 15804 19712
rect 19432 19660 19484 19712
rect 20260 19660 20312 19712
rect 20444 19703 20496 19712
rect 20444 19669 20453 19703
rect 20453 19669 20487 19703
rect 20487 19669 20496 19703
rect 20444 19660 20496 19669
rect 27252 19660 27304 19712
rect 27712 19660 27764 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 9772 19456 9824 19508
rect 12532 19456 12584 19508
rect 14372 19456 14424 19508
rect 10232 19320 10284 19372
rect 10508 19388 10560 19440
rect 10876 19388 10928 19440
rect 11796 19388 11848 19440
rect 13084 19388 13136 19440
rect 14924 19431 14976 19440
rect 14924 19397 14933 19431
rect 14933 19397 14967 19431
rect 14967 19397 14976 19431
rect 14924 19388 14976 19397
rect 15476 19388 15528 19440
rect 15660 19388 15712 19440
rect 10600 19363 10652 19372
rect 10600 19329 10609 19363
rect 10609 19329 10643 19363
rect 10643 19329 10652 19363
rect 10600 19320 10652 19329
rect 10692 19320 10744 19372
rect 11520 19363 11572 19372
rect 10968 19295 11020 19304
rect 10968 19261 10977 19295
rect 10977 19261 11011 19295
rect 11011 19261 11020 19295
rect 10968 19252 11020 19261
rect 11520 19329 11529 19363
rect 11529 19329 11563 19363
rect 11563 19329 11572 19363
rect 11520 19320 11572 19329
rect 15752 19363 15804 19372
rect 15752 19329 15761 19363
rect 15761 19329 15795 19363
rect 15795 19329 15804 19363
rect 15752 19320 15804 19329
rect 15844 19363 15896 19372
rect 15844 19329 15853 19363
rect 15853 19329 15887 19363
rect 15887 19329 15896 19363
rect 17316 19388 17368 19440
rect 17592 19388 17644 19440
rect 18144 19388 18196 19440
rect 15844 19320 15896 19329
rect 16396 19320 16448 19372
rect 17868 19363 17920 19372
rect 17868 19329 17877 19363
rect 17877 19329 17911 19363
rect 17911 19329 17920 19363
rect 17868 19320 17920 19329
rect 19340 19320 19392 19372
rect 16028 19252 16080 19304
rect 18696 19252 18748 19304
rect 19156 19295 19208 19304
rect 8484 19184 8536 19236
rect 14096 19184 14148 19236
rect 19156 19261 19165 19295
rect 19165 19261 19199 19295
rect 19199 19261 19208 19295
rect 19156 19252 19208 19261
rect 20996 19320 21048 19372
rect 21732 19320 21784 19372
rect 21916 19363 21968 19372
rect 21916 19329 21925 19363
rect 21925 19329 21959 19363
rect 21959 19329 21968 19363
rect 21916 19320 21968 19329
rect 22100 19363 22152 19372
rect 22100 19329 22109 19363
rect 22109 19329 22143 19363
rect 22143 19329 22152 19363
rect 22100 19320 22152 19329
rect 23020 19456 23072 19508
rect 26240 19456 26292 19508
rect 27160 19456 27212 19508
rect 22376 19320 22428 19372
rect 23204 19320 23256 19372
rect 25780 19363 25832 19372
rect 25780 19329 25790 19363
rect 25790 19329 25824 19363
rect 25824 19329 25832 19363
rect 25780 19320 25832 19329
rect 26056 19363 26108 19372
rect 26056 19329 26085 19363
rect 26085 19329 26108 19363
rect 26056 19320 26108 19329
rect 26240 19320 26292 19372
rect 26976 19320 27028 19372
rect 27712 19320 27764 19372
rect 9772 19159 9824 19168
rect 9772 19125 9781 19159
rect 9781 19125 9815 19159
rect 9815 19125 9824 19159
rect 9772 19116 9824 19125
rect 10600 19116 10652 19168
rect 13544 19159 13596 19168
rect 13544 19125 13553 19159
rect 13553 19125 13587 19159
rect 13587 19125 13596 19159
rect 13544 19116 13596 19125
rect 14464 19116 14516 19168
rect 15108 19116 15160 19168
rect 21916 19184 21968 19236
rect 22192 19184 22244 19236
rect 22468 19184 22520 19236
rect 18144 19116 18196 19168
rect 19064 19116 19116 19168
rect 20168 19116 20220 19168
rect 21732 19116 21784 19168
rect 22376 19116 22428 19168
rect 23388 19116 23440 19168
rect 24952 19116 25004 19168
rect 27344 19252 27396 19304
rect 26240 19116 26292 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 9772 18912 9824 18964
rect 10232 18912 10284 18964
rect 10784 18912 10836 18964
rect 11520 18912 11572 18964
rect 12164 18912 12216 18964
rect 14372 18912 14424 18964
rect 17684 18955 17736 18964
rect 10416 18751 10468 18760
rect 10416 18717 10425 18751
rect 10425 18717 10459 18751
rect 10459 18717 10468 18751
rect 10416 18708 10468 18717
rect 10508 18708 10560 18760
rect 10600 18640 10652 18692
rect 13084 18751 13136 18760
rect 13084 18717 13093 18751
rect 13093 18717 13127 18751
rect 13127 18717 13136 18751
rect 13084 18708 13136 18717
rect 13820 18776 13872 18828
rect 10876 18640 10928 18692
rect 14372 18708 14424 18760
rect 14924 18844 14976 18896
rect 15476 18776 15528 18828
rect 16580 18776 16632 18828
rect 14924 18751 14976 18760
rect 14924 18717 14933 18751
rect 14933 18717 14967 18751
rect 14967 18717 14976 18751
rect 14924 18708 14976 18717
rect 15292 18708 15344 18760
rect 15844 18708 15896 18760
rect 16028 18751 16080 18760
rect 16028 18717 16037 18751
rect 16037 18717 16071 18751
rect 16071 18717 16080 18751
rect 16028 18708 16080 18717
rect 16856 18751 16908 18760
rect 16856 18717 16865 18751
rect 16865 18717 16899 18751
rect 16899 18717 16908 18751
rect 16856 18708 16908 18717
rect 17132 18776 17184 18828
rect 17684 18921 17693 18955
rect 17693 18921 17727 18955
rect 17727 18921 17736 18955
rect 17684 18912 17736 18921
rect 17868 18912 17920 18964
rect 20536 18844 20588 18896
rect 21364 18912 21416 18964
rect 26700 18912 26752 18964
rect 27712 18912 27764 18964
rect 22284 18844 22336 18896
rect 27804 18844 27856 18896
rect 18512 18776 18564 18828
rect 19984 18776 20036 18828
rect 22468 18819 22520 18828
rect 22468 18785 22477 18819
rect 22477 18785 22511 18819
rect 22511 18785 22520 18819
rect 22468 18776 22520 18785
rect 26424 18776 26476 18828
rect 18144 18751 18196 18760
rect 18144 18717 18153 18751
rect 18153 18717 18187 18751
rect 18187 18717 18196 18751
rect 18144 18708 18196 18717
rect 18328 18751 18380 18760
rect 18328 18717 18337 18751
rect 18337 18717 18371 18751
rect 18371 18717 18380 18751
rect 18328 18708 18380 18717
rect 19156 18708 19208 18760
rect 22560 18708 22612 18760
rect 23940 18708 23992 18760
rect 24492 18751 24544 18760
rect 24492 18717 24501 18751
rect 24501 18717 24535 18751
rect 24535 18717 24544 18751
rect 24492 18708 24544 18717
rect 26240 18708 26292 18760
rect 26884 18708 26936 18760
rect 27160 18751 27212 18760
rect 27160 18717 27167 18751
rect 27167 18717 27212 18751
rect 27160 18708 27212 18717
rect 27436 18751 27488 18760
rect 27436 18717 27450 18751
rect 27450 18717 27484 18751
rect 27484 18717 27488 18751
rect 27436 18708 27488 18717
rect 15200 18640 15252 18692
rect 17132 18640 17184 18692
rect 18512 18640 18564 18692
rect 19432 18640 19484 18692
rect 21824 18640 21876 18692
rect 25780 18640 25832 18692
rect 12808 18615 12860 18624
rect 12808 18581 12817 18615
rect 12817 18581 12851 18615
rect 12851 18581 12860 18615
rect 12808 18572 12860 18581
rect 14372 18572 14424 18624
rect 16580 18615 16632 18624
rect 16580 18581 16589 18615
rect 16589 18581 16623 18615
rect 16623 18581 16632 18615
rect 16580 18572 16632 18581
rect 16948 18572 17000 18624
rect 17316 18572 17368 18624
rect 23664 18572 23716 18624
rect 23848 18615 23900 18624
rect 23848 18581 23857 18615
rect 23857 18581 23891 18615
rect 23891 18581 23900 18615
rect 23848 18572 23900 18581
rect 26240 18572 26292 18624
rect 27160 18572 27212 18624
rect 27896 18640 27948 18692
rect 28540 18751 28592 18760
rect 28540 18717 28549 18751
rect 28549 18717 28583 18751
rect 28583 18717 28592 18751
rect 28540 18708 28592 18717
rect 28632 18640 28684 18692
rect 27436 18572 27488 18624
rect 28080 18615 28132 18624
rect 28080 18581 28089 18615
rect 28089 18581 28123 18615
rect 28123 18581 28132 18615
rect 28080 18572 28132 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 10508 18368 10560 18420
rect 10692 18411 10744 18420
rect 10692 18377 10701 18411
rect 10701 18377 10735 18411
rect 10735 18377 10744 18411
rect 10692 18368 10744 18377
rect 13084 18368 13136 18420
rect 16580 18300 16632 18352
rect 8484 18232 8536 18284
rect 10968 18232 11020 18284
rect 13084 18275 13136 18284
rect 13084 18241 13093 18275
rect 13093 18241 13127 18275
rect 13127 18241 13136 18275
rect 13084 18232 13136 18241
rect 13268 18275 13320 18284
rect 13268 18241 13277 18275
rect 13277 18241 13311 18275
rect 13311 18241 13320 18275
rect 13268 18232 13320 18241
rect 13544 18232 13596 18284
rect 14188 18275 14240 18284
rect 14188 18241 14197 18275
rect 14197 18241 14231 18275
rect 14231 18241 14240 18275
rect 14188 18232 14240 18241
rect 13820 18164 13872 18216
rect 14464 18232 14516 18284
rect 14556 18275 14608 18284
rect 14556 18241 14565 18275
rect 14565 18241 14599 18275
rect 14599 18241 14608 18275
rect 14556 18232 14608 18241
rect 15476 18232 15528 18284
rect 15752 18275 15804 18284
rect 15752 18241 15761 18275
rect 15761 18241 15795 18275
rect 15795 18241 15804 18275
rect 15752 18232 15804 18241
rect 19064 18300 19116 18352
rect 22008 18368 22060 18420
rect 16028 18207 16080 18216
rect 16028 18173 16037 18207
rect 16037 18173 16071 18207
rect 16071 18173 16080 18207
rect 16028 18164 16080 18173
rect 19892 18232 19944 18284
rect 20444 18300 20496 18352
rect 22100 18300 22152 18352
rect 22928 18300 22980 18352
rect 22836 18232 22888 18284
rect 23112 18275 23164 18284
rect 23112 18241 23121 18275
rect 23121 18241 23155 18275
rect 23155 18241 23164 18275
rect 23112 18232 23164 18241
rect 25320 18300 25372 18352
rect 17224 18207 17276 18216
rect 17224 18173 17233 18207
rect 17233 18173 17267 18207
rect 17267 18173 17276 18207
rect 17224 18164 17276 18173
rect 18696 18096 18748 18148
rect 12348 18028 12400 18080
rect 14188 18028 14240 18080
rect 16856 18028 16908 18080
rect 18236 18028 18288 18080
rect 18788 18028 18840 18080
rect 20444 18028 20496 18080
rect 21916 18164 21968 18216
rect 20996 18096 21048 18148
rect 21272 18096 21324 18148
rect 23480 18207 23532 18216
rect 23480 18173 23489 18207
rect 23489 18173 23523 18207
rect 23523 18173 23532 18207
rect 23480 18164 23532 18173
rect 24768 18232 24820 18284
rect 25044 18232 25096 18284
rect 26792 18368 26844 18420
rect 26332 18232 26384 18284
rect 24216 18164 24268 18216
rect 25596 18164 25648 18216
rect 26148 18164 26200 18216
rect 26976 18207 27028 18216
rect 26976 18173 26985 18207
rect 26985 18173 27019 18207
rect 27019 18173 27028 18207
rect 26976 18164 27028 18173
rect 28356 18164 28408 18216
rect 24492 18096 24544 18148
rect 21180 18071 21232 18080
rect 21180 18037 21189 18071
rect 21189 18037 21223 18071
rect 21223 18037 21232 18071
rect 21180 18028 21232 18037
rect 22100 18028 22152 18080
rect 27252 18028 27304 18080
rect 28264 18028 28316 18080
rect 28632 18028 28684 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 10416 17824 10468 17876
rect 10968 17824 11020 17876
rect 15476 17824 15528 17876
rect 16396 17824 16448 17876
rect 17960 17824 18012 17876
rect 15568 17756 15620 17808
rect 16488 17756 16540 17808
rect 8484 17688 8536 17740
rect 12808 17688 12860 17740
rect 15844 17688 15896 17740
rect 16396 17688 16448 17740
rect 11796 17620 11848 17672
rect 12256 17620 12308 17672
rect 13176 17663 13228 17672
rect 13176 17629 13185 17663
rect 13185 17629 13219 17663
rect 13219 17629 13228 17663
rect 13176 17620 13228 17629
rect 11980 17552 12032 17604
rect 13360 17663 13412 17672
rect 13360 17629 13369 17663
rect 13369 17629 13403 17663
rect 13403 17629 13412 17663
rect 13360 17620 13412 17629
rect 13544 17663 13596 17672
rect 13544 17629 13553 17663
rect 13553 17629 13587 17663
rect 13587 17629 13596 17663
rect 14096 17663 14148 17672
rect 13544 17620 13596 17629
rect 13820 17552 13872 17604
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 14188 17620 14240 17672
rect 16028 17620 16080 17672
rect 17868 17688 17920 17740
rect 14924 17552 14976 17604
rect 17776 17620 17828 17672
rect 17960 17663 18012 17672
rect 17960 17629 17969 17663
rect 17969 17629 18003 17663
rect 18003 17629 18012 17663
rect 18328 17731 18380 17740
rect 18328 17697 18337 17731
rect 18337 17697 18371 17731
rect 18371 17697 18380 17731
rect 20628 17824 20680 17876
rect 21824 17867 21876 17876
rect 21824 17833 21833 17867
rect 21833 17833 21867 17867
rect 21867 17833 21876 17867
rect 21824 17824 21876 17833
rect 23296 17824 23348 17876
rect 23480 17824 23532 17876
rect 26424 17867 26476 17876
rect 19432 17756 19484 17808
rect 19524 17756 19576 17808
rect 20168 17756 20220 17808
rect 18328 17688 18380 17697
rect 17960 17620 18012 17629
rect 18236 17663 18288 17672
rect 18236 17629 18248 17663
rect 18248 17629 18282 17663
rect 18282 17629 18288 17663
rect 18236 17620 18288 17629
rect 18880 17620 18932 17672
rect 19248 17663 19300 17672
rect 19248 17629 19257 17663
rect 19257 17629 19291 17663
rect 19291 17629 19300 17663
rect 19248 17620 19300 17629
rect 19984 17688 20036 17740
rect 20260 17688 20312 17740
rect 23204 17756 23256 17808
rect 23848 17756 23900 17808
rect 19708 17620 19760 17672
rect 20352 17620 20404 17672
rect 20444 17620 20496 17672
rect 24676 17731 24728 17740
rect 24676 17697 24685 17731
rect 24685 17697 24719 17731
rect 24719 17697 24728 17731
rect 24676 17688 24728 17697
rect 26424 17833 26433 17867
rect 26433 17833 26467 17867
rect 26467 17833 26476 17867
rect 26424 17824 26476 17833
rect 25596 17756 25648 17808
rect 25504 17688 25556 17740
rect 21456 17620 21508 17672
rect 22100 17620 22152 17672
rect 22284 17663 22336 17672
rect 22284 17629 22293 17663
rect 22293 17629 22327 17663
rect 22327 17629 22336 17663
rect 22284 17620 22336 17629
rect 22560 17620 22612 17672
rect 22928 17620 22980 17672
rect 23112 17620 23164 17672
rect 24860 17620 24912 17672
rect 24952 17663 25004 17672
rect 24952 17629 24961 17663
rect 24961 17629 24995 17663
rect 24995 17629 25004 17663
rect 24952 17620 25004 17629
rect 25320 17620 25372 17672
rect 25872 17663 25924 17672
rect 26148 17756 26200 17808
rect 27068 17756 27120 17808
rect 26976 17688 27028 17740
rect 25872 17629 25885 17663
rect 25885 17629 25919 17663
rect 25919 17629 25924 17663
rect 25872 17620 25924 17629
rect 26148 17620 26200 17672
rect 26516 17620 26568 17672
rect 27528 17620 27580 17672
rect 28080 17620 28132 17672
rect 28172 17552 28224 17604
rect 10784 17484 10836 17536
rect 11796 17527 11848 17536
rect 11796 17493 11805 17527
rect 11805 17493 11839 17527
rect 11839 17493 11848 17527
rect 11796 17484 11848 17493
rect 11888 17484 11940 17536
rect 15844 17484 15896 17536
rect 18604 17484 18656 17536
rect 19248 17484 19300 17536
rect 19340 17484 19392 17536
rect 20352 17484 20404 17536
rect 22744 17484 22796 17536
rect 25320 17484 25372 17536
rect 25964 17484 26016 17536
rect 27620 17484 27672 17536
rect 27712 17484 27764 17536
rect 28540 17484 28592 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 10600 17280 10652 17332
rect 13360 17280 13412 17332
rect 15660 17280 15712 17332
rect 20904 17323 20956 17332
rect 8484 17212 8536 17264
rect 13268 17212 13320 17264
rect 15108 17212 15160 17264
rect 7932 17144 7984 17196
rect 10508 17187 10560 17196
rect 10508 17153 10517 17187
rect 10517 17153 10551 17187
rect 10551 17153 10560 17187
rect 10508 17144 10560 17153
rect 12072 17187 12124 17196
rect 12072 17153 12081 17187
rect 12081 17153 12115 17187
rect 12115 17153 12124 17187
rect 12072 17144 12124 17153
rect 12256 17076 12308 17128
rect 12716 17187 12768 17196
rect 12716 17153 12725 17187
rect 12725 17153 12759 17187
rect 12759 17153 12768 17187
rect 12716 17144 12768 17153
rect 15200 17144 15252 17196
rect 17500 17187 17552 17196
rect 17500 17153 17509 17187
rect 17509 17153 17543 17187
rect 17543 17153 17552 17187
rect 17500 17144 17552 17153
rect 13360 17076 13412 17128
rect 13820 17076 13872 17128
rect 15476 17076 15528 17128
rect 16672 17076 16724 17128
rect 16948 17076 17000 17128
rect 17684 17187 17736 17196
rect 17684 17153 17693 17187
rect 17693 17153 17727 17187
rect 17727 17153 17736 17187
rect 17684 17144 17736 17153
rect 18144 17144 18196 17196
rect 18604 17144 18656 17196
rect 19616 17144 19668 17196
rect 20076 17144 20128 17196
rect 20352 17187 20404 17196
rect 20352 17153 20361 17187
rect 20361 17153 20395 17187
rect 20395 17153 20404 17187
rect 20352 17144 20404 17153
rect 18328 17076 18380 17128
rect 19984 17076 20036 17128
rect 20444 17119 20496 17128
rect 20444 17085 20453 17119
rect 20453 17085 20487 17119
rect 20487 17085 20496 17119
rect 20444 17076 20496 17085
rect 20904 17289 20913 17323
rect 20913 17289 20947 17323
rect 20947 17289 20956 17323
rect 20904 17280 20956 17289
rect 20996 17280 21048 17332
rect 22100 17280 22152 17332
rect 23388 17280 23440 17332
rect 23480 17280 23532 17332
rect 25780 17323 25832 17332
rect 21088 17212 21140 17264
rect 22192 17212 22244 17264
rect 22284 17212 22336 17264
rect 23204 17212 23256 17264
rect 25780 17289 25789 17323
rect 25789 17289 25823 17323
rect 25823 17289 25832 17323
rect 25780 17280 25832 17289
rect 26424 17280 26476 17332
rect 27160 17280 27212 17332
rect 27252 17280 27304 17332
rect 20720 17187 20772 17196
rect 20720 17153 20729 17187
rect 20729 17153 20763 17187
rect 20763 17153 20772 17187
rect 20720 17144 20772 17153
rect 21456 17144 21508 17196
rect 21824 17119 21876 17128
rect 16120 17008 16172 17060
rect 17132 17008 17184 17060
rect 9220 16983 9272 16992
rect 9220 16949 9229 16983
rect 9229 16949 9263 16983
rect 9263 16949 9272 16983
rect 9220 16940 9272 16949
rect 13084 16940 13136 16992
rect 15660 16940 15712 16992
rect 17408 16940 17460 16992
rect 17776 16940 17828 16992
rect 20352 16940 20404 16992
rect 20996 17008 21048 17060
rect 21824 17085 21833 17119
rect 21833 17085 21867 17119
rect 21867 17085 21876 17119
rect 21824 17076 21876 17085
rect 23940 17187 23992 17196
rect 23940 17153 23949 17187
rect 23949 17153 23983 17187
rect 23983 17153 23992 17187
rect 23940 17144 23992 17153
rect 23572 17008 23624 17060
rect 25964 17187 26016 17196
rect 25964 17153 25973 17187
rect 25973 17153 26007 17187
rect 26007 17153 26016 17187
rect 25964 17144 26016 17153
rect 26332 17076 26384 17128
rect 26884 17144 26936 17196
rect 26792 17076 26844 17128
rect 27252 17187 27304 17196
rect 27252 17153 27261 17187
rect 27261 17153 27295 17187
rect 27295 17153 27304 17187
rect 27528 17187 27580 17196
rect 27252 17144 27304 17153
rect 27528 17153 27537 17187
rect 27537 17153 27571 17187
rect 27571 17153 27580 17187
rect 27528 17144 27580 17153
rect 27344 17119 27396 17128
rect 27344 17085 27353 17119
rect 27353 17085 27387 17119
rect 27387 17085 27396 17119
rect 27344 17076 27396 17085
rect 27620 17076 27672 17128
rect 21088 16940 21140 16992
rect 22928 16940 22980 16992
rect 25136 16940 25188 16992
rect 25320 16983 25372 16992
rect 25320 16949 25329 16983
rect 25329 16949 25363 16983
rect 25363 16949 25372 16983
rect 25320 16940 25372 16949
rect 25412 16940 25464 16992
rect 28080 16940 28132 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 11980 16779 12032 16788
rect 11980 16745 11989 16779
rect 11989 16745 12023 16779
rect 12023 16745 12032 16779
rect 11980 16736 12032 16745
rect 15108 16779 15160 16788
rect 15108 16745 15117 16779
rect 15117 16745 15151 16779
rect 15151 16745 15160 16779
rect 15108 16736 15160 16745
rect 15660 16736 15712 16788
rect 19708 16736 19760 16788
rect 7748 16668 7800 16720
rect 8484 16600 8536 16652
rect 9220 16532 9272 16584
rect 11888 16532 11940 16584
rect 12808 16532 12860 16584
rect 13820 16532 13872 16584
rect 15752 16600 15804 16652
rect 16396 16668 16448 16720
rect 16304 16600 16356 16652
rect 14556 16532 14608 16584
rect 8208 16439 8260 16448
rect 8208 16405 8217 16439
rect 8217 16405 8251 16439
rect 8251 16405 8260 16439
rect 8208 16396 8260 16405
rect 10048 16464 10100 16516
rect 14832 16464 14884 16516
rect 15292 16464 15344 16516
rect 15660 16507 15712 16516
rect 15660 16473 15669 16507
rect 15669 16473 15703 16507
rect 15703 16473 15712 16507
rect 15660 16464 15712 16473
rect 16488 16600 16540 16652
rect 17224 16600 17276 16652
rect 16764 16532 16816 16584
rect 17408 16532 17460 16584
rect 19340 16532 19392 16584
rect 21824 16736 21876 16788
rect 22468 16532 22520 16584
rect 26792 16736 26844 16788
rect 28356 16736 28408 16788
rect 24860 16643 24912 16652
rect 24860 16609 24869 16643
rect 24869 16609 24903 16643
rect 24903 16609 24912 16643
rect 24860 16600 24912 16609
rect 25780 16600 25832 16652
rect 27068 16668 27120 16720
rect 26148 16575 26200 16584
rect 16120 16507 16172 16516
rect 16120 16473 16129 16507
rect 16129 16473 16163 16507
rect 16163 16473 16172 16507
rect 16120 16464 16172 16473
rect 16488 16464 16540 16516
rect 16672 16507 16724 16516
rect 16672 16473 16681 16507
rect 16681 16473 16715 16507
rect 16715 16473 16724 16507
rect 16672 16464 16724 16473
rect 16856 16507 16908 16516
rect 16856 16473 16865 16507
rect 16865 16473 16899 16507
rect 16899 16473 16908 16507
rect 16856 16464 16908 16473
rect 17316 16464 17368 16516
rect 19800 16464 19852 16516
rect 22192 16464 22244 16516
rect 9680 16396 9732 16448
rect 12440 16439 12492 16448
rect 12440 16405 12449 16439
rect 12449 16405 12483 16439
rect 12483 16405 12492 16439
rect 12440 16396 12492 16405
rect 14464 16396 14516 16448
rect 15108 16396 15160 16448
rect 15844 16396 15896 16448
rect 17500 16396 17552 16448
rect 17592 16396 17644 16448
rect 17960 16396 18012 16448
rect 20352 16396 20404 16448
rect 21548 16396 21600 16448
rect 22100 16396 22152 16448
rect 24584 16464 24636 16516
rect 26148 16541 26157 16575
rect 26157 16541 26191 16575
rect 26191 16541 26200 16575
rect 26148 16532 26200 16541
rect 26792 16600 26844 16652
rect 26976 16600 27028 16652
rect 26240 16464 26292 16516
rect 28724 16532 28776 16584
rect 27344 16464 27396 16516
rect 28172 16464 28224 16516
rect 22652 16396 22704 16448
rect 23020 16439 23072 16448
rect 23020 16405 23029 16439
rect 23029 16405 23063 16439
rect 23063 16405 23072 16439
rect 23020 16396 23072 16405
rect 23756 16396 23808 16448
rect 27804 16396 27856 16448
rect 27988 16396 28040 16448
rect 28632 16396 28684 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 8208 16124 8260 16176
rect 9220 16056 9272 16108
rect 9680 16099 9732 16108
rect 9680 16065 9689 16099
rect 9689 16065 9723 16099
rect 9723 16065 9732 16099
rect 9680 16056 9732 16065
rect 9772 16056 9824 16108
rect 11060 16192 11112 16244
rect 13544 16192 13596 16244
rect 12440 16124 12492 16176
rect 12624 16056 12676 16108
rect 14004 16056 14056 16108
rect 15752 16192 15804 16244
rect 17776 16192 17828 16244
rect 18512 16235 18564 16244
rect 18512 16201 18521 16235
rect 18521 16201 18555 16235
rect 18555 16201 18564 16235
rect 18512 16192 18564 16201
rect 15660 16124 15712 16176
rect 16028 16124 16080 16176
rect 20260 16192 20312 16244
rect 24676 16192 24728 16244
rect 26608 16192 26660 16244
rect 28172 16235 28224 16244
rect 15292 16099 15344 16108
rect 7840 16031 7892 16040
rect 7840 15997 7849 16031
rect 7849 15997 7883 16031
rect 7883 15997 7892 16031
rect 7840 15988 7892 15997
rect 10324 15988 10376 16040
rect 13360 16031 13412 16040
rect 13360 15997 13369 16031
rect 13369 15997 13403 16031
rect 13403 15997 13412 16031
rect 13360 15988 13412 15997
rect 8852 15920 8904 15972
rect 10876 15963 10928 15972
rect 10876 15929 10885 15963
rect 10885 15929 10919 15963
rect 10919 15929 10928 15963
rect 10876 15920 10928 15929
rect 8024 15852 8076 15904
rect 9864 15852 9916 15904
rect 11060 15852 11112 15904
rect 12256 15852 12308 15904
rect 14740 15920 14792 15972
rect 15292 16065 15301 16099
rect 15301 16065 15335 16099
rect 15335 16065 15344 16099
rect 15292 16056 15344 16065
rect 15752 16099 15804 16108
rect 15752 16065 15761 16099
rect 15761 16065 15795 16099
rect 15795 16065 15804 16099
rect 15752 16056 15804 16065
rect 16580 16056 16632 16108
rect 16764 16056 16816 16108
rect 15476 15988 15528 16040
rect 17500 16099 17552 16108
rect 17500 16065 17509 16099
rect 17509 16065 17543 16099
rect 17543 16065 17552 16099
rect 17500 16056 17552 16065
rect 19340 16124 19392 16176
rect 19248 16099 19300 16108
rect 19248 16065 19257 16099
rect 19257 16065 19291 16099
rect 19291 16065 19300 16099
rect 19248 16056 19300 16065
rect 17868 15988 17920 16040
rect 19892 16056 19944 16108
rect 20168 16056 20220 16108
rect 22652 16167 22704 16176
rect 22652 16133 22686 16167
rect 22686 16133 22704 16167
rect 22652 16124 22704 16133
rect 23388 16056 23440 16108
rect 24952 16056 25004 16108
rect 25780 16099 25832 16108
rect 25780 16065 25789 16099
rect 25789 16065 25823 16099
rect 25823 16065 25832 16099
rect 25780 16056 25832 16065
rect 26240 16056 26292 16108
rect 26884 16056 26936 16108
rect 27068 16056 27120 16108
rect 27344 16099 27396 16108
rect 27344 16065 27353 16099
rect 27353 16065 27387 16099
rect 27387 16065 27396 16099
rect 27344 16056 27396 16065
rect 28172 16201 28181 16235
rect 28181 16201 28215 16235
rect 28215 16201 28224 16235
rect 28172 16192 28224 16201
rect 28356 16099 28408 16108
rect 28356 16065 28365 16099
rect 28365 16065 28399 16099
rect 28399 16065 28408 16099
rect 28356 16056 28408 16065
rect 28632 16099 28684 16108
rect 28632 16065 28641 16099
rect 28641 16065 28675 16099
rect 28675 16065 28684 16099
rect 28632 16056 28684 16065
rect 21640 15988 21692 16040
rect 22008 15988 22060 16040
rect 16856 15920 16908 15972
rect 17684 15920 17736 15972
rect 22284 15920 22336 15972
rect 23388 15920 23440 15972
rect 24308 15920 24360 15972
rect 24584 15988 24636 16040
rect 26516 15988 26568 16040
rect 25412 15920 25464 15972
rect 26332 15920 26384 15972
rect 27344 15920 27396 15972
rect 12624 15852 12676 15904
rect 13084 15852 13136 15904
rect 16396 15852 16448 15904
rect 20168 15852 20220 15904
rect 27620 15852 27672 15904
rect 28540 15895 28592 15904
rect 28540 15861 28549 15895
rect 28549 15861 28583 15895
rect 28583 15861 28592 15895
rect 28540 15852 28592 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 9772 15648 9824 15700
rect 12624 15691 12676 15700
rect 12624 15657 12633 15691
rect 12633 15657 12667 15691
rect 12667 15657 12676 15691
rect 12624 15648 12676 15657
rect 12808 15691 12860 15700
rect 12808 15657 12817 15691
rect 12817 15657 12851 15691
rect 12851 15657 12860 15691
rect 12808 15648 12860 15657
rect 10324 15555 10376 15564
rect 10324 15521 10333 15555
rect 10333 15521 10367 15555
rect 10367 15521 10376 15555
rect 10324 15512 10376 15521
rect 15660 15648 15712 15700
rect 17500 15691 17552 15700
rect 17500 15657 17509 15691
rect 17509 15657 17543 15691
rect 17543 15657 17552 15691
rect 17684 15691 17736 15700
rect 17500 15648 17552 15657
rect 17684 15657 17693 15691
rect 17693 15657 17727 15691
rect 17727 15657 17736 15691
rect 17684 15648 17736 15657
rect 18696 15648 18748 15700
rect 20444 15648 20496 15700
rect 22652 15648 22704 15700
rect 23296 15648 23348 15700
rect 23572 15691 23624 15700
rect 23572 15657 23581 15691
rect 23581 15657 23615 15691
rect 23615 15657 23624 15691
rect 23572 15648 23624 15657
rect 16948 15580 17000 15632
rect 7840 15444 7892 15496
rect 9680 15444 9732 15496
rect 12532 15444 12584 15496
rect 13360 15444 13412 15496
rect 17316 15512 17368 15564
rect 19524 15512 19576 15564
rect 14832 15487 14884 15496
rect 14832 15453 14841 15487
rect 14841 15453 14875 15487
rect 14875 15453 14884 15487
rect 14832 15444 14884 15453
rect 15292 15444 15344 15496
rect 15476 15487 15528 15496
rect 15476 15453 15485 15487
rect 15485 15453 15519 15487
rect 15519 15453 15528 15487
rect 15476 15444 15528 15453
rect 17224 15444 17276 15496
rect 7288 15419 7340 15428
rect 7288 15385 7322 15419
rect 7322 15385 7340 15419
rect 9128 15419 9180 15428
rect 7288 15376 7340 15385
rect 9128 15385 9137 15419
rect 9137 15385 9171 15419
rect 9171 15385 9180 15419
rect 9128 15376 9180 15385
rect 10784 15376 10836 15428
rect 12440 15419 12492 15428
rect 12440 15385 12449 15419
rect 12449 15385 12483 15419
rect 12483 15385 12492 15419
rect 12440 15376 12492 15385
rect 15108 15376 15160 15428
rect 16028 15376 16080 15428
rect 9312 15351 9364 15360
rect 9312 15317 9321 15351
rect 9321 15317 9355 15351
rect 9355 15317 9364 15351
rect 9312 15308 9364 15317
rect 11704 15351 11756 15360
rect 11704 15317 11713 15351
rect 11713 15317 11747 15351
rect 11747 15317 11756 15351
rect 11704 15308 11756 15317
rect 12256 15308 12308 15360
rect 13268 15351 13320 15360
rect 13268 15317 13277 15351
rect 13277 15317 13311 15351
rect 13311 15317 13320 15351
rect 13268 15308 13320 15317
rect 14280 15308 14332 15360
rect 14740 15308 14792 15360
rect 16580 15308 16632 15360
rect 17684 15308 17736 15360
rect 19064 15444 19116 15496
rect 18696 15376 18748 15428
rect 19524 15376 19576 15428
rect 21640 15580 21692 15632
rect 22100 15580 22152 15632
rect 22284 15580 22336 15632
rect 25596 15580 25648 15632
rect 21088 15512 21140 15564
rect 21548 15512 21600 15564
rect 22468 15512 22520 15564
rect 23388 15512 23440 15564
rect 21916 15444 21968 15496
rect 22744 15487 22796 15496
rect 20168 15376 20220 15428
rect 21548 15376 21600 15428
rect 22744 15453 22753 15487
rect 22753 15453 22787 15487
rect 22787 15453 22796 15487
rect 22744 15444 22796 15453
rect 23480 15487 23532 15496
rect 23480 15453 23489 15487
rect 23489 15453 23523 15487
rect 23523 15453 23532 15487
rect 23480 15444 23532 15453
rect 22560 15376 22612 15428
rect 24860 15512 24912 15564
rect 25044 15512 25096 15564
rect 28540 15580 28592 15632
rect 27896 15555 27948 15564
rect 27896 15521 27905 15555
rect 27905 15521 27939 15555
rect 27939 15521 27948 15555
rect 27896 15512 27948 15521
rect 28448 15512 28500 15564
rect 24584 15487 24636 15496
rect 24584 15453 24615 15487
rect 24615 15453 24636 15487
rect 24584 15444 24636 15453
rect 24676 15487 24728 15496
rect 24676 15453 24685 15487
rect 24685 15453 24719 15487
rect 24719 15453 24728 15487
rect 24676 15444 24728 15453
rect 25228 15444 25280 15496
rect 27620 15487 27672 15496
rect 27620 15453 27629 15487
rect 27629 15453 27663 15487
rect 27663 15453 27672 15487
rect 27620 15444 27672 15453
rect 28080 15444 28132 15496
rect 26240 15376 26292 15428
rect 25044 15308 25096 15360
rect 27436 15351 27488 15360
rect 27436 15317 27445 15351
rect 27445 15317 27479 15351
rect 27479 15317 27488 15351
rect 27436 15308 27488 15317
rect 28356 15351 28408 15360
rect 28356 15317 28365 15351
rect 28365 15317 28399 15351
rect 28399 15317 28408 15351
rect 28356 15308 28408 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 7288 15104 7340 15156
rect 9128 15104 9180 15156
rect 10048 15147 10100 15156
rect 10048 15113 10057 15147
rect 10057 15113 10091 15147
rect 10091 15113 10100 15147
rect 10048 15104 10100 15113
rect 10784 15147 10836 15156
rect 10784 15113 10793 15147
rect 10793 15113 10827 15147
rect 10827 15113 10836 15147
rect 10784 15104 10836 15113
rect 12256 15104 12308 15156
rect 12348 15104 12400 15156
rect 17408 15104 17460 15156
rect 18420 15104 18472 15156
rect 8852 15036 8904 15088
rect 9864 15079 9916 15088
rect 9864 15045 9873 15079
rect 9873 15045 9907 15079
rect 9907 15045 9916 15079
rect 9864 15036 9916 15045
rect 11520 15079 11572 15088
rect 11520 15045 11529 15079
rect 11529 15045 11563 15079
rect 11563 15045 11572 15079
rect 11520 15036 11572 15045
rect 13084 15036 13136 15088
rect 8116 15011 8168 15020
rect 8116 14977 8150 15011
rect 8150 14977 8168 15011
rect 9680 15011 9732 15020
rect 8116 14968 8168 14977
rect 9680 14977 9689 15011
rect 9689 14977 9723 15011
rect 9723 14977 9732 15011
rect 9680 14968 9732 14977
rect 10508 14968 10560 15020
rect 15476 15036 15528 15088
rect 7840 14943 7892 14952
rect 7840 14909 7849 14943
rect 7849 14909 7883 14943
rect 7883 14909 7892 14943
rect 7840 14900 7892 14909
rect 12716 14943 12768 14952
rect 12716 14909 12725 14943
rect 12725 14909 12759 14943
rect 12759 14909 12768 14943
rect 12716 14900 12768 14909
rect 14280 14900 14332 14952
rect 14004 14832 14056 14884
rect 11704 14807 11756 14816
rect 11704 14773 11713 14807
rect 11713 14773 11747 14807
rect 11747 14773 11756 14807
rect 11704 14764 11756 14773
rect 16028 14832 16080 14884
rect 16580 14764 16632 14816
rect 17224 15011 17276 15020
rect 17224 14977 17234 15011
rect 17234 14977 17268 15011
rect 17268 14977 17276 15011
rect 17224 14968 17276 14977
rect 17224 14832 17276 14884
rect 17684 14968 17736 15020
rect 18144 14968 18196 15020
rect 18236 14968 18288 15020
rect 18604 15011 18656 15020
rect 18604 14977 18613 15011
rect 18613 14977 18647 15011
rect 18647 14977 18656 15011
rect 18604 14968 18656 14977
rect 20536 15104 20588 15156
rect 22192 15147 22244 15156
rect 22192 15113 22201 15147
rect 22201 15113 22235 15147
rect 22235 15113 22244 15147
rect 22192 15104 22244 15113
rect 26056 15104 26108 15156
rect 27896 15104 27948 15156
rect 21364 15036 21416 15088
rect 27436 15036 27488 15088
rect 17868 14832 17920 14884
rect 19248 14900 19300 14952
rect 20168 14900 20220 14952
rect 20720 14968 20772 15020
rect 22376 15011 22428 15020
rect 22376 14977 22385 15011
rect 22385 14977 22419 15011
rect 22419 14977 22428 15011
rect 22376 14968 22428 14977
rect 23020 14968 23072 15020
rect 23572 14968 23624 15020
rect 24124 15011 24176 15020
rect 24124 14977 24133 15011
rect 24133 14977 24167 15011
rect 24167 14977 24176 15011
rect 24124 14968 24176 14977
rect 24860 15011 24912 15020
rect 24860 14977 24894 15011
rect 24894 14977 24912 15011
rect 26976 15011 27028 15020
rect 24860 14968 24912 14977
rect 26976 14977 26985 15011
rect 26985 14977 27019 15011
rect 27019 14977 27028 15011
rect 26976 14968 27028 14977
rect 21824 14900 21876 14952
rect 23296 14900 23348 14952
rect 24584 14943 24636 14952
rect 24584 14909 24593 14943
rect 24593 14909 24627 14943
rect 24627 14909 24636 14943
rect 24584 14900 24636 14909
rect 18880 14832 18932 14884
rect 22100 14832 22152 14884
rect 19248 14764 19300 14816
rect 20812 14807 20864 14816
rect 20812 14773 20821 14807
rect 20821 14773 20855 14807
rect 20855 14773 20864 14807
rect 20812 14764 20864 14773
rect 23296 14807 23348 14816
rect 23296 14773 23305 14807
rect 23305 14773 23339 14807
rect 23339 14773 23348 14807
rect 23296 14764 23348 14773
rect 23940 14807 23992 14816
rect 23940 14773 23949 14807
rect 23949 14773 23983 14807
rect 23983 14773 23992 14807
rect 23940 14764 23992 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 7932 14560 7984 14612
rect 8116 14560 8168 14612
rect 9220 14560 9272 14612
rect 10692 14560 10744 14612
rect 13544 14603 13596 14612
rect 13544 14569 13553 14603
rect 13553 14569 13587 14603
rect 13587 14569 13596 14603
rect 13544 14560 13596 14569
rect 13176 14492 13228 14544
rect 17316 14560 17368 14612
rect 17408 14560 17460 14612
rect 18788 14492 18840 14544
rect 10324 14424 10376 14476
rect 14096 14467 14148 14476
rect 7748 14399 7800 14408
rect 7748 14365 7757 14399
rect 7757 14365 7791 14399
rect 7791 14365 7800 14399
rect 7748 14356 7800 14365
rect 9312 14356 9364 14408
rect 11612 14356 11664 14408
rect 12532 14399 12584 14408
rect 12532 14365 12541 14399
rect 12541 14365 12575 14399
rect 12575 14365 12584 14399
rect 12532 14356 12584 14365
rect 14096 14433 14105 14467
rect 14105 14433 14139 14467
rect 14139 14433 14148 14467
rect 14096 14424 14148 14433
rect 16212 14424 16264 14476
rect 13268 14356 13320 14408
rect 13360 14399 13412 14408
rect 13360 14365 13369 14399
rect 13369 14365 13403 14399
rect 13403 14365 13412 14399
rect 13360 14356 13412 14365
rect 14188 14356 14240 14408
rect 14372 14399 14424 14408
rect 14372 14365 14406 14399
rect 14406 14365 14424 14399
rect 14372 14356 14424 14365
rect 9220 14288 9272 14340
rect 10508 14288 10560 14340
rect 10876 14288 10928 14340
rect 13728 14288 13780 14340
rect 15108 14288 15160 14340
rect 16580 14399 16632 14408
rect 16580 14365 16589 14399
rect 16589 14365 16623 14399
rect 16623 14365 16632 14399
rect 16580 14356 16632 14365
rect 16856 14424 16908 14476
rect 22008 14560 22060 14612
rect 24860 14603 24912 14612
rect 24860 14569 24869 14603
rect 24869 14569 24903 14603
rect 24903 14569 24912 14603
rect 24860 14560 24912 14569
rect 24952 14560 25004 14612
rect 21364 14492 21416 14544
rect 15568 14288 15620 14340
rect 17132 14356 17184 14408
rect 17224 14288 17276 14340
rect 10600 14220 10652 14272
rect 11704 14220 11756 14272
rect 15476 14263 15528 14272
rect 15476 14229 15485 14263
rect 15485 14229 15519 14263
rect 15519 14229 15528 14263
rect 15476 14220 15528 14229
rect 16028 14263 16080 14272
rect 16028 14229 16037 14263
rect 16037 14229 16071 14263
rect 16071 14229 16080 14263
rect 16028 14220 16080 14229
rect 20352 14424 20404 14476
rect 22468 14467 22520 14476
rect 17776 14356 17828 14408
rect 20812 14356 20864 14408
rect 21824 14399 21876 14408
rect 21824 14365 21833 14399
rect 21833 14365 21867 14399
rect 21867 14365 21876 14399
rect 21824 14356 21876 14365
rect 22468 14433 22477 14467
rect 22477 14433 22511 14467
rect 22511 14433 22520 14467
rect 22468 14424 22520 14433
rect 25688 14424 25740 14476
rect 26056 14424 26108 14476
rect 26976 14560 27028 14612
rect 28080 14603 28132 14612
rect 28080 14569 28089 14603
rect 28089 14569 28123 14603
rect 28123 14569 28132 14603
rect 28080 14560 28132 14569
rect 28448 14560 28500 14612
rect 22652 14399 22704 14408
rect 22652 14365 22661 14399
rect 22661 14365 22695 14399
rect 22695 14365 22704 14399
rect 22652 14356 22704 14365
rect 23480 14356 23532 14408
rect 25044 14399 25096 14408
rect 25044 14365 25053 14399
rect 25053 14365 25087 14399
rect 25087 14365 25096 14399
rect 25044 14356 25096 14365
rect 28356 14356 28408 14408
rect 17868 14331 17920 14340
rect 17868 14297 17893 14331
rect 17893 14297 17920 14331
rect 17868 14288 17920 14297
rect 21732 14288 21784 14340
rect 23848 14288 23900 14340
rect 18512 14263 18564 14272
rect 18512 14229 18521 14263
rect 18521 14229 18555 14263
rect 18555 14229 18564 14263
rect 18512 14220 18564 14229
rect 20076 14220 20128 14272
rect 22468 14220 22520 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 9220 14059 9272 14068
rect 9220 14025 9229 14059
rect 9229 14025 9263 14059
rect 9263 14025 9272 14059
rect 9220 14016 9272 14025
rect 10324 14059 10376 14068
rect 10324 14025 10333 14059
rect 10333 14025 10367 14059
rect 10367 14025 10376 14059
rect 10324 14016 10376 14025
rect 14832 14016 14884 14068
rect 14924 14016 14976 14068
rect 7840 13923 7892 13932
rect 7840 13889 7849 13923
rect 7849 13889 7883 13923
rect 7883 13889 7892 13923
rect 8208 13948 8260 14000
rect 11520 13991 11572 14000
rect 11520 13957 11529 13991
rect 11529 13957 11563 13991
rect 11563 13957 11572 13991
rect 11520 13948 11572 13957
rect 12440 13948 12492 14000
rect 13268 13948 13320 14000
rect 14648 13948 14700 14000
rect 8116 13923 8168 13932
rect 7840 13880 7892 13889
rect 8116 13889 8150 13923
rect 8150 13889 8168 13923
rect 8116 13880 8168 13889
rect 10968 13880 11020 13932
rect 12624 13923 12676 13932
rect 12624 13889 12633 13923
rect 12633 13889 12667 13923
rect 12667 13889 12676 13923
rect 12624 13880 12676 13889
rect 12808 13923 12860 13932
rect 12808 13889 12817 13923
rect 12817 13889 12851 13923
rect 12851 13889 12860 13923
rect 12808 13880 12860 13889
rect 14464 13880 14516 13932
rect 16580 14016 16632 14068
rect 25320 14016 25372 14068
rect 26424 14016 26476 14068
rect 14372 13812 14424 13864
rect 15660 13880 15712 13932
rect 16120 13880 16172 13932
rect 17040 13880 17092 13932
rect 17500 13991 17552 14000
rect 17500 13957 17509 13991
rect 17509 13957 17543 13991
rect 17543 13957 17552 13991
rect 17500 13948 17552 13957
rect 18144 13948 18196 14000
rect 18052 13880 18104 13932
rect 20536 13948 20588 14000
rect 19248 13923 19300 13932
rect 19248 13889 19257 13923
rect 19257 13889 19291 13923
rect 19291 13889 19300 13923
rect 19248 13880 19300 13889
rect 20076 13880 20128 13932
rect 15476 13812 15528 13864
rect 15200 13744 15252 13796
rect 16304 13812 16356 13864
rect 17500 13812 17552 13864
rect 18420 13812 18472 13864
rect 19340 13812 19392 13864
rect 20628 13812 20680 13864
rect 21916 13880 21968 13932
rect 23296 13948 23348 14000
rect 22652 13880 22704 13932
rect 24584 13948 24636 14000
rect 27528 13948 27580 14000
rect 23940 13923 23992 13932
rect 23940 13889 23974 13923
rect 23974 13889 23992 13923
rect 23940 13880 23992 13889
rect 25596 13923 25648 13932
rect 25596 13889 25605 13923
rect 25605 13889 25639 13923
rect 25639 13889 25648 13923
rect 25596 13880 25648 13889
rect 25688 13923 25740 13932
rect 25688 13889 25698 13923
rect 25698 13889 25732 13923
rect 25732 13889 25740 13923
rect 25688 13880 25740 13889
rect 25872 13923 25924 13932
rect 25872 13889 25881 13923
rect 25881 13889 25915 13923
rect 25915 13889 25924 13923
rect 25872 13880 25924 13889
rect 26056 13923 26108 13932
rect 26056 13889 26070 13923
rect 26070 13889 26104 13923
rect 26104 13889 26108 13923
rect 26056 13880 26108 13889
rect 20904 13812 20956 13864
rect 11704 13719 11756 13728
rect 11704 13685 11713 13719
rect 11713 13685 11747 13719
rect 11747 13685 11756 13719
rect 11704 13676 11756 13685
rect 11888 13719 11940 13728
rect 11888 13685 11897 13719
rect 11897 13685 11931 13719
rect 11931 13685 11940 13719
rect 11888 13676 11940 13685
rect 13912 13676 13964 13728
rect 14280 13676 14332 13728
rect 25780 13744 25832 13796
rect 17040 13676 17092 13728
rect 17500 13676 17552 13728
rect 17868 13719 17920 13728
rect 17868 13685 17877 13719
rect 17877 13685 17911 13719
rect 17911 13685 17920 13719
rect 17868 13676 17920 13685
rect 18144 13676 18196 13728
rect 18420 13676 18472 13728
rect 19524 13676 19576 13728
rect 21088 13676 21140 13728
rect 21824 13676 21876 13728
rect 22192 13676 22244 13728
rect 24952 13676 25004 13728
rect 26240 13676 26292 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 12532 13472 12584 13524
rect 14280 13515 14332 13524
rect 11428 13404 11480 13456
rect 14280 13481 14289 13515
rect 14289 13481 14323 13515
rect 14323 13481 14332 13515
rect 14280 13472 14332 13481
rect 14648 13472 14700 13524
rect 15844 13472 15896 13524
rect 16672 13472 16724 13524
rect 17040 13515 17092 13524
rect 17040 13481 17049 13515
rect 17049 13481 17083 13515
rect 17083 13481 17092 13515
rect 17040 13472 17092 13481
rect 17592 13472 17644 13524
rect 18512 13472 18564 13524
rect 19524 13472 19576 13524
rect 20628 13472 20680 13524
rect 15108 13404 15160 13456
rect 9404 13336 9456 13388
rect 10324 13336 10376 13388
rect 12808 13336 12860 13388
rect 12164 13268 12216 13320
rect 13176 13311 13228 13320
rect 13176 13277 13185 13311
rect 13185 13277 13219 13311
rect 13219 13277 13228 13311
rect 13176 13268 13228 13277
rect 14096 13311 14148 13320
rect 14096 13277 14105 13311
rect 14105 13277 14139 13311
rect 14139 13277 14148 13311
rect 14096 13268 14148 13277
rect 16304 13336 16356 13388
rect 14464 13268 14516 13320
rect 15384 13311 15436 13320
rect 15384 13277 15393 13311
rect 15393 13277 15427 13311
rect 15427 13277 15436 13311
rect 15384 13268 15436 13277
rect 9312 13243 9364 13252
rect 9312 13209 9321 13243
rect 9321 13209 9355 13243
rect 9355 13209 9364 13243
rect 9312 13200 9364 13209
rect 9864 13200 9916 13252
rect 10784 13200 10836 13252
rect 11520 13200 11572 13252
rect 12256 13243 12308 13252
rect 12256 13209 12265 13243
rect 12265 13209 12299 13243
rect 12299 13209 12308 13243
rect 12256 13200 12308 13209
rect 12440 13243 12492 13252
rect 12440 13209 12465 13243
rect 12465 13209 12492 13243
rect 12440 13200 12492 13209
rect 13268 13200 13320 13252
rect 14556 13200 14608 13252
rect 14924 13200 14976 13252
rect 17868 13404 17920 13456
rect 22560 13472 22612 13524
rect 24584 13472 24636 13524
rect 16580 13336 16632 13388
rect 17132 13336 17184 13388
rect 8024 13132 8076 13184
rect 9680 13175 9732 13184
rect 9680 13141 9689 13175
rect 9689 13141 9723 13175
rect 9723 13141 9732 13175
rect 9680 13132 9732 13141
rect 15476 13175 15528 13184
rect 15476 13141 15485 13175
rect 15485 13141 15519 13175
rect 15519 13141 15528 13175
rect 15476 13132 15528 13141
rect 16580 13132 16632 13184
rect 16948 13132 17000 13184
rect 18052 13268 18104 13320
rect 20168 13336 20220 13388
rect 19984 13268 20036 13320
rect 21180 13404 21232 13456
rect 21640 13336 21692 13388
rect 26976 13472 27028 13524
rect 27436 13404 27488 13456
rect 28264 13404 28316 13456
rect 17960 13243 18012 13252
rect 17960 13209 17969 13243
rect 17969 13209 18003 13243
rect 18003 13209 18012 13243
rect 17960 13200 18012 13209
rect 18144 13243 18196 13252
rect 18144 13209 18169 13243
rect 18169 13209 18196 13243
rect 19248 13243 19300 13252
rect 18144 13200 18196 13209
rect 19248 13209 19257 13243
rect 19257 13209 19291 13243
rect 19291 13209 19300 13243
rect 19248 13200 19300 13209
rect 19340 13200 19392 13252
rect 20076 13200 20128 13252
rect 20168 13200 20220 13252
rect 18052 13132 18104 13184
rect 21180 13268 21232 13320
rect 21732 13268 21784 13320
rect 22192 13311 22244 13320
rect 22192 13277 22201 13311
rect 22201 13277 22235 13311
rect 22235 13277 22244 13311
rect 22192 13268 22244 13277
rect 22560 13268 22612 13320
rect 23296 13311 23348 13320
rect 23296 13277 23306 13311
rect 23306 13277 23340 13311
rect 23340 13277 23348 13311
rect 27068 13336 27120 13388
rect 23296 13268 23348 13277
rect 20996 13243 21048 13252
rect 20996 13209 21005 13243
rect 21005 13209 21039 13243
rect 21039 13209 21048 13243
rect 20996 13200 21048 13209
rect 21456 13132 21508 13184
rect 22008 13132 22060 13184
rect 24952 13200 25004 13252
rect 26240 13268 26292 13320
rect 26700 13268 26752 13320
rect 27620 13268 27672 13320
rect 25964 13200 26016 13252
rect 23664 13132 23716 13184
rect 24032 13132 24084 13184
rect 25688 13132 25740 13184
rect 27252 13132 27304 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 9864 12971 9916 12980
rect 8300 12860 8352 12912
rect 8668 12860 8720 12912
rect 9404 12860 9456 12912
rect 9864 12937 9873 12971
rect 9873 12937 9907 12971
rect 9907 12937 9916 12971
rect 9864 12928 9916 12937
rect 10508 12971 10560 12980
rect 10508 12937 10517 12971
rect 10517 12937 10551 12971
rect 10551 12937 10560 12971
rect 10508 12928 10560 12937
rect 11612 12928 11664 12980
rect 13176 12928 13228 12980
rect 13912 12928 13964 12980
rect 11060 12860 11112 12912
rect 11520 12903 11572 12912
rect 11520 12869 11529 12903
rect 11529 12869 11563 12903
rect 11563 12869 11572 12903
rect 11520 12860 11572 12869
rect 12440 12860 12492 12912
rect 12624 12860 12676 12912
rect 15752 12903 15804 12912
rect 9128 12792 9180 12844
rect 9312 12792 9364 12844
rect 10692 12835 10744 12844
rect 10692 12801 10701 12835
rect 10701 12801 10735 12835
rect 10735 12801 10744 12835
rect 10692 12792 10744 12801
rect 15752 12869 15761 12903
rect 15761 12869 15795 12903
rect 15795 12869 15804 12903
rect 15752 12860 15804 12869
rect 16948 12860 17000 12912
rect 17224 12860 17276 12912
rect 18696 12903 18748 12912
rect 18696 12869 18705 12903
rect 18705 12869 18739 12903
rect 18739 12869 18748 12903
rect 20996 12928 21048 12980
rect 23572 12928 23624 12980
rect 24124 12928 24176 12980
rect 18696 12860 18748 12869
rect 14280 12835 14332 12844
rect 14280 12801 14289 12835
rect 14289 12801 14323 12835
rect 14323 12801 14332 12835
rect 14280 12792 14332 12801
rect 15476 12792 15528 12844
rect 17684 12792 17736 12844
rect 18236 12792 18288 12844
rect 18512 12835 18564 12844
rect 18512 12801 18519 12835
rect 18519 12801 18564 12835
rect 18512 12792 18564 12801
rect 18880 12792 18932 12844
rect 21364 12860 21416 12912
rect 20444 12792 20496 12844
rect 20720 12792 20772 12844
rect 21916 12792 21968 12844
rect 23664 12860 23716 12912
rect 22652 12792 22704 12844
rect 13912 12656 13964 12708
rect 16856 12724 16908 12776
rect 17500 12724 17552 12776
rect 20904 12724 20956 12776
rect 21180 12724 21232 12776
rect 22008 12724 22060 12776
rect 23020 12724 23072 12776
rect 24032 12792 24084 12844
rect 24584 12792 24636 12844
rect 25320 12835 25372 12844
rect 25320 12801 25329 12835
rect 25329 12801 25363 12835
rect 25363 12801 25372 12835
rect 25320 12792 25372 12801
rect 27436 12928 27488 12980
rect 27528 12928 27580 12980
rect 25688 12903 25740 12912
rect 25688 12869 25697 12903
rect 25697 12869 25731 12903
rect 25731 12869 25740 12903
rect 25688 12860 25740 12869
rect 25964 12792 26016 12844
rect 26976 12835 27028 12844
rect 26976 12801 26985 12835
rect 26985 12801 27019 12835
rect 27019 12801 27028 12835
rect 26976 12792 27028 12801
rect 27712 12792 27764 12844
rect 19064 12656 19116 12708
rect 24124 12656 24176 12708
rect 25872 12724 25924 12776
rect 11704 12631 11756 12640
rect 11704 12597 11713 12631
rect 11713 12597 11747 12631
rect 11747 12597 11756 12631
rect 11704 12588 11756 12597
rect 13452 12588 13504 12640
rect 14372 12588 14424 12640
rect 15660 12588 15712 12640
rect 17040 12588 17092 12640
rect 20628 12588 20680 12640
rect 22376 12588 22428 12640
rect 25872 12588 25924 12640
rect 26792 12588 26844 12640
rect 26976 12588 27028 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 6000 12384 6052 12436
rect 8852 12384 8904 12436
rect 9128 12427 9180 12436
rect 9128 12393 9137 12427
rect 9137 12393 9171 12427
rect 9171 12393 9180 12427
rect 9128 12384 9180 12393
rect 11704 12384 11756 12436
rect 13452 12427 13504 12436
rect 13452 12393 13461 12427
rect 13461 12393 13495 12427
rect 13495 12393 13504 12427
rect 13452 12384 13504 12393
rect 10140 12316 10192 12368
rect 10232 12248 10284 12300
rect 13084 12248 13136 12300
rect 15016 12384 15068 12436
rect 15292 12384 15344 12436
rect 16488 12384 16540 12436
rect 18236 12384 18288 12436
rect 20904 12384 20956 12436
rect 21088 12384 21140 12436
rect 21548 12384 21600 12436
rect 23664 12384 23716 12436
rect 25780 12384 25832 12436
rect 26148 12384 26200 12436
rect 13728 12316 13780 12368
rect 14556 12316 14608 12368
rect 21640 12316 21692 12368
rect 13820 12248 13872 12300
rect 15660 12291 15712 12300
rect 15660 12257 15669 12291
rect 15669 12257 15703 12291
rect 15703 12257 15712 12291
rect 15660 12248 15712 12257
rect 16028 12248 16080 12300
rect 16948 12248 17000 12300
rect 17132 12291 17184 12300
rect 17132 12257 17141 12291
rect 17141 12257 17175 12291
rect 17175 12257 17184 12291
rect 17132 12248 17184 12257
rect 20352 12248 20404 12300
rect 20444 12248 20496 12300
rect 24308 12316 24360 12368
rect 28080 12316 28132 12368
rect 22100 12248 22152 12300
rect 9680 12180 9732 12232
rect 9956 12223 10008 12232
rect 9956 12189 9965 12223
rect 9965 12189 9999 12223
rect 9999 12189 10008 12223
rect 9956 12180 10008 12189
rect 10416 12223 10468 12232
rect 10416 12189 10425 12223
rect 10425 12189 10459 12223
rect 10459 12189 10468 12223
rect 10416 12180 10468 12189
rect 10692 12223 10744 12232
rect 10692 12189 10726 12223
rect 10726 12189 10744 12223
rect 10692 12180 10744 12189
rect 10968 12180 11020 12232
rect 12808 12180 12860 12232
rect 15476 12223 15528 12232
rect 15476 12189 15485 12223
rect 15485 12189 15519 12223
rect 15519 12189 15528 12223
rect 15476 12180 15528 12189
rect 15844 12223 15896 12232
rect 15844 12189 15853 12223
rect 15853 12189 15887 12223
rect 15887 12189 15896 12223
rect 15844 12180 15896 12189
rect 17500 12180 17552 12232
rect 19984 12180 20036 12232
rect 22376 12223 22428 12232
rect 10324 12112 10376 12164
rect 12440 12112 12492 12164
rect 12992 12112 13044 12164
rect 8944 12044 8996 12096
rect 9772 12087 9824 12096
rect 9772 12053 9781 12087
rect 9781 12053 9815 12087
rect 9815 12053 9824 12087
rect 9772 12044 9824 12053
rect 12532 12044 12584 12096
rect 14188 12112 14240 12164
rect 18972 12112 19024 12164
rect 20444 12112 20496 12164
rect 22376 12189 22385 12223
rect 22385 12189 22419 12223
rect 22419 12189 22428 12223
rect 22376 12180 22428 12189
rect 23664 12248 23716 12300
rect 24216 12248 24268 12300
rect 23296 12180 23348 12232
rect 23112 12112 23164 12164
rect 24216 12112 24268 12164
rect 25412 12248 25464 12300
rect 25964 12248 26016 12300
rect 13820 12044 13872 12096
rect 19340 12044 19392 12096
rect 20260 12044 20312 12096
rect 20812 12044 20864 12096
rect 21456 12044 21508 12096
rect 22652 12044 22704 12096
rect 25688 12112 25740 12164
rect 25872 12112 25924 12164
rect 26240 12223 26292 12232
rect 26240 12189 26249 12223
rect 26249 12189 26283 12223
rect 26283 12189 26292 12223
rect 26240 12180 26292 12189
rect 27436 12180 27488 12232
rect 27988 12223 28040 12232
rect 27988 12189 27997 12223
rect 27997 12189 28031 12223
rect 28031 12189 28040 12223
rect 27988 12180 28040 12189
rect 24860 12044 24912 12096
rect 27160 12044 27212 12096
rect 27528 12044 27580 12096
rect 28080 12112 28132 12164
rect 28264 12155 28316 12164
rect 28264 12121 28273 12155
rect 28273 12121 28307 12155
rect 28307 12121 28316 12155
rect 28264 12112 28316 12121
rect 28448 12044 28500 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 5908 11840 5960 11892
rect 10784 11883 10836 11892
rect 8760 11772 8812 11824
rect 10784 11849 10793 11883
rect 10793 11849 10827 11883
rect 10827 11849 10836 11883
rect 10784 11840 10836 11849
rect 10876 11840 10928 11892
rect 12532 11840 12584 11892
rect 12256 11772 12308 11824
rect 12348 11815 12400 11824
rect 12348 11781 12357 11815
rect 12357 11781 12391 11815
rect 12391 11781 12400 11815
rect 15384 11840 15436 11892
rect 15936 11840 15988 11892
rect 12348 11772 12400 11781
rect 6460 11704 6512 11756
rect 9772 11704 9824 11756
rect 11428 11704 11480 11756
rect 11888 11704 11940 11756
rect 7472 11500 7524 11552
rect 10416 11568 10468 11620
rect 12808 11704 12860 11756
rect 13728 11772 13780 11824
rect 14464 11772 14516 11824
rect 13084 11747 13136 11756
rect 13084 11713 13093 11747
rect 13093 11713 13127 11747
rect 13127 11713 13136 11747
rect 13084 11704 13136 11713
rect 14832 11704 14884 11756
rect 15660 11704 15712 11756
rect 16580 11772 16632 11824
rect 18512 11840 18564 11892
rect 19524 11772 19576 11824
rect 16856 11747 16908 11756
rect 16856 11713 16865 11747
rect 16865 11713 16899 11747
rect 16899 11713 16908 11747
rect 16856 11704 16908 11713
rect 9588 11500 9640 11552
rect 15476 11568 15528 11620
rect 15660 11568 15712 11620
rect 12900 11500 12952 11552
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 13820 11500 13872 11509
rect 14832 11500 14884 11552
rect 16672 11543 16724 11552
rect 16672 11509 16681 11543
rect 16681 11509 16715 11543
rect 16715 11509 16724 11543
rect 16672 11500 16724 11509
rect 22928 11840 22980 11892
rect 23296 11883 23348 11892
rect 23296 11849 23305 11883
rect 23305 11849 23339 11883
rect 23339 11849 23348 11883
rect 23296 11840 23348 11849
rect 23848 11840 23900 11892
rect 24860 11772 24912 11824
rect 27712 11840 27764 11892
rect 28264 11840 28316 11892
rect 26516 11772 26568 11824
rect 27252 11815 27304 11824
rect 27252 11781 27286 11815
rect 27286 11781 27304 11815
rect 27252 11772 27304 11781
rect 20352 11704 20404 11756
rect 21456 11704 21508 11756
rect 21916 11747 21968 11756
rect 21916 11713 21925 11747
rect 21925 11713 21959 11747
rect 21959 11713 21968 11747
rect 21916 11704 21968 11713
rect 23756 11704 23808 11756
rect 23112 11636 23164 11688
rect 26424 11704 26476 11756
rect 26792 11704 26844 11756
rect 23940 11679 23992 11688
rect 23940 11645 23949 11679
rect 23949 11645 23983 11679
rect 23983 11645 23992 11679
rect 24216 11679 24268 11688
rect 23940 11636 23992 11645
rect 24216 11645 24225 11679
rect 24225 11645 24259 11679
rect 24259 11645 24268 11679
rect 24216 11636 24268 11645
rect 25044 11636 25096 11688
rect 28080 11704 28132 11756
rect 29000 11747 29052 11756
rect 29000 11713 29009 11747
rect 29009 11713 29043 11747
rect 29043 11713 29052 11747
rect 29000 11704 29052 11713
rect 21732 11568 21784 11620
rect 20720 11500 20772 11552
rect 21548 11500 21600 11552
rect 22192 11500 22244 11552
rect 22284 11500 22336 11552
rect 26884 11568 26936 11620
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 9956 11296 10008 11348
rect 8300 11228 8352 11280
rect 9404 11228 9456 11280
rect 11336 11228 11388 11280
rect 12348 11296 12400 11348
rect 14188 11339 14240 11348
rect 14188 11305 14197 11339
rect 14197 11305 14231 11339
rect 14231 11305 14240 11339
rect 14188 11296 14240 11305
rect 14924 11339 14976 11348
rect 14924 11305 14933 11339
rect 14933 11305 14967 11339
rect 14967 11305 14976 11339
rect 14924 11296 14976 11305
rect 16764 11296 16816 11348
rect 17224 11296 17276 11348
rect 18052 11296 18104 11348
rect 13084 11228 13136 11280
rect 7196 11160 7248 11212
rect 6920 11135 6972 11144
rect 5448 11024 5500 11076
rect 6920 11101 6929 11135
rect 6929 11101 6963 11135
rect 6963 11101 6972 11135
rect 6920 11092 6972 11101
rect 7104 11092 7156 11144
rect 7840 11135 7892 11144
rect 7840 11101 7849 11135
rect 7849 11101 7883 11135
rect 7883 11101 7892 11135
rect 7840 11092 7892 11101
rect 8024 11160 8076 11212
rect 8116 11092 8168 11144
rect 12348 11160 12400 11212
rect 12532 11203 12584 11212
rect 12532 11169 12541 11203
rect 12541 11169 12575 11203
rect 12575 11169 12584 11203
rect 12900 11203 12952 11212
rect 12532 11160 12584 11169
rect 12900 11169 12909 11203
rect 12909 11169 12943 11203
rect 12943 11169 12952 11203
rect 12900 11160 12952 11169
rect 10968 11135 11020 11144
rect 10968 11101 10977 11135
rect 10977 11101 11011 11135
rect 11011 11101 11020 11135
rect 10968 11092 11020 11101
rect 12440 11092 12492 11144
rect 15844 11228 15896 11280
rect 19524 11228 19576 11280
rect 14464 11092 14516 11144
rect 14924 11092 14976 11144
rect 15476 11092 15528 11144
rect 16672 11160 16724 11212
rect 17132 11160 17184 11212
rect 17316 11160 17368 11212
rect 17684 11160 17736 11212
rect 15844 11135 15896 11144
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 15844 11092 15896 11101
rect 16580 11135 16632 11144
rect 7288 11024 7340 11076
rect 9680 11024 9732 11076
rect 11796 11024 11848 11076
rect 14832 11067 14884 11076
rect 14832 11033 14841 11067
rect 14841 11033 14875 11067
rect 14875 11033 14884 11067
rect 14832 11024 14884 11033
rect 16580 11101 16589 11135
rect 16589 11101 16623 11135
rect 16623 11101 16632 11135
rect 16580 11092 16632 11101
rect 16856 11135 16908 11144
rect 16856 11101 16865 11135
rect 16865 11101 16899 11135
rect 16899 11101 16908 11135
rect 16856 11092 16908 11101
rect 4620 10999 4672 11008
rect 4620 10965 4629 10999
rect 4629 10965 4663 10999
rect 4663 10965 4672 10999
rect 4620 10956 4672 10965
rect 7012 10956 7064 11008
rect 7104 10956 7156 11008
rect 9588 10956 9640 11008
rect 11060 10956 11112 11008
rect 12532 10956 12584 11008
rect 12624 10956 12676 11008
rect 17868 11024 17920 11076
rect 17132 10956 17184 11008
rect 18420 11024 18472 11076
rect 19984 11092 20036 11144
rect 20996 11296 21048 11348
rect 21640 11296 21692 11348
rect 26240 11296 26292 11348
rect 27068 11339 27120 11348
rect 27068 11305 27077 11339
rect 27077 11305 27111 11339
rect 27111 11305 27120 11339
rect 27068 11296 27120 11305
rect 21364 11228 21416 11280
rect 23112 11160 23164 11212
rect 20904 11092 20956 11144
rect 20996 11024 21048 11076
rect 21640 11092 21692 11144
rect 20904 10956 20956 11008
rect 22652 11024 22704 11076
rect 22928 11024 22980 11076
rect 23296 11228 23348 11280
rect 24216 11228 24268 11280
rect 29552 11271 29604 11280
rect 24308 11160 24360 11212
rect 29552 11237 29561 11271
rect 29561 11237 29595 11271
rect 29595 11237 29604 11271
rect 29552 11228 29604 11237
rect 23572 11135 23624 11144
rect 23572 11101 23581 11135
rect 23581 11101 23615 11135
rect 23615 11101 23624 11135
rect 23572 11092 23624 11101
rect 24216 11092 24268 11144
rect 24400 11135 24452 11144
rect 24400 11101 24409 11135
rect 24409 11101 24443 11135
rect 24443 11101 24452 11135
rect 24400 11092 24452 11101
rect 26516 11092 26568 11144
rect 27620 11135 27672 11144
rect 27620 11101 27629 11135
rect 27629 11101 27663 11135
rect 27663 11101 27672 11135
rect 27620 11092 27672 11101
rect 28448 11135 28500 11144
rect 28448 11101 28457 11135
rect 28457 11101 28491 11135
rect 28491 11101 28500 11135
rect 28448 11092 28500 11101
rect 29736 11135 29788 11144
rect 29736 11101 29745 11135
rect 29745 11101 29779 11135
rect 29779 11101 29788 11135
rect 29736 11092 29788 11101
rect 23756 11024 23808 11076
rect 24124 11024 24176 11076
rect 24308 11024 24360 11076
rect 25780 10999 25832 11008
rect 25780 10965 25789 10999
rect 25789 10965 25823 10999
rect 25823 10965 25832 10999
rect 25780 10956 25832 10965
rect 26148 11024 26200 11076
rect 27068 11024 27120 11076
rect 36268 10956 36320 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 204 10752 256 10804
rect 6460 10795 6512 10804
rect 6460 10761 6469 10795
rect 6469 10761 6503 10795
rect 6503 10761 6512 10795
rect 6460 10752 6512 10761
rect 6920 10752 6972 10804
rect 7288 10752 7340 10804
rect 7840 10752 7892 10804
rect 11796 10752 11848 10804
rect 23572 10752 23624 10804
rect 1860 10548 1912 10600
rect 5448 10591 5500 10600
rect 5448 10557 5457 10591
rect 5457 10557 5491 10591
rect 5491 10557 5500 10591
rect 5448 10548 5500 10557
rect 6368 10616 6420 10668
rect 6920 10616 6972 10668
rect 7104 10659 7156 10668
rect 7104 10625 7113 10659
rect 7113 10625 7147 10659
rect 7147 10625 7156 10659
rect 7104 10616 7156 10625
rect 7288 10659 7340 10668
rect 7288 10625 7297 10659
rect 7297 10625 7331 10659
rect 7331 10625 7340 10659
rect 7288 10616 7340 10625
rect 7564 10616 7616 10668
rect 8392 10659 8444 10668
rect 8392 10625 8401 10659
rect 8401 10625 8435 10659
rect 8435 10625 8444 10659
rect 8392 10616 8444 10625
rect 8944 10616 8996 10668
rect 11796 10616 11848 10668
rect 12072 10659 12124 10668
rect 12072 10625 12081 10659
rect 12081 10625 12115 10659
rect 12115 10625 12124 10659
rect 12072 10616 12124 10625
rect 12900 10616 12952 10668
rect 4712 10455 4764 10464
rect 4712 10421 4721 10455
rect 4721 10421 4755 10455
rect 4755 10421 4764 10455
rect 4712 10412 4764 10421
rect 8208 10455 8260 10464
rect 8208 10421 8217 10455
rect 8217 10421 8251 10455
rect 8251 10421 8260 10455
rect 8208 10412 8260 10421
rect 12716 10548 12768 10600
rect 10416 10480 10468 10532
rect 10968 10523 11020 10532
rect 10968 10489 10977 10523
rect 10977 10489 11011 10523
rect 11011 10489 11020 10523
rect 10968 10480 11020 10489
rect 11336 10480 11388 10532
rect 15660 10659 15712 10668
rect 15660 10625 15669 10659
rect 15669 10625 15703 10659
rect 15703 10625 15712 10659
rect 15660 10616 15712 10625
rect 15844 10659 15896 10668
rect 15844 10625 15853 10659
rect 15853 10625 15887 10659
rect 15887 10625 15896 10659
rect 15844 10616 15896 10625
rect 17132 10659 17184 10668
rect 17132 10625 17141 10659
rect 17141 10625 17175 10659
rect 17175 10625 17184 10659
rect 17132 10616 17184 10625
rect 19432 10684 19484 10736
rect 18512 10659 18564 10668
rect 18512 10625 18521 10659
rect 18521 10625 18555 10659
rect 18555 10625 18564 10659
rect 18512 10616 18564 10625
rect 20720 10684 20772 10736
rect 19892 10659 19944 10668
rect 19892 10625 19926 10659
rect 19926 10625 19944 10659
rect 19892 10616 19944 10625
rect 23296 10684 23348 10736
rect 24216 10727 24268 10736
rect 24216 10693 24225 10727
rect 24225 10693 24259 10727
rect 24259 10693 24268 10727
rect 24216 10684 24268 10693
rect 22284 10659 22336 10668
rect 22284 10625 22318 10659
rect 22318 10625 22336 10659
rect 22284 10616 22336 10625
rect 24860 10659 24912 10668
rect 24860 10625 24869 10659
rect 24869 10625 24903 10659
rect 24903 10625 24912 10659
rect 24860 10616 24912 10625
rect 26516 10684 26568 10736
rect 9956 10412 10008 10464
rect 12440 10412 12492 10464
rect 12716 10412 12768 10464
rect 17868 10548 17920 10600
rect 24492 10548 24544 10600
rect 25044 10548 25096 10600
rect 14832 10480 14884 10532
rect 18144 10480 18196 10532
rect 19616 10480 19668 10532
rect 20996 10523 21048 10532
rect 20996 10489 21005 10523
rect 21005 10489 21039 10523
rect 21039 10489 21048 10523
rect 20996 10480 21048 10489
rect 25320 10616 25372 10668
rect 27436 10659 27488 10668
rect 27436 10625 27445 10659
rect 27445 10625 27479 10659
rect 27479 10625 27488 10659
rect 27436 10616 27488 10625
rect 27712 10616 27764 10668
rect 28448 10616 28500 10668
rect 29000 10684 29052 10736
rect 28632 10548 28684 10600
rect 30196 10659 30248 10668
rect 30196 10625 30205 10659
rect 30205 10625 30239 10659
rect 30239 10625 30248 10659
rect 30196 10616 30248 10625
rect 30288 10616 30340 10668
rect 25780 10480 25832 10532
rect 28724 10523 28776 10532
rect 28724 10489 28733 10523
rect 28733 10489 28767 10523
rect 28767 10489 28776 10523
rect 28724 10480 28776 10489
rect 28816 10480 28868 10532
rect 17868 10412 17920 10464
rect 18604 10412 18656 10464
rect 24308 10412 24360 10464
rect 25412 10455 25464 10464
rect 25412 10421 25421 10455
rect 25421 10421 25455 10455
rect 25455 10421 25464 10455
rect 25412 10412 25464 10421
rect 25872 10412 25924 10464
rect 26240 10412 26292 10464
rect 27620 10412 27672 10464
rect 29368 10455 29420 10464
rect 29368 10421 29377 10455
rect 29377 10421 29411 10455
rect 29411 10421 29420 10455
rect 29368 10412 29420 10421
rect 30656 10455 30708 10464
rect 30656 10421 30665 10455
rect 30665 10421 30699 10455
rect 30699 10421 30708 10455
rect 30656 10412 30708 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 6368 10251 6420 10260
rect 6368 10217 6377 10251
rect 6377 10217 6411 10251
rect 6411 10217 6420 10251
rect 6368 10208 6420 10217
rect 7012 10208 7064 10260
rect 8116 10251 8168 10260
rect 8116 10217 8125 10251
rect 8125 10217 8159 10251
rect 8159 10217 8168 10251
rect 8116 10208 8168 10217
rect 8392 10208 8444 10260
rect 3976 10047 4028 10056
rect 3976 10013 3985 10047
rect 3985 10013 4019 10047
rect 4019 10013 4028 10047
rect 3976 10004 4028 10013
rect 4712 10004 4764 10056
rect 2964 9936 3016 9988
rect 5540 10004 5592 10056
rect 7288 10140 7340 10192
rect 12164 10140 12216 10192
rect 17040 10208 17092 10260
rect 18512 10208 18564 10260
rect 21088 10208 21140 10260
rect 7104 10047 7156 10056
rect 7104 10013 7113 10047
rect 7113 10013 7147 10047
rect 7147 10013 7156 10047
rect 7104 10004 7156 10013
rect 7288 10047 7340 10056
rect 7288 10013 7297 10047
rect 7297 10013 7331 10047
rect 7331 10013 7340 10047
rect 7288 10004 7340 10013
rect 8208 10072 8260 10124
rect 7564 10004 7616 10056
rect 8852 10004 8904 10056
rect 6920 9936 6972 9988
rect 12440 10115 12492 10124
rect 12440 10081 12449 10115
rect 12449 10081 12483 10115
rect 12483 10081 12492 10115
rect 12440 10072 12492 10081
rect 13636 10072 13688 10124
rect 12624 10047 12676 10056
rect 12624 10013 12633 10047
rect 12633 10013 12667 10047
rect 12667 10013 12676 10047
rect 12624 10004 12676 10013
rect 15200 10072 15252 10124
rect 17132 10072 17184 10124
rect 23296 10208 23348 10260
rect 23480 10251 23532 10260
rect 23480 10217 23489 10251
rect 23489 10217 23523 10251
rect 23523 10217 23532 10251
rect 23480 10208 23532 10217
rect 22652 10140 22704 10192
rect 14464 10047 14516 10056
rect 10968 9936 11020 9988
rect 14464 10013 14473 10047
rect 14473 10013 14507 10047
rect 14507 10013 14516 10047
rect 14464 10004 14516 10013
rect 14832 10047 14884 10056
rect 14832 10013 14841 10047
rect 14841 10013 14875 10047
rect 14875 10013 14884 10047
rect 14832 10004 14884 10013
rect 17776 10004 17828 10056
rect 20352 10072 20404 10124
rect 23756 10072 23808 10124
rect 19432 10047 19484 10056
rect 19432 10013 19441 10047
rect 19441 10013 19475 10047
rect 19475 10013 19484 10047
rect 19432 10004 19484 10013
rect 22376 10004 22428 10056
rect 26700 10208 26752 10260
rect 26976 10208 27028 10260
rect 27252 10208 27304 10260
rect 27988 10208 28040 10260
rect 28908 10208 28960 10260
rect 29184 10140 29236 10192
rect 26884 10072 26936 10124
rect 28724 10072 28776 10124
rect 24952 10047 25004 10056
rect 13544 9979 13596 9988
rect 13544 9945 13553 9979
rect 13553 9945 13587 9979
rect 13587 9945 13596 9979
rect 14648 9979 14700 9988
rect 13544 9936 13596 9945
rect 14648 9945 14657 9979
rect 14657 9945 14691 9979
rect 14691 9945 14700 9979
rect 14648 9936 14700 9945
rect 11244 9868 11296 9920
rect 12348 9868 12400 9920
rect 13728 9868 13780 9920
rect 14096 9868 14148 9920
rect 16396 9936 16448 9988
rect 18604 9936 18656 9988
rect 19984 9936 20036 9988
rect 20444 9936 20496 9988
rect 21548 9936 21600 9988
rect 24952 10013 24961 10047
rect 24961 10013 24995 10047
rect 24995 10013 25004 10047
rect 24952 10004 25004 10013
rect 25412 10004 25464 10056
rect 23848 9936 23900 9988
rect 25044 9936 25096 9988
rect 29368 10004 29420 10056
rect 29736 10047 29788 10056
rect 29736 10013 29745 10047
rect 29745 10013 29779 10047
rect 29779 10013 29788 10047
rect 29736 10004 29788 10013
rect 26884 9936 26936 9988
rect 27436 9936 27488 9988
rect 19340 9911 19392 9920
rect 19340 9877 19349 9911
rect 19349 9877 19383 9911
rect 19383 9877 19392 9911
rect 19340 9868 19392 9877
rect 20904 9868 20956 9920
rect 21180 9911 21232 9920
rect 21180 9877 21189 9911
rect 21189 9877 21223 9911
rect 21223 9877 21232 9911
rect 21180 9868 21232 9877
rect 23572 9868 23624 9920
rect 26976 9868 27028 9920
rect 29000 9911 29052 9920
rect 29000 9877 29009 9911
rect 29009 9877 29043 9911
rect 29043 9877 29052 9911
rect 29000 9868 29052 9877
rect 30104 9868 30156 9920
rect 31024 9911 31076 9920
rect 31024 9877 31033 9911
rect 31033 9877 31067 9911
rect 31067 9877 31076 9911
rect 31024 9868 31076 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 7104 9664 7156 9716
rect 7380 9664 7432 9716
rect 9128 9664 9180 9716
rect 12072 9664 12124 9716
rect 3976 9596 4028 9648
rect 9680 9596 9732 9648
rect 10232 9596 10284 9648
rect 11796 9639 11848 9648
rect 11796 9605 11805 9639
rect 11805 9605 11839 9639
rect 11839 9605 11848 9639
rect 11796 9596 11848 9605
rect 4620 9528 4672 9580
rect 6368 9571 6420 9580
rect 6368 9537 6377 9571
rect 6377 9537 6411 9571
rect 6411 9537 6420 9571
rect 6368 9528 6420 9537
rect 8116 9528 8168 9580
rect 5264 9367 5316 9376
rect 5264 9333 5273 9367
rect 5273 9333 5307 9367
rect 5307 9333 5316 9367
rect 5264 9324 5316 9333
rect 5632 9324 5684 9376
rect 9496 9528 9548 9580
rect 10600 9571 10652 9580
rect 8760 9503 8812 9512
rect 8760 9469 8769 9503
rect 8769 9469 8803 9503
rect 8803 9469 8812 9503
rect 8760 9460 8812 9469
rect 10600 9537 10609 9571
rect 10609 9537 10643 9571
rect 10643 9537 10652 9571
rect 10600 9528 10652 9537
rect 10784 9571 10836 9580
rect 10784 9537 10793 9571
rect 10793 9537 10827 9571
rect 10827 9537 10836 9571
rect 10784 9528 10836 9537
rect 9864 9460 9916 9512
rect 11244 9528 11296 9580
rect 24308 9664 24360 9716
rect 25320 9664 25372 9716
rect 25412 9664 25464 9716
rect 26884 9664 26936 9716
rect 27160 9664 27212 9716
rect 32496 9664 32548 9716
rect 13728 9596 13780 9648
rect 14832 9596 14884 9648
rect 17684 9596 17736 9648
rect 19340 9596 19392 9648
rect 19432 9596 19484 9648
rect 20168 9596 20220 9648
rect 11152 9460 11204 9512
rect 12716 9571 12768 9580
rect 12716 9537 12725 9571
rect 12725 9537 12759 9571
rect 12759 9537 12768 9571
rect 12716 9528 12768 9537
rect 14096 9571 14148 9580
rect 14096 9537 14105 9571
rect 14105 9537 14139 9571
rect 14139 9537 14148 9571
rect 14096 9528 14148 9537
rect 15292 9571 15344 9580
rect 15292 9537 15301 9571
rect 15301 9537 15335 9571
rect 15335 9537 15344 9571
rect 15292 9528 15344 9537
rect 16396 9528 16448 9580
rect 17960 9528 18012 9580
rect 18236 9528 18288 9580
rect 18604 9528 18656 9580
rect 18788 9528 18840 9580
rect 19800 9528 19852 9580
rect 20536 9596 20588 9648
rect 20720 9596 20772 9648
rect 20352 9571 20404 9580
rect 20352 9537 20361 9571
rect 20361 9537 20395 9571
rect 20395 9537 20404 9571
rect 20352 9528 20404 9537
rect 21180 9528 21232 9580
rect 21272 9571 21324 9580
rect 21272 9537 21281 9571
rect 21281 9537 21315 9571
rect 21315 9537 21324 9571
rect 22468 9571 22520 9580
rect 21272 9528 21324 9537
rect 22468 9537 22477 9571
rect 22477 9537 22511 9571
rect 22511 9537 22520 9571
rect 22468 9528 22520 9537
rect 23480 9596 23532 9648
rect 24400 9596 24452 9648
rect 24860 9596 24912 9648
rect 22836 9571 22888 9580
rect 22836 9537 22845 9571
rect 22845 9537 22879 9571
rect 22879 9537 22888 9571
rect 22836 9528 22888 9537
rect 24492 9528 24544 9580
rect 24768 9528 24820 9580
rect 25320 9571 25372 9580
rect 25320 9537 25329 9571
rect 25329 9537 25363 9571
rect 25363 9537 25372 9571
rect 25320 9528 25372 9537
rect 26056 9528 26108 9580
rect 26976 9528 27028 9580
rect 13728 9460 13780 9512
rect 11796 9392 11848 9444
rect 12624 9392 12676 9444
rect 10232 9324 10284 9376
rect 11244 9324 11296 9376
rect 16672 9503 16724 9512
rect 16672 9469 16681 9503
rect 16681 9469 16715 9503
rect 16715 9469 16724 9503
rect 16672 9460 16724 9469
rect 16948 9392 17000 9444
rect 17960 9392 18012 9444
rect 18696 9392 18748 9444
rect 15660 9324 15712 9376
rect 17592 9324 17644 9376
rect 18972 9367 19024 9376
rect 18972 9333 18981 9367
rect 18981 9333 19015 9367
rect 19015 9333 19024 9367
rect 18972 9324 19024 9333
rect 19248 9367 19300 9376
rect 19248 9333 19257 9367
rect 19257 9333 19291 9367
rect 19291 9333 19300 9367
rect 19248 9324 19300 9333
rect 20076 9367 20128 9376
rect 20076 9333 20085 9367
rect 20085 9333 20119 9367
rect 20119 9333 20128 9367
rect 20076 9324 20128 9333
rect 20720 9392 20772 9444
rect 22100 9460 22152 9512
rect 22192 9392 22244 9444
rect 22928 9392 22980 9444
rect 24676 9460 24728 9512
rect 26700 9460 26752 9512
rect 27988 9596 28040 9648
rect 27896 9571 27948 9580
rect 27896 9537 27905 9571
rect 27905 9537 27939 9571
rect 27939 9537 27948 9571
rect 27896 9528 27948 9537
rect 28080 9571 28132 9580
rect 28080 9537 28089 9571
rect 28089 9537 28123 9571
rect 28123 9537 28132 9571
rect 28080 9528 28132 9537
rect 29000 9596 29052 9648
rect 28632 9571 28684 9580
rect 28632 9537 28641 9571
rect 28641 9537 28675 9571
rect 28675 9537 28684 9571
rect 28632 9528 28684 9537
rect 29276 9571 29328 9580
rect 29276 9537 29285 9571
rect 29285 9537 29319 9571
rect 29319 9537 29328 9571
rect 29276 9528 29328 9537
rect 29368 9528 29420 9580
rect 30932 9528 30984 9580
rect 31208 9571 31260 9580
rect 31208 9537 31217 9571
rect 31217 9537 31251 9571
rect 31251 9537 31260 9571
rect 31208 9528 31260 9537
rect 24952 9392 25004 9444
rect 25136 9392 25188 9444
rect 25596 9392 25648 9444
rect 21364 9324 21416 9376
rect 22744 9367 22796 9376
rect 22744 9333 22753 9367
rect 22753 9333 22787 9367
rect 22787 9333 22796 9367
rect 22744 9324 22796 9333
rect 23940 9324 23992 9376
rect 25504 9324 25556 9376
rect 25964 9367 26016 9376
rect 25964 9333 25973 9367
rect 25973 9333 26007 9367
rect 26007 9333 26016 9367
rect 25964 9324 26016 9333
rect 26056 9324 26108 9376
rect 30748 9324 30800 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 7196 9120 7248 9172
rect 8024 9163 8076 9172
rect 8024 9129 8033 9163
rect 8033 9129 8067 9163
rect 8067 9129 8076 9163
rect 8024 9120 8076 9129
rect 13728 9120 13780 9172
rect 18696 9163 18748 9172
rect 16212 9052 16264 9104
rect 6276 8984 6328 9036
rect 2136 8848 2188 8900
rect 5264 8916 5316 8968
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 5540 8959 5592 8968
rect 5356 8916 5408 8925
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 5816 8959 5868 8968
rect 5816 8925 5825 8959
rect 5825 8925 5859 8959
rect 5859 8925 5868 8959
rect 5816 8916 5868 8925
rect 5908 8959 5960 8968
rect 5908 8925 5917 8959
rect 5917 8925 5951 8959
rect 5951 8925 5960 8959
rect 7564 8984 7616 9036
rect 5908 8916 5960 8925
rect 3148 8780 3200 8832
rect 4988 8780 5040 8832
rect 7472 8959 7524 8968
rect 7472 8925 7481 8959
rect 7481 8925 7515 8959
rect 7515 8925 7524 8959
rect 7472 8916 7524 8925
rect 8576 8916 8628 8968
rect 10048 8916 10100 8968
rect 10968 8916 11020 8968
rect 14280 8984 14332 9036
rect 7288 8848 7340 8900
rect 9036 8848 9088 8900
rect 9404 8848 9456 8900
rect 10140 8848 10192 8900
rect 13728 8916 13780 8968
rect 15108 8959 15160 8968
rect 15108 8925 15117 8959
rect 15117 8925 15151 8959
rect 15151 8925 15160 8959
rect 15108 8916 15160 8925
rect 15292 8916 15344 8968
rect 17316 9052 17368 9104
rect 18696 9129 18705 9163
rect 18705 9129 18739 9163
rect 18739 9129 18748 9163
rect 18696 9120 18748 9129
rect 21180 9163 21232 9172
rect 21180 9129 21189 9163
rect 21189 9129 21223 9163
rect 21223 9129 21232 9163
rect 21180 9120 21232 9129
rect 21364 9120 21416 9172
rect 22284 9120 22336 9172
rect 22744 9120 22796 9172
rect 22836 9120 22888 9172
rect 23756 9120 23808 9172
rect 32772 9120 32824 9172
rect 21916 9052 21968 9104
rect 25504 9052 25556 9104
rect 26240 9052 26292 9104
rect 16672 9027 16724 9036
rect 16672 8993 16681 9027
rect 16681 8993 16715 9027
rect 16715 8993 16724 9027
rect 16672 8984 16724 8993
rect 24400 9027 24452 9036
rect 24400 8993 24409 9027
rect 24409 8993 24443 9027
rect 24443 8993 24452 9027
rect 24400 8984 24452 8993
rect 16580 8916 16632 8968
rect 17132 8916 17184 8968
rect 17868 8916 17920 8968
rect 20628 8916 20680 8968
rect 25964 8916 26016 8968
rect 7840 8780 7892 8832
rect 8484 8780 8536 8832
rect 12532 8848 12584 8900
rect 11336 8780 11388 8832
rect 11796 8780 11848 8832
rect 13360 8780 13412 8832
rect 16396 8848 16448 8900
rect 16672 8848 16724 8900
rect 17592 8891 17644 8900
rect 17592 8857 17626 8891
rect 17626 8857 17644 8891
rect 17592 8848 17644 8857
rect 17684 8848 17736 8900
rect 14924 8823 14976 8832
rect 14924 8789 14933 8823
rect 14933 8789 14967 8823
rect 14967 8789 14976 8823
rect 14924 8780 14976 8789
rect 17960 8780 18012 8832
rect 21824 8848 21876 8900
rect 29184 8984 29236 9036
rect 26332 8916 26384 8968
rect 26608 8959 26660 8968
rect 26608 8925 26617 8959
rect 26617 8925 26651 8959
rect 26651 8925 26660 8959
rect 26608 8916 26660 8925
rect 26700 8916 26752 8968
rect 27344 8916 27396 8968
rect 27804 8959 27856 8968
rect 27804 8925 27813 8959
rect 27813 8925 27847 8959
rect 27847 8925 27856 8959
rect 27804 8916 27856 8925
rect 28080 8959 28132 8968
rect 28080 8925 28089 8959
rect 28089 8925 28123 8959
rect 28123 8925 28132 8959
rect 28080 8916 28132 8925
rect 28356 8959 28408 8968
rect 28356 8925 28365 8959
rect 28365 8925 28399 8959
rect 28399 8925 28408 8959
rect 28356 8916 28408 8925
rect 28632 8959 28684 8968
rect 28632 8925 28641 8959
rect 28641 8925 28675 8959
rect 28675 8925 28684 8959
rect 28632 8916 28684 8925
rect 30196 8916 30248 8968
rect 30656 8916 30708 8968
rect 31208 8959 31260 8968
rect 31208 8925 31217 8959
rect 31217 8925 31251 8959
rect 31251 8925 31260 8959
rect 31208 8916 31260 8925
rect 31852 8959 31904 8968
rect 31852 8925 31861 8959
rect 31861 8925 31895 8959
rect 31895 8925 31904 8959
rect 31852 8916 31904 8925
rect 24308 8780 24360 8832
rect 24860 8780 24912 8832
rect 26608 8780 26660 8832
rect 26884 8780 26936 8832
rect 27436 8780 27488 8832
rect 28172 8891 28224 8900
rect 28172 8857 28181 8891
rect 28181 8857 28215 8891
rect 28215 8857 28224 8891
rect 28172 8848 28224 8857
rect 29920 8848 29972 8900
rect 29736 8780 29788 8832
rect 30564 8780 30616 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 5172 8576 5224 8628
rect 5632 8619 5684 8628
rect 5632 8585 5641 8619
rect 5641 8585 5675 8619
rect 5675 8585 5684 8619
rect 5632 8576 5684 8585
rect 5724 8508 5776 8560
rect 1308 8440 1360 8492
rect 3976 8440 4028 8492
rect 4896 8440 4948 8492
rect 5632 8440 5684 8492
rect 10324 8619 10376 8628
rect 10324 8585 10333 8619
rect 10333 8585 10367 8619
rect 10367 8585 10376 8619
rect 10324 8576 10376 8585
rect 7012 8440 7064 8492
rect 5080 8415 5132 8424
rect 1952 8236 2004 8288
rect 5080 8381 5089 8415
rect 5089 8381 5123 8415
rect 5123 8381 5132 8415
rect 5080 8372 5132 8381
rect 5264 8372 5316 8424
rect 8484 8508 8536 8560
rect 9864 8508 9916 8560
rect 10876 8508 10928 8560
rect 13912 8619 13964 8628
rect 13912 8585 13921 8619
rect 13921 8585 13955 8619
rect 13955 8585 13964 8619
rect 13912 8576 13964 8585
rect 16580 8576 16632 8628
rect 16672 8576 16724 8628
rect 18604 8576 18656 8628
rect 24492 8619 24544 8628
rect 11704 8551 11756 8560
rect 11704 8517 11713 8551
rect 11713 8517 11747 8551
rect 11747 8517 11756 8551
rect 11704 8508 11756 8517
rect 7380 8483 7432 8492
rect 7380 8449 7389 8483
rect 7389 8449 7423 8483
rect 7423 8449 7432 8483
rect 7380 8440 7432 8449
rect 8300 8483 8352 8492
rect 8300 8449 8309 8483
rect 8309 8449 8343 8483
rect 8343 8449 8352 8483
rect 8300 8440 8352 8449
rect 8392 8440 8444 8492
rect 9312 8483 9364 8492
rect 9312 8449 9321 8483
rect 9321 8449 9355 8483
rect 9355 8449 9364 8483
rect 9312 8440 9364 8449
rect 9496 8440 9548 8492
rect 10140 8483 10192 8492
rect 10140 8449 10149 8483
rect 10149 8449 10183 8483
rect 10183 8449 10192 8483
rect 10140 8440 10192 8449
rect 9772 8372 9824 8424
rect 11244 8440 11296 8492
rect 11520 8483 11572 8492
rect 11520 8449 11529 8483
rect 11529 8449 11563 8483
rect 11563 8449 11572 8483
rect 11520 8440 11572 8449
rect 12716 8483 12768 8492
rect 12716 8449 12725 8483
rect 12725 8449 12759 8483
rect 12759 8449 12768 8483
rect 12716 8440 12768 8449
rect 14464 8508 14516 8560
rect 14924 8508 14976 8560
rect 13544 8483 13596 8492
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 13728 8483 13780 8492
rect 13728 8449 13737 8483
rect 13737 8449 13771 8483
rect 13771 8449 13780 8483
rect 13728 8440 13780 8449
rect 16580 8440 16632 8492
rect 14648 8372 14700 8424
rect 19432 8508 19484 8560
rect 20260 8551 20312 8560
rect 20260 8517 20269 8551
rect 20269 8517 20303 8551
rect 20303 8517 20312 8551
rect 20260 8508 20312 8517
rect 24492 8585 24501 8619
rect 24501 8585 24535 8619
rect 24535 8585 24544 8619
rect 24492 8576 24544 8585
rect 26056 8576 26108 8628
rect 26332 8619 26384 8628
rect 26332 8585 26341 8619
rect 26341 8585 26375 8619
rect 26375 8585 26384 8619
rect 26332 8576 26384 8585
rect 17132 8483 17184 8492
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 17224 8483 17276 8492
rect 17224 8449 17233 8483
rect 17233 8449 17267 8483
rect 17267 8449 17276 8483
rect 17868 8483 17920 8492
rect 17224 8440 17276 8449
rect 17868 8449 17877 8483
rect 17877 8449 17911 8483
rect 17911 8449 17920 8483
rect 17868 8440 17920 8449
rect 18144 8483 18196 8492
rect 18144 8449 18178 8483
rect 18178 8449 18196 8483
rect 18144 8440 18196 8449
rect 20076 8483 20128 8492
rect 20076 8449 20085 8483
rect 20085 8449 20119 8483
rect 20119 8449 20128 8483
rect 20076 8440 20128 8449
rect 17776 8372 17828 8424
rect 18972 8372 19024 8424
rect 22100 8483 22152 8492
rect 22100 8449 22134 8483
rect 22134 8449 22152 8483
rect 22100 8440 22152 8449
rect 23940 8483 23992 8492
rect 23940 8449 23949 8483
rect 23949 8449 23983 8483
rect 23983 8449 23992 8483
rect 23940 8440 23992 8449
rect 20628 8372 20680 8424
rect 25964 8508 26016 8560
rect 24308 8483 24360 8492
rect 24308 8449 24317 8483
rect 24317 8449 24351 8483
rect 24351 8449 24360 8483
rect 24308 8440 24360 8449
rect 25044 8440 25096 8492
rect 25596 8440 25648 8492
rect 25780 8440 25832 8492
rect 28172 8576 28224 8628
rect 28356 8576 28408 8628
rect 29184 8619 29236 8628
rect 29184 8585 29193 8619
rect 29193 8585 29227 8619
rect 29227 8585 29236 8619
rect 29184 8576 29236 8585
rect 29736 8576 29788 8628
rect 32680 8576 32732 8628
rect 24860 8372 24912 8424
rect 25964 8372 26016 8424
rect 27436 8440 27488 8492
rect 29828 8483 29880 8492
rect 29828 8449 29837 8483
rect 29837 8449 29871 8483
rect 29871 8449 29880 8483
rect 29828 8440 29880 8449
rect 28356 8372 28408 8424
rect 30840 8440 30892 8492
rect 33140 8483 33192 8492
rect 7564 8347 7616 8356
rect 7564 8313 7573 8347
rect 7573 8313 7607 8347
rect 7607 8313 7616 8347
rect 7564 8304 7616 8313
rect 8116 8347 8168 8356
rect 8116 8313 8125 8347
rect 8125 8313 8159 8347
rect 8159 8313 8168 8347
rect 8116 8304 8168 8313
rect 9312 8304 9364 8356
rect 10140 8304 10192 8356
rect 10692 8304 10744 8356
rect 6460 8279 6512 8288
rect 6460 8245 6469 8279
rect 6469 8245 6503 8279
rect 6503 8245 6512 8279
rect 6460 8236 6512 8245
rect 6644 8236 6696 8288
rect 7656 8236 7708 8288
rect 14924 8304 14976 8356
rect 15200 8304 15252 8356
rect 16396 8304 16448 8356
rect 18880 8304 18932 8356
rect 13084 8279 13136 8288
rect 13084 8245 13093 8279
rect 13093 8245 13127 8279
rect 13127 8245 13136 8279
rect 13084 8236 13136 8245
rect 13452 8236 13504 8288
rect 16028 8236 16080 8288
rect 16120 8236 16172 8288
rect 21456 8236 21508 8288
rect 22192 8236 22244 8288
rect 28264 8236 28316 8288
rect 30012 8304 30064 8356
rect 32404 8304 32456 8356
rect 33140 8449 33149 8483
rect 33149 8449 33183 8483
rect 33183 8449 33192 8483
rect 33140 8440 33192 8449
rect 34704 8440 34756 8492
rect 32956 8372 33008 8424
rect 33600 8304 33652 8356
rect 35440 8236 35492 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 2044 8032 2096 8084
rect 4620 7964 4672 8016
rect 9496 8032 9548 8084
rect 9772 8032 9824 8084
rect 9864 8032 9916 8084
rect 10416 8075 10468 8084
rect 10416 8041 10425 8075
rect 10425 8041 10459 8075
rect 10459 8041 10468 8075
rect 10416 8032 10468 8041
rect 10600 8032 10652 8084
rect 12440 8032 12492 8084
rect 13544 8032 13596 8084
rect 16120 8075 16172 8084
rect 16120 8041 16129 8075
rect 16129 8041 16163 8075
rect 16163 8041 16172 8075
rect 16120 8032 16172 8041
rect 16580 8075 16632 8084
rect 16580 8041 16589 8075
rect 16589 8041 16623 8075
rect 16623 8041 16632 8075
rect 16580 8032 16632 8041
rect 17500 8075 17552 8084
rect 17500 8041 17509 8075
rect 17509 8041 17543 8075
rect 17543 8041 17552 8075
rect 17500 8032 17552 8041
rect 18144 8032 18196 8084
rect 21272 8032 21324 8084
rect 22100 8032 22152 8084
rect 22284 8075 22336 8084
rect 22284 8041 22293 8075
rect 22293 8041 22327 8075
rect 22327 8041 22336 8075
rect 22284 8032 22336 8041
rect 27436 8032 27488 8084
rect 29092 8032 29144 8084
rect 34704 8075 34756 8084
rect 34704 8041 34713 8075
rect 34713 8041 34747 8075
rect 34747 8041 34756 8075
rect 34704 8032 34756 8041
rect 9312 7964 9364 8016
rect 9404 8007 9456 8016
rect 9404 7973 9413 8007
rect 9413 7973 9447 8007
rect 9447 7973 9456 8007
rect 9404 7964 9456 7973
rect 12256 7964 12308 8016
rect 16488 7964 16540 8016
rect 4712 7896 4764 7948
rect 1768 7871 1820 7880
rect 1768 7837 1777 7871
rect 1777 7837 1811 7871
rect 1811 7837 1820 7871
rect 1952 7871 2004 7880
rect 1768 7828 1820 7837
rect 1952 7837 1961 7871
rect 1961 7837 1995 7871
rect 1995 7837 2004 7871
rect 1952 7828 2004 7837
rect 3516 7828 3568 7880
rect 5448 7871 5500 7880
rect 2320 7760 2372 7812
rect 5080 7760 5132 7812
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 5448 7828 5500 7837
rect 6092 7871 6144 7880
rect 6092 7837 6101 7871
rect 6101 7837 6135 7871
rect 6135 7837 6144 7871
rect 6092 7828 6144 7837
rect 6184 7828 6236 7880
rect 6736 7828 6788 7880
rect 5632 7760 5684 7812
rect 7656 7828 7708 7880
rect 8116 7828 8168 7880
rect 8852 7760 8904 7812
rect 8944 7804 8996 7856
rect 9312 7828 9364 7880
rect 9404 7828 9456 7880
rect 9864 7896 9916 7948
rect 10140 7871 10192 7880
rect 10140 7837 10149 7871
rect 10149 7837 10183 7871
rect 10183 7837 10192 7871
rect 10140 7828 10192 7837
rect 10232 7871 10284 7880
rect 10232 7837 10241 7871
rect 10241 7837 10275 7871
rect 10275 7837 10284 7871
rect 10508 7871 10560 7880
rect 10232 7828 10284 7837
rect 10508 7837 10517 7871
rect 10517 7837 10551 7871
rect 10551 7837 10560 7871
rect 10508 7828 10560 7837
rect 9772 7760 9824 7812
rect 10692 7760 10744 7812
rect 11336 7828 11388 7880
rect 11612 7896 11664 7948
rect 12440 7939 12492 7948
rect 12440 7905 12449 7939
rect 12449 7905 12483 7939
rect 12483 7905 12492 7939
rect 12440 7896 12492 7905
rect 14464 7939 14516 7948
rect 12256 7871 12308 7880
rect 12256 7837 12265 7871
rect 12265 7837 12299 7871
rect 12299 7837 12308 7871
rect 12532 7871 12584 7880
rect 12256 7828 12308 7837
rect 12532 7837 12541 7871
rect 12541 7837 12575 7871
rect 12575 7837 12584 7871
rect 12532 7828 12584 7837
rect 12992 7828 13044 7880
rect 13360 7828 13412 7880
rect 13544 7871 13596 7880
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 14464 7905 14473 7939
rect 14473 7905 14507 7939
rect 14507 7905 14516 7939
rect 14464 7896 14516 7905
rect 13912 7828 13964 7880
rect 16304 7896 16356 7948
rect 20168 7964 20220 8016
rect 20720 7964 20772 8016
rect 21548 7964 21600 8016
rect 15108 7828 15160 7880
rect 16948 7828 17000 7880
rect 17500 7896 17552 7948
rect 18052 7871 18104 7880
rect 18052 7837 18061 7871
rect 18061 7837 18095 7871
rect 18095 7837 18104 7871
rect 18052 7828 18104 7837
rect 18236 7871 18288 7880
rect 18236 7837 18245 7871
rect 18245 7837 18279 7871
rect 18279 7837 18288 7871
rect 18236 7828 18288 7837
rect 19248 7828 19300 7880
rect 20444 7871 20496 7880
rect 20444 7837 20453 7871
rect 20453 7837 20487 7871
rect 20487 7837 20496 7871
rect 20444 7828 20496 7837
rect 22192 7896 22244 7948
rect 22928 7871 22980 7880
rect 22928 7837 22937 7871
rect 22937 7837 22971 7871
rect 22971 7837 22980 7871
rect 22928 7828 22980 7837
rect 23480 7896 23532 7948
rect 23664 7896 23716 7948
rect 4344 7692 4396 7744
rect 4804 7692 4856 7744
rect 5816 7692 5868 7744
rect 6460 7692 6512 7744
rect 8484 7692 8536 7744
rect 9588 7692 9640 7744
rect 10048 7692 10100 7744
rect 10140 7692 10192 7744
rect 15476 7760 15528 7812
rect 13728 7692 13780 7744
rect 17960 7760 18012 7812
rect 19432 7803 19484 7812
rect 19432 7769 19441 7803
rect 19441 7769 19475 7803
rect 19475 7769 19484 7803
rect 19432 7760 19484 7769
rect 16028 7692 16080 7744
rect 16580 7692 16632 7744
rect 17408 7692 17460 7744
rect 20352 7760 20404 7812
rect 22468 7760 22520 7812
rect 23940 7828 23992 7880
rect 25136 7871 25188 7880
rect 25136 7837 25145 7871
rect 25145 7837 25179 7871
rect 25179 7837 25188 7871
rect 25136 7828 25188 7837
rect 26608 7896 26660 7948
rect 25412 7828 25464 7880
rect 26700 7828 26752 7880
rect 20536 7692 20588 7744
rect 20720 7692 20772 7744
rect 24492 7760 24544 7812
rect 25044 7760 25096 7812
rect 27344 7896 27396 7948
rect 27620 7964 27672 8016
rect 28632 7964 28684 8016
rect 29000 7964 29052 8016
rect 29276 7896 29328 7948
rect 29460 7896 29512 7948
rect 27528 7871 27580 7880
rect 27528 7837 27537 7871
rect 27537 7837 27571 7871
rect 27571 7837 27580 7871
rect 27528 7828 27580 7837
rect 27620 7828 27672 7880
rect 28080 7760 28132 7812
rect 28264 7760 28316 7812
rect 30472 7828 30524 7880
rect 31024 7871 31076 7880
rect 31024 7837 31033 7871
rect 31033 7837 31067 7871
rect 31067 7837 31076 7871
rect 31024 7828 31076 7837
rect 31668 7871 31720 7880
rect 31668 7837 31677 7871
rect 31677 7837 31711 7871
rect 31711 7837 31720 7871
rect 31668 7828 31720 7837
rect 32956 7828 33008 7880
rect 29828 7760 29880 7812
rect 23756 7692 23808 7744
rect 25504 7692 25556 7744
rect 26700 7692 26752 7744
rect 28908 7692 28960 7744
rect 30380 7692 30432 7744
rect 32864 7760 32916 7812
rect 35164 7871 35216 7880
rect 35164 7837 35173 7871
rect 35173 7837 35207 7871
rect 35207 7837 35216 7871
rect 35164 7828 35216 7837
rect 33048 7692 33100 7744
rect 34704 7692 34756 7744
rect 35440 7692 35492 7744
rect 35624 7735 35676 7744
rect 35624 7701 35633 7735
rect 35633 7701 35667 7735
rect 35667 7701 35676 7735
rect 35624 7692 35676 7701
rect 36084 7692 36136 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 1768 7488 1820 7540
rect 2320 7531 2372 7540
rect 2320 7497 2329 7531
rect 2329 7497 2363 7531
rect 2363 7497 2372 7531
rect 2320 7488 2372 7497
rect 2964 7531 3016 7540
rect 940 7352 992 7404
rect 2964 7497 2973 7531
rect 2973 7497 3007 7531
rect 3007 7497 3016 7531
rect 2964 7488 3016 7497
rect 4068 7488 4120 7540
rect 5816 7488 5868 7540
rect 3884 7395 3936 7404
rect 3884 7361 3918 7395
rect 3918 7361 3936 7395
rect 4344 7420 4396 7472
rect 6184 7420 6236 7472
rect 8484 7463 8536 7472
rect 3884 7352 3936 7361
rect 3608 7327 3660 7336
rect 3608 7293 3617 7327
rect 3617 7293 3651 7327
rect 3651 7293 3660 7327
rect 3608 7284 3660 7293
rect 4804 7352 4856 7404
rect 6368 7395 6420 7404
rect 6368 7361 6377 7395
rect 6377 7361 6411 7395
rect 6411 7361 6420 7395
rect 6368 7352 6420 7361
rect 6460 7352 6512 7404
rect 8484 7429 8518 7463
rect 8518 7429 8536 7463
rect 8484 7420 8536 7429
rect 9496 7488 9548 7540
rect 10048 7488 10100 7540
rect 10416 7488 10468 7540
rect 4620 7216 4672 7268
rect 5264 7216 5316 7268
rect 5448 7148 5500 7200
rect 8116 7284 8168 7336
rect 9496 7352 9548 7404
rect 10140 7352 10192 7404
rect 10968 7352 11020 7404
rect 15108 7488 15160 7540
rect 15476 7531 15528 7540
rect 15476 7497 15485 7531
rect 15485 7497 15519 7531
rect 15519 7497 15528 7531
rect 15476 7488 15528 7497
rect 18236 7488 18288 7540
rect 18604 7488 18656 7540
rect 12348 7420 12400 7472
rect 9772 7284 9824 7336
rect 12440 7352 12492 7404
rect 13084 7352 13136 7404
rect 9404 7216 9456 7268
rect 13452 7284 13504 7336
rect 15752 7395 15804 7404
rect 15752 7361 15761 7395
rect 15761 7361 15795 7395
rect 15795 7361 15804 7395
rect 16028 7395 16080 7404
rect 15752 7352 15804 7361
rect 16028 7361 16037 7395
rect 16037 7361 16071 7395
rect 16071 7361 16080 7395
rect 16028 7352 16080 7361
rect 16580 7352 16632 7404
rect 17132 7352 17184 7404
rect 20352 7488 20404 7540
rect 22376 7531 22428 7540
rect 22376 7497 22385 7531
rect 22385 7497 22419 7531
rect 22419 7497 22428 7531
rect 22376 7488 22428 7497
rect 22744 7488 22796 7540
rect 27344 7488 27396 7540
rect 24032 7420 24084 7472
rect 24216 7420 24268 7472
rect 20904 7395 20956 7404
rect 20904 7361 20913 7395
rect 20913 7361 20947 7395
rect 20947 7361 20956 7395
rect 20904 7352 20956 7361
rect 22100 7352 22152 7404
rect 23020 7395 23072 7404
rect 23020 7361 23029 7395
rect 23029 7361 23063 7395
rect 23063 7361 23072 7395
rect 23020 7352 23072 7361
rect 23664 7395 23716 7404
rect 23664 7361 23673 7395
rect 23673 7361 23707 7395
rect 23707 7361 23716 7395
rect 23664 7352 23716 7361
rect 24308 7395 24360 7404
rect 24308 7361 24317 7395
rect 24317 7361 24351 7395
rect 24351 7361 24360 7395
rect 24308 7352 24360 7361
rect 24492 7420 24544 7472
rect 24768 7352 24820 7404
rect 25320 7395 25372 7404
rect 25320 7361 25329 7395
rect 25329 7361 25363 7395
rect 25363 7361 25372 7395
rect 25320 7352 25372 7361
rect 25964 7395 26016 7404
rect 25964 7361 25973 7395
rect 25973 7361 26007 7395
rect 26007 7361 26016 7395
rect 25964 7352 26016 7361
rect 27068 7352 27120 7404
rect 28080 7420 28132 7472
rect 29276 7488 29328 7540
rect 30840 7531 30892 7540
rect 30840 7497 30849 7531
rect 30849 7497 30883 7531
rect 30883 7497 30892 7531
rect 30840 7488 30892 7497
rect 32864 7531 32916 7540
rect 32864 7497 32873 7531
rect 32873 7497 32907 7531
rect 32907 7497 32916 7531
rect 32864 7488 32916 7497
rect 34704 7488 34756 7540
rect 36084 7488 36136 7540
rect 29184 7395 29236 7404
rect 29184 7361 29193 7395
rect 29193 7361 29227 7395
rect 29227 7361 29236 7395
rect 32772 7420 32824 7472
rect 29184 7352 29236 7361
rect 16120 7284 16172 7336
rect 17408 7284 17460 7336
rect 6552 7148 6604 7200
rect 6644 7148 6696 7200
rect 9220 7148 9272 7200
rect 10692 7148 10744 7200
rect 14924 7216 14976 7268
rect 20444 7284 20496 7336
rect 23940 7284 23992 7336
rect 28080 7284 28132 7336
rect 28908 7284 28960 7336
rect 20260 7216 20312 7268
rect 24400 7216 24452 7268
rect 31208 7352 31260 7404
rect 30196 7284 30248 7336
rect 32496 7352 32548 7404
rect 33048 7395 33100 7404
rect 33048 7361 33057 7395
rect 33057 7361 33091 7395
rect 33091 7361 33100 7395
rect 33048 7352 33100 7361
rect 35624 7420 35676 7472
rect 35164 7352 35216 7404
rect 35716 7352 35768 7404
rect 36452 7395 36504 7404
rect 36452 7361 36461 7395
rect 36461 7361 36495 7395
rect 36495 7361 36504 7395
rect 36452 7352 36504 7361
rect 32956 7284 33008 7336
rect 31944 7216 31996 7268
rect 34796 7216 34848 7268
rect 13268 7191 13320 7200
rect 13268 7157 13277 7191
rect 13277 7157 13311 7191
rect 13311 7157 13320 7191
rect 13268 7148 13320 7157
rect 13452 7148 13504 7200
rect 15660 7148 15712 7200
rect 23204 7148 23256 7200
rect 24124 7191 24176 7200
rect 24124 7157 24133 7191
rect 24133 7157 24167 7191
rect 24167 7157 24176 7191
rect 24124 7148 24176 7157
rect 24952 7148 25004 7200
rect 29184 7148 29236 7200
rect 32128 7148 32180 7200
rect 33416 7148 33468 7200
rect 35440 7148 35492 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 2136 6944 2188 6996
rect 2964 6944 3016 6996
rect 3056 6808 3108 6860
rect 2964 6740 3016 6792
rect 3608 6808 3660 6860
rect 5632 6851 5684 6860
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 5632 6808 5684 6817
rect 4068 6783 4120 6792
rect 4068 6749 4102 6783
rect 4102 6749 4120 6783
rect 4068 6740 4120 6749
rect 6000 6808 6052 6860
rect 7656 6876 7708 6928
rect 9220 6987 9272 6996
rect 9220 6953 9229 6987
rect 9229 6953 9263 6987
rect 9263 6953 9272 6987
rect 9220 6944 9272 6953
rect 9404 6987 9456 6996
rect 9404 6953 9413 6987
rect 9413 6953 9447 6987
rect 9447 6953 9456 6987
rect 9404 6944 9456 6953
rect 12256 6944 12308 6996
rect 14004 6944 14056 6996
rect 12348 6876 12400 6928
rect 12808 6876 12860 6928
rect 7564 6808 7616 6860
rect 6184 6783 6236 6792
rect 4528 6672 4580 6724
rect 6184 6749 6193 6783
rect 6193 6749 6227 6783
rect 6227 6749 6236 6783
rect 6184 6740 6236 6749
rect 6828 6740 6880 6792
rect 8208 6740 8260 6792
rect 8668 6740 8720 6792
rect 8760 6740 8812 6792
rect 16028 6944 16080 6996
rect 16304 6944 16356 6996
rect 16672 6944 16724 6996
rect 18052 6876 18104 6928
rect 18788 6876 18840 6928
rect 7932 6672 7984 6724
rect 9036 6672 9088 6724
rect 9404 6740 9456 6792
rect 15200 6808 15252 6860
rect 21732 6944 21784 6996
rect 25964 6944 26016 6996
rect 29184 6944 29236 6996
rect 34612 6944 34664 6996
rect 24032 6876 24084 6928
rect 24400 6876 24452 6928
rect 24676 6876 24728 6928
rect 24952 6876 25004 6928
rect 25044 6876 25096 6928
rect 29460 6876 29512 6928
rect 11980 6740 12032 6792
rect 12992 6783 13044 6792
rect 12992 6749 13001 6783
rect 13001 6749 13035 6783
rect 13035 6749 13044 6783
rect 12992 6740 13044 6749
rect 13176 6740 13228 6792
rect 13544 6740 13596 6792
rect 16120 6783 16172 6792
rect 16120 6749 16129 6783
rect 16129 6749 16163 6783
rect 16163 6749 16172 6783
rect 16120 6740 16172 6749
rect 21456 6808 21508 6860
rect 24308 6808 24360 6860
rect 16488 6783 16540 6792
rect 16488 6749 16497 6783
rect 16497 6749 16531 6783
rect 16531 6749 16540 6783
rect 16488 6740 16540 6749
rect 10600 6715 10652 6724
rect 10600 6681 10634 6715
rect 10634 6681 10652 6715
rect 10600 6672 10652 6681
rect 10876 6672 10928 6724
rect 5632 6604 5684 6656
rect 6460 6604 6512 6656
rect 9588 6604 9640 6656
rect 10692 6604 10744 6656
rect 12164 6672 12216 6724
rect 14556 6672 14608 6724
rect 14740 6672 14792 6724
rect 17868 6740 17920 6792
rect 19064 6740 19116 6792
rect 19340 6740 19392 6792
rect 20628 6740 20680 6792
rect 21824 6783 21876 6792
rect 21824 6749 21833 6783
rect 21833 6749 21867 6783
rect 21867 6749 21876 6783
rect 21824 6740 21876 6749
rect 23756 6740 23808 6792
rect 24492 6740 24544 6792
rect 24768 6740 24820 6792
rect 29092 6808 29144 6860
rect 25596 6783 25648 6792
rect 25596 6749 25605 6783
rect 25605 6749 25639 6783
rect 25639 6749 25648 6783
rect 25596 6740 25648 6749
rect 26148 6740 26200 6792
rect 26332 6740 26384 6792
rect 28080 6783 28132 6792
rect 28080 6749 28089 6783
rect 28089 6749 28123 6783
rect 28123 6749 28132 6783
rect 28080 6740 28132 6749
rect 20168 6715 20220 6724
rect 15108 6604 15160 6656
rect 15200 6604 15252 6656
rect 15936 6647 15988 6656
rect 15936 6613 15945 6647
rect 15945 6613 15979 6647
rect 15979 6613 15988 6647
rect 15936 6604 15988 6613
rect 16304 6604 16356 6656
rect 20168 6681 20202 6715
rect 20202 6681 20220 6715
rect 20168 6672 20220 6681
rect 23296 6672 23348 6724
rect 20720 6604 20772 6656
rect 21272 6647 21324 6656
rect 21272 6613 21281 6647
rect 21281 6613 21315 6647
rect 21315 6613 21324 6647
rect 21272 6604 21324 6613
rect 21364 6604 21416 6656
rect 23388 6604 23440 6656
rect 25136 6672 25188 6724
rect 24400 6647 24452 6656
rect 24400 6613 24409 6647
rect 24409 6613 24443 6647
rect 24443 6613 24452 6647
rect 24400 6604 24452 6613
rect 25228 6604 25280 6656
rect 26516 6672 26568 6724
rect 28540 6715 28592 6724
rect 28540 6681 28549 6715
rect 28549 6681 28583 6715
rect 28583 6681 28592 6715
rect 28540 6672 28592 6681
rect 29276 6740 29328 6792
rect 29736 6783 29788 6792
rect 29736 6749 29745 6783
rect 29745 6749 29779 6783
rect 29779 6749 29788 6783
rect 29736 6740 29788 6749
rect 26424 6604 26476 6656
rect 29828 6672 29880 6724
rect 30012 6715 30064 6724
rect 30012 6681 30046 6715
rect 30046 6681 30064 6715
rect 30012 6672 30064 6681
rect 31760 6783 31812 6792
rect 31760 6749 31769 6783
rect 31769 6749 31803 6783
rect 31803 6749 31812 6783
rect 31760 6740 31812 6749
rect 32128 6672 32180 6724
rect 32496 6808 32548 6860
rect 37556 6808 37608 6860
rect 32312 6740 32364 6792
rect 32772 6740 32824 6792
rect 34060 6783 34112 6792
rect 34060 6749 34069 6783
rect 34069 6749 34103 6783
rect 34103 6749 34112 6783
rect 34060 6740 34112 6749
rect 35808 6783 35860 6792
rect 35808 6749 35817 6783
rect 35817 6749 35851 6783
rect 35851 6749 35860 6783
rect 35808 6740 35860 6749
rect 33508 6672 33560 6724
rect 34704 6715 34756 6724
rect 34704 6681 34713 6715
rect 34713 6681 34747 6715
rect 34747 6681 34756 6715
rect 34704 6672 34756 6681
rect 30472 6604 30524 6656
rect 31208 6604 31260 6656
rect 32864 6604 32916 6656
rect 33876 6604 33928 6656
rect 34888 6647 34940 6656
rect 34888 6613 34913 6647
rect 34913 6613 34940 6647
rect 34888 6604 34940 6613
rect 37648 6604 37700 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 1768 6443 1820 6452
rect 1768 6409 1777 6443
rect 1777 6409 1811 6443
rect 1811 6409 1820 6443
rect 1768 6400 1820 6409
rect 3884 6400 3936 6452
rect 3976 6400 4028 6452
rect 4712 6400 4764 6452
rect 6092 6400 6144 6452
rect 4436 6332 4488 6384
rect 3884 6307 3936 6316
rect 2780 6196 2832 6248
rect 3884 6273 3893 6307
rect 3893 6273 3927 6307
rect 3927 6273 3936 6307
rect 3884 6264 3936 6273
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 4804 6264 4856 6316
rect 5540 6264 5592 6316
rect 7288 6332 7340 6384
rect 7380 6332 7432 6384
rect 8484 6332 8536 6384
rect 8944 6332 8996 6384
rect 9496 6400 9548 6452
rect 10140 6400 10192 6452
rect 10600 6443 10652 6452
rect 10600 6409 10609 6443
rect 10609 6409 10643 6443
rect 10643 6409 10652 6443
rect 10600 6400 10652 6409
rect 10692 6400 10744 6452
rect 6644 6307 6696 6316
rect 6644 6273 6653 6307
rect 6653 6273 6687 6307
rect 6687 6273 6696 6307
rect 6644 6264 6696 6273
rect 5816 6196 5868 6248
rect 7012 6264 7064 6316
rect 8668 6264 8720 6316
rect 8392 6196 8444 6248
rect 8852 6196 8904 6248
rect 10232 6332 10284 6384
rect 12716 6400 12768 6452
rect 12992 6400 13044 6452
rect 15108 6400 15160 6452
rect 16488 6400 16540 6452
rect 9956 6264 10008 6316
rect 10508 6264 10560 6316
rect 10784 6307 10836 6316
rect 10784 6273 10793 6307
rect 10793 6273 10827 6307
rect 10827 6273 10836 6307
rect 10784 6264 10836 6273
rect 11704 6264 11756 6316
rect 13176 6332 13228 6384
rect 15292 6332 15344 6384
rect 24676 6400 24728 6452
rect 18880 6332 18932 6384
rect 19248 6332 19300 6384
rect 20168 6332 20220 6384
rect 21180 6332 21232 6384
rect 31852 6400 31904 6452
rect 36452 6400 36504 6452
rect 12348 6264 12400 6316
rect 12992 6307 13044 6316
rect 12992 6273 13001 6307
rect 13001 6273 13035 6307
rect 13035 6273 13044 6307
rect 12992 6264 13044 6273
rect 13268 6264 13320 6316
rect 14096 6307 14148 6316
rect 11612 6239 11664 6248
rect 11612 6205 11621 6239
rect 11621 6205 11655 6239
rect 11655 6205 11664 6239
rect 11612 6196 11664 6205
rect 14096 6273 14105 6307
rect 14105 6273 14139 6307
rect 14139 6273 14148 6307
rect 14096 6264 14148 6273
rect 14740 6307 14792 6316
rect 14740 6273 14749 6307
rect 14749 6273 14783 6307
rect 14783 6273 14792 6307
rect 14740 6264 14792 6273
rect 15016 6307 15068 6316
rect 15016 6273 15050 6307
rect 15050 6273 15068 6307
rect 15016 6264 15068 6273
rect 17224 6264 17276 6316
rect 19984 6264 20036 6316
rect 20444 6307 20496 6316
rect 20444 6273 20453 6307
rect 20453 6273 20487 6307
rect 20487 6273 20496 6307
rect 20444 6264 20496 6273
rect 2412 6060 2464 6112
rect 2872 6128 2924 6180
rect 3332 6060 3384 6112
rect 4068 6060 4120 6112
rect 5540 6060 5592 6112
rect 6828 6103 6880 6112
rect 6828 6069 6837 6103
rect 6837 6069 6871 6103
rect 6871 6069 6880 6103
rect 6828 6060 6880 6069
rect 7748 6060 7800 6112
rect 9588 6060 9640 6112
rect 10048 6103 10100 6112
rect 10048 6069 10057 6103
rect 10057 6069 10091 6103
rect 10091 6069 10100 6103
rect 10048 6060 10100 6069
rect 10232 6128 10284 6180
rect 13820 6196 13872 6248
rect 16120 6196 16172 6248
rect 17684 6196 17736 6248
rect 11980 6171 12032 6180
rect 11980 6137 11989 6171
rect 11989 6137 12023 6171
rect 12023 6137 12032 6171
rect 11980 6128 12032 6137
rect 11428 6060 11480 6112
rect 11520 6103 11572 6112
rect 11520 6069 11529 6103
rect 11529 6069 11563 6103
rect 11563 6069 11572 6103
rect 11520 6060 11572 6069
rect 13360 6060 13412 6112
rect 13912 6060 13964 6112
rect 16120 6103 16172 6112
rect 16120 6069 16129 6103
rect 16129 6069 16163 6103
rect 16163 6069 16172 6103
rect 16120 6060 16172 6069
rect 19248 6196 19300 6248
rect 21640 6264 21692 6316
rect 21824 6264 21876 6316
rect 22284 6307 22336 6316
rect 22284 6273 22293 6307
rect 22293 6273 22327 6307
rect 22327 6273 22336 6307
rect 22284 6264 22336 6273
rect 22836 6264 22888 6316
rect 24308 6307 24360 6316
rect 21456 6196 21508 6248
rect 24308 6273 24317 6307
rect 24317 6273 24351 6307
rect 24351 6273 24360 6307
rect 24308 6264 24360 6273
rect 26240 6332 26292 6384
rect 25504 6264 25556 6316
rect 27068 6264 27120 6316
rect 27528 6264 27580 6316
rect 29000 6264 29052 6316
rect 29736 6332 29788 6384
rect 29828 6332 29880 6384
rect 30380 6264 30432 6316
rect 24860 6196 24912 6248
rect 32956 6332 33008 6384
rect 32404 6307 32456 6316
rect 32404 6273 32438 6307
rect 32438 6273 32456 6307
rect 32404 6264 32456 6273
rect 34796 6332 34848 6384
rect 32128 6239 32180 6248
rect 19156 6128 19208 6180
rect 23480 6128 23532 6180
rect 19340 6060 19392 6112
rect 19616 6060 19668 6112
rect 24768 6128 24820 6180
rect 32128 6205 32137 6239
rect 32137 6205 32171 6239
rect 32171 6205 32180 6239
rect 32128 6196 32180 6205
rect 26148 6128 26200 6180
rect 27252 6060 27304 6112
rect 35900 6332 35952 6384
rect 37280 6264 37332 6316
rect 27804 6060 27856 6112
rect 28540 6060 28592 6112
rect 29460 6060 29512 6112
rect 31852 6060 31904 6112
rect 33048 6060 33100 6112
rect 35348 6103 35400 6112
rect 35348 6069 35357 6103
rect 35357 6069 35391 6103
rect 35391 6069 35400 6103
rect 35348 6060 35400 6069
rect 35992 6103 36044 6112
rect 35992 6069 36001 6103
rect 36001 6069 36035 6103
rect 36035 6069 36044 6103
rect 35992 6060 36044 6069
rect 37924 6060 37976 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 3884 5856 3936 5908
rect 4620 5856 4672 5908
rect 7748 5856 7800 5908
rect 8208 5856 8260 5908
rect 11888 5856 11940 5908
rect 12256 5856 12308 5908
rect 12348 5856 12400 5908
rect 15292 5856 15344 5908
rect 15752 5856 15804 5908
rect 16120 5856 16172 5908
rect 16580 5899 16632 5908
rect 16580 5865 16589 5899
rect 16589 5865 16623 5899
rect 16623 5865 16632 5899
rect 16580 5856 16632 5865
rect 10232 5788 10284 5840
rect 11704 5788 11756 5840
rect 12164 5831 12216 5840
rect 12164 5797 12173 5831
rect 12173 5797 12207 5831
rect 12207 5797 12216 5831
rect 12164 5788 12216 5797
rect 12900 5788 12952 5840
rect 14004 5788 14056 5840
rect 6184 5720 6236 5772
rect 6276 5720 6328 5772
rect 1768 5695 1820 5704
rect 1768 5661 1777 5695
rect 1777 5661 1811 5695
rect 1811 5661 1820 5695
rect 1768 5652 1820 5661
rect 2596 5695 2648 5704
rect 2596 5661 2605 5695
rect 2605 5661 2639 5695
rect 2639 5661 2648 5695
rect 2596 5652 2648 5661
rect 4160 5695 4212 5704
rect 4160 5661 4169 5695
rect 4169 5661 4203 5695
rect 4203 5661 4212 5695
rect 4160 5652 4212 5661
rect 3056 5516 3108 5568
rect 5080 5584 5132 5636
rect 6092 5584 6144 5636
rect 5908 5516 5960 5568
rect 6460 5584 6512 5636
rect 8944 5652 8996 5704
rect 7012 5516 7064 5568
rect 7288 5559 7340 5568
rect 7288 5525 7297 5559
rect 7297 5525 7331 5559
rect 7331 5525 7340 5559
rect 7288 5516 7340 5525
rect 9772 5652 9824 5704
rect 9956 5652 10008 5704
rect 11520 5720 11572 5772
rect 11796 5763 11848 5772
rect 11796 5729 11805 5763
rect 11805 5729 11839 5763
rect 11839 5729 11848 5763
rect 11796 5720 11848 5729
rect 11244 5695 11296 5704
rect 11244 5661 11253 5695
rect 11253 5661 11287 5695
rect 11287 5661 11296 5695
rect 11244 5652 11296 5661
rect 11336 5652 11388 5704
rect 12808 5720 12860 5772
rect 15108 5720 15160 5772
rect 15292 5763 15344 5772
rect 15292 5729 15301 5763
rect 15301 5729 15335 5763
rect 15335 5729 15344 5763
rect 15292 5720 15344 5729
rect 13636 5652 13688 5704
rect 10876 5516 10928 5568
rect 14004 5584 14056 5636
rect 12900 5516 12952 5568
rect 13268 5516 13320 5568
rect 13728 5516 13780 5568
rect 16672 5720 16724 5772
rect 18052 5856 18104 5908
rect 18420 5856 18472 5908
rect 19156 5856 19208 5908
rect 19432 5856 19484 5908
rect 17132 5788 17184 5840
rect 16488 5652 16540 5704
rect 18604 5763 18656 5772
rect 18604 5729 18613 5763
rect 18613 5729 18647 5763
rect 18647 5729 18656 5763
rect 18604 5720 18656 5729
rect 19616 5856 19668 5908
rect 20904 5856 20956 5908
rect 23848 5899 23900 5908
rect 23848 5865 23857 5899
rect 23857 5865 23891 5899
rect 23891 5865 23900 5899
rect 23848 5856 23900 5865
rect 26608 5899 26660 5908
rect 26608 5865 26617 5899
rect 26617 5865 26651 5899
rect 26651 5865 26660 5899
rect 26608 5856 26660 5865
rect 26884 5856 26936 5908
rect 30748 5856 30800 5908
rect 33416 5899 33468 5908
rect 33416 5865 33425 5899
rect 33425 5865 33459 5899
rect 33459 5865 33468 5899
rect 33416 5856 33468 5865
rect 33600 5899 33652 5908
rect 33600 5865 33609 5899
rect 33609 5865 33643 5899
rect 33643 5865 33652 5899
rect 33600 5856 33652 5865
rect 34612 5856 34664 5908
rect 35808 5856 35860 5908
rect 15200 5627 15252 5636
rect 15200 5593 15209 5627
rect 15209 5593 15243 5627
rect 15243 5593 15252 5627
rect 15200 5584 15252 5593
rect 16304 5627 16356 5636
rect 16304 5593 16313 5627
rect 16313 5593 16347 5627
rect 16347 5593 16356 5627
rect 16304 5584 16356 5593
rect 17684 5652 17736 5704
rect 18420 5695 18472 5704
rect 18420 5661 18429 5695
rect 18429 5661 18463 5695
rect 18463 5661 18472 5695
rect 18420 5652 18472 5661
rect 21272 5788 21324 5840
rect 21456 5831 21508 5840
rect 21456 5797 21465 5831
rect 21465 5797 21499 5831
rect 21499 5797 21508 5831
rect 21456 5788 21508 5797
rect 24952 5788 25004 5840
rect 29000 5788 29052 5840
rect 29276 5788 29328 5840
rect 34428 5788 34480 5840
rect 35992 5788 36044 5840
rect 37372 5788 37424 5840
rect 19984 5720 20036 5772
rect 20444 5652 20496 5704
rect 20720 5652 20772 5704
rect 21364 5652 21416 5704
rect 21916 5652 21968 5704
rect 28264 5720 28316 5772
rect 28356 5720 28408 5772
rect 29552 5720 29604 5772
rect 31944 5763 31996 5772
rect 31944 5729 31953 5763
rect 31953 5729 31987 5763
rect 31987 5729 31996 5763
rect 31944 5720 31996 5729
rect 32036 5720 32088 5772
rect 32312 5720 32364 5772
rect 34060 5720 34112 5772
rect 35808 5720 35860 5772
rect 22100 5627 22152 5636
rect 22100 5593 22109 5627
rect 22109 5593 22143 5627
rect 22143 5593 22152 5627
rect 22100 5584 22152 5593
rect 22652 5695 22704 5704
rect 22652 5661 22661 5695
rect 22661 5661 22695 5695
rect 22695 5661 22704 5695
rect 22652 5652 22704 5661
rect 24124 5652 24176 5704
rect 24400 5695 24452 5704
rect 24400 5661 24409 5695
rect 24409 5661 24443 5695
rect 24443 5661 24452 5695
rect 24400 5652 24452 5661
rect 26240 5652 26292 5704
rect 27712 5652 27764 5704
rect 23296 5584 23348 5636
rect 23388 5584 23440 5636
rect 24308 5584 24360 5636
rect 24768 5627 24820 5636
rect 24768 5593 24777 5627
rect 24777 5593 24811 5627
rect 24811 5593 24820 5627
rect 24768 5584 24820 5593
rect 26700 5584 26752 5636
rect 15108 5516 15160 5568
rect 16948 5559 17000 5568
rect 16948 5525 16957 5559
rect 16957 5525 16991 5559
rect 16991 5525 17000 5559
rect 16948 5516 17000 5525
rect 18144 5559 18196 5568
rect 18144 5525 18153 5559
rect 18153 5525 18187 5559
rect 18187 5525 18196 5559
rect 18144 5516 18196 5525
rect 18604 5516 18656 5568
rect 19984 5516 20036 5568
rect 21824 5516 21876 5568
rect 22376 5516 22428 5568
rect 29736 5652 29788 5704
rect 30380 5627 30432 5636
rect 30380 5593 30414 5627
rect 30414 5593 30432 5627
rect 30380 5584 30432 5593
rect 32128 5584 32180 5636
rect 28908 5516 28960 5568
rect 30012 5516 30064 5568
rect 30288 5516 30340 5568
rect 31576 5516 31628 5568
rect 34152 5652 34204 5704
rect 36912 5652 36964 5704
rect 37096 5695 37148 5704
rect 37096 5661 37105 5695
rect 37105 5661 37139 5695
rect 37139 5661 37148 5695
rect 37096 5652 37148 5661
rect 37740 5695 37792 5704
rect 37740 5661 37749 5695
rect 37749 5661 37783 5695
rect 37783 5661 37792 5695
rect 37740 5652 37792 5661
rect 32404 5584 32456 5636
rect 33048 5584 33100 5636
rect 32956 5516 33008 5568
rect 34612 5584 34664 5636
rect 35348 5584 35400 5636
rect 34520 5516 34572 5568
rect 34796 5516 34848 5568
rect 35532 5559 35584 5568
rect 35532 5525 35541 5559
rect 35541 5525 35575 5559
rect 35575 5525 35584 5559
rect 35532 5516 35584 5525
rect 37464 5516 37516 5568
rect 37832 5516 37884 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 3056 5312 3108 5364
rect 4620 5312 4672 5364
rect 5080 5312 5132 5364
rect 5356 5312 5408 5364
rect 2872 5244 2924 5296
rect 5632 5312 5684 5364
rect 6920 5312 6972 5364
rect 7932 5312 7984 5364
rect 8024 5312 8076 5364
rect 9772 5312 9824 5364
rect 10324 5312 10376 5364
rect 2780 5176 2832 5228
rect 3424 5176 3476 5228
rect 3700 5176 3752 5228
rect 4620 5176 4672 5228
rect 5632 5185 5649 5212
rect 5649 5185 5683 5212
rect 5683 5185 5684 5212
rect 5632 5160 5684 5185
rect 7104 5244 7156 5296
rect 6460 5176 6512 5228
rect 5816 5108 5868 5160
rect 10048 5244 10100 5296
rect 10968 5312 11020 5364
rect 11336 5312 11388 5364
rect 11060 5244 11112 5296
rect 15108 5312 15160 5364
rect 17500 5312 17552 5364
rect 18972 5312 19024 5364
rect 20352 5312 20404 5364
rect 24216 5312 24268 5364
rect 24860 5312 24912 5364
rect 16948 5244 17000 5296
rect 18144 5287 18196 5296
rect 18144 5253 18153 5287
rect 18153 5253 18187 5287
rect 18187 5253 18196 5287
rect 18144 5244 18196 5253
rect 20260 5244 20312 5296
rect 23572 5287 23624 5296
rect 23572 5253 23606 5287
rect 23606 5253 23624 5287
rect 23572 5244 23624 5253
rect 27896 5312 27948 5364
rect 7380 5219 7432 5228
rect 7380 5185 7389 5219
rect 7389 5185 7423 5219
rect 7423 5185 7432 5219
rect 7380 5176 7432 5185
rect 8024 5176 8076 5228
rect 9128 5176 9180 5228
rect 9588 5219 9640 5228
rect 9588 5185 9597 5219
rect 9597 5185 9631 5219
rect 9631 5185 9640 5219
rect 9588 5176 9640 5185
rect 7472 5151 7524 5160
rect 7472 5117 7481 5151
rect 7481 5117 7515 5151
rect 7515 5117 7524 5151
rect 7472 5108 7524 5117
rect 10232 5176 10284 5228
rect 10508 5219 10560 5228
rect 10508 5185 10517 5219
rect 10517 5185 10551 5219
rect 10551 5185 10560 5219
rect 10508 5176 10560 5185
rect 10876 5176 10928 5228
rect 3608 5040 3660 5092
rect 2320 5015 2372 5024
rect 2320 4981 2329 5015
rect 2329 4981 2363 5015
rect 2363 4981 2372 5015
rect 2320 4972 2372 4981
rect 4988 4972 5040 5024
rect 5264 4972 5316 5024
rect 9772 5040 9824 5092
rect 10600 5040 10652 5092
rect 6000 4972 6052 5024
rect 7656 5015 7708 5024
rect 7656 4981 7665 5015
rect 7665 4981 7699 5015
rect 7699 4981 7708 5015
rect 7656 4972 7708 4981
rect 8944 4972 8996 5024
rect 9220 4972 9272 5024
rect 9588 4972 9640 5024
rect 10692 4972 10744 5024
rect 10968 5108 11020 5160
rect 12164 5176 12216 5228
rect 12808 5108 12860 5160
rect 13268 5176 13320 5228
rect 14648 5176 14700 5228
rect 15568 5176 15620 5228
rect 15844 5219 15896 5228
rect 15844 5185 15853 5219
rect 15853 5185 15887 5219
rect 15887 5185 15896 5219
rect 15844 5176 15896 5185
rect 17408 5176 17460 5228
rect 19340 5219 19392 5228
rect 19340 5185 19349 5219
rect 19349 5185 19383 5219
rect 19383 5185 19392 5219
rect 19340 5176 19392 5185
rect 21824 5219 21876 5228
rect 21824 5185 21833 5219
rect 21833 5185 21867 5219
rect 21867 5185 21876 5219
rect 21824 5176 21876 5185
rect 24676 5176 24728 5228
rect 26608 5244 26660 5296
rect 29460 5312 29512 5364
rect 30380 5355 30432 5364
rect 30380 5321 30389 5355
rect 30389 5321 30423 5355
rect 30423 5321 30432 5355
rect 30380 5312 30432 5321
rect 22284 5108 22336 5160
rect 24952 5108 25004 5160
rect 25780 5176 25832 5228
rect 27344 5176 27396 5228
rect 29000 5287 29052 5296
rect 29000 5253 29025 5287
rect 29025 5253 29052 5287
rect 34520 5312 34572 5364
rect 37280 5312 37332 5364
rect 29000 5244 29052 5253
rect 31576 5244 31628 5296
rect 29276 5176 29328 5228
rect 25872 5108 25924 5160
rect 27712 5108 27764 5160
rect 28724 5108 28776 5160
rect 30288 5176 30340 5228
rect 32496 5244 32548 5296
rect 34612 5287 34664 5296
rect 30196 5108 30248 5160
rect 32772 5176 32824 5228
rect 33416 5176 33468 5228
rect 34612 5253 34653 5287
rect 34653 5253 34664 5287
rect 34612 5244 34664 5253
rect 35900 5244 35952 5296
rect 34796 5176 34848 5228
rect 35348 5176 35400 5228
rect 34520 5108 34572 5160
rect 36268 5176 36320 5228
rect 37648 5176 37700 5228
rect 18604 5040 18656 5092
rect 24400 5040 24452 5092
rect 11336 4972 11388 5024
rect 12440 4972 12492 5024
rect 14004 4972 14056 5024
rect 14280 4972 14332 5024
rect 15200 4972 15252 5024
rect 15384 4972 15436 5024
rect 20904 4972 20956 5024
rect 22192 4972 22244 5024
rect 23940 4972 23992 5024
rect 24216 4972 24268 5024
rect 26056 5040 26108 5092
rect 31024 5040 31076 5092
rect 34704 5040 34756 5092
rect 27620 5015 27672 5024
rect 27620 4981 27629 5015
rect 27629 4981 27663 5015
rect 27663 4981 27672 5015
rect 27620 4972 27672 4981
rect 29092 4972 29144 5024
rect 29552 4972 29604 5024
rect 29736 4972 29788 5024
rect 31392 4972 31444 5024
rect 32220 4972 32272 5024
rect 33324 5015 33376 5024
rect 33324 4981 33333 5015
rect 33333 4981 33367 5015
rect 33367 4981 33376 5015
rect 33324 4972 33376 4981
rect 34428 4972 34480 5024
rect 35900 5015 35952 5024
rect 35900 4981 35909 5015
rect 35909 4981 35943 5015
rect 35943 4981 35952 5015
rect 35900 4972 35952 4981
rect 37280 4972 37332 5024
rect 39764 4972 39816 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 2320 4768 2372 4820
rect 3056 4743 3108 4752
rect 2688 4632 2740 4684
rect 3056 4709 3065 4743
rect 3065 4709 3099 4743
rect 3099 4709 3108 4743
rect 3056 4700 3108 4709
rect 4160 4700 4212 4752
rect 5632 4768 5684 4820
rect 7012 4768 7064 4820
rect 7932 4768 7984 4820
rect 8116 4811 8168 4820
rect 8116 4777 8125 4811
rect 8125 4777 8159 4811
rect 8159 4777 8168 4811
rect 8116 4768 8168 4777
rect 8208 4768 8260 4820
rect 9312 4768 9364 4820
rect 11796 4811 11848 4820
rect 11796 4777 11805 4811
rect 11805 4777 11839 4811
rect 11839 4777 11848 4811
rect 11796 4768 11848 4777
rect 14648 4811 14700 4820
rect 14648 4777 14657 4811
rect 14657 4777 14691 4811
rect 14691 4777 14700 4811
rect 14648 4768 14700 4777
rect 18604 4811 18656 4820
rect 18604 4777 18613 4811
rect 18613 4777 18647 4811
rect 18647 4777 18656 4811
rect 18604 4768 18656 4777
rect 21732 4768 21784 4820
rect 22100 4768 22152 4820
rect 22468 4768 22520 4820
rect 22652 4768 22704 4820
rect 28448 4768 28500 4820
rect 29736 4811 29788 4820
rect 29736 4777 29745 4811
rect 29745 4777 29779 4811
rect 29779 4777 29788 4811
rect 29736 4768 29788 4777
rect 5540 4700 5592 4752
rect 3884 4564 3936 4616
rect 4988 4607 5040 4616
rect 4988 4573 4997 4607
rect 4997 4573 5031 4607
rect 5031 4573 5040 4607
rect 4988 4564 5040 4573
rect 5080 4607 5132 4616
rect 5080 4573 5089 4607
rect 5089 4573 5123 4607
rect 5123 4573 5132 4607
rect 5080 4564 5132 4573
rect 5264 4564 5316 4616
rect 2872 4496 2924 4548
rect 4068 4496 4120 4548
rect 4620 4496 4672 4548
rect 7656 4632 7708 4684
rect 5816 4607 5868 4616
rect 5816 4573 5825 4607
rect 5825 4573 5859 4607
rect 5859 4573 5868 4607
rect 5816 4564 5868 4573
rect 5908 4564 5960 4616
rect 6552 4564 6604 4616
rect 7288 4564 7340 4616
rect 9496 4700 9548 4752
rect 9772 4743 9824 4752
rect 9772 4709 9781 4743
rect 9781 4709 9815 4743
rect 9815 4709 9824 4743
rect 9772 4700 9824 4709
rect 8944 4675 8996 4684
rect 8944 4641 8953 4675
rect 8953 4641 8987 4675
rect 8987 4641 8996 4675
rect 8944 4632 8996 4641
rect 8208 4607 8260 4616
rect 8208 4573 8217 4607
rect 8217 4573 8251 4607
rect 8251 4573 8260 4607
rect 8208 4564 8260 4573
rect 9404 4428 9456 4480
rect 10324 4632 10376 4684
rect 13912 4632 13964 4684
rect 12440 4607 12492 4616
rect 12440 4573 12449 4607
rect 12449 4573 12483 4607
rect 12483 4573 12492 4607
rect 12440 4564 12492 4573
rect 12624 4564 12676 4616
rect 12900 4607 12952 4616
rect 12900 4573 12909 4607
rect 12909 4573 12943 4607
rect 12943 4573 12952 4607
rect 12900 4564 12952 4573
rect 13084 4607 13136 4616
rect 13084 4573 13093 4607
rect 13093 4573 13127 4607
rect 13127 4573 13136 4607
rect 13084 4564 13136 4573
rect 14096 4607 14148 4616
rect 14096 4573 14105 4607
rect 14105 4573 14139 4607
rect 14139 4573 14148 4607
rect 14096 4564 14148 4573
rect 14740 4632 14792 4684
rect 17132 4632 17184 4684
rect 19340 4632 19392 4684
rect 20536 4700 20588 4752
rect 21824 4700 21876 4752
rect 23572 4700 23624 4752
rect 25872 4700 25924 4752
rect 30564 4768 30616 4820
rect 31392 4811 31444 4820
rect 31392 4777 31401 4811
rect 31401 4777 31435 4811
rect 31435 4777 31444 4811
rect 31392 4768 31444 4777
rect 31760 4768 31812 4820
rect 32220 4811 32272 4820
rect 32220 4777 32229 4811
rect 32229 4777 32263 4811
rect 32263 4777 32272 4811
rect 32220 4768 32272 4777
rect 33048 4811 33100 4820
rect 33048 4777 33057 4811
rect 33057 4777 33091 4811
rect 33091 4777 33100 4811
rect 33048 4768 33100 4777
rect 33140 4768 33192 4820
rect 23664 4632 23716 4684
rect 14464 4607 14516 4616
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 14648 4564 14700 4616
rect 17592 4564 17644 4616
rect 18420 4607 18472 4616
rect 18420 4573 18429 4607
rect 18429 4573 18463 4607
rect 18463 4573 18472 4607
rect 18420 4564 18472 4573
rect 19984 4564 20036 4616
rect 14280 4539 14332 4548
rect 10600 4428 10652 4480
rect 14280 4505 14289 4539
rect 14289 4505 14323 4539
rect 14323 4505 14332 4539
rect 14280 4496 14332 4505
rect 13268 4471 13320 4480
rect 13268 4437 13277 4471
rect 13277 4437 13311 4471
rect 13311 4437 13320 4471
rect 13268 4428 13320 4437
rect 13636 4428 13688 4480
rect 16580 4496 16632 4548
rect 20536 4564 20588 4616
rect 22376 4564 22428 4616
rect 23204 4607 23256 4616
rect 23204 4573 23213 4607
rect 23213 4573 23247 4607
rect 23247 4573 23256 4607
rect 23204 4564 23256 4573
rect 27620 4632 27672 4684
rect 25136 4607 25188 4616
rect 25136 4573 25145 4607
rect 25145 4573 25179 4607
rect 25179 4573 25188 4607
rect 25136 4564 25188 4573
rect 26056 4564 26108 4616
rect 26792 4564 26844 4616
rect 27712 4564 27764 4616
rect 28724 4607 28776 4616
rect 28724 4573 28733 4607
rect 28733 4573 28767 4607
rect 28767 4573 28776 4607
rect 28724 4564 28776 4573
rect 29000 4607 29052 4616
rect 29000 4573 29009 4607
rect 29009 4573 29043 4607
rect 29043 4573 29052 4607
rect 29000 4564 29052 4573
rect 24768 4496 24820 4548
rect 34428 4700 34480 4752
rect 35716 4768 35768 4820
rect 34612 4700 34664 4752
rect 35348 4700 35400 4752
rect 35808 4700 35860 4752
rect 33968 4564 34020 4616
rect 35716 4607 35768 4616
rect 29460 4496 29512 4548
rect 31208 4539 31260 4548
rect 31208 4505 31217 4539
rect 31217 4505 31251 4539
rect 31251 4505 31260 4539
rect 31208 4496 31260 4505
rect 16488 4471 16540 4480
rect 16488 4437 16497 4471
rect 16497 4437 16531 4471
rect 16531 4437 16540 4471
rect 16488 4428 16540 4437
rect 18144 4428 18196 4480
rect 20628 4428 20680 4480
rect 23480 4428 23532 4480
rect 27620 4471 27672 4480
rect 27620 4437 27629 4471
rect 27629 4437 27663 4471
rect 27663 4437 27672 4471
rect 27620 4428 27672 4437
rect 28356 4428 28408 4480
rect 28448 4428 28500 4480
rect 28816 4428 28868 4480
rect 29092 4428 29144 4480
rect 30380 4471 30432 4480
rect 30380 4437 30389 4471
rect 30389 4437 30423 4471
rect 30423 4437 30432 4471
rect 30380 4428 30432 4437
rect 31668 4496 31720 4548
rect 33508 4496 33560 4548
rect 34336 4496 34388 4548
rect 32220 4471 32272 4480
rect 32220 4437 32245 4471
rect 32245 4437 32272 4471
rect 32220 4428 32272 4437
rect 32956 4428 33008 4480
rect 33232 4428 33284 4480
rect 34888 4471 34940 4480
rect 35716 4573 35725 4607
rect 35725 4573 35759 4607
rect 35759 4573 35768 4607
rect 35716 4564 35768 4573
rect 37556 4564 37608 4616
rect 34888 4437 34913 4471
rect 34913 4437 34940 4471
rect 34888 4428 34940 4437
rect 36176 4471 36228 4480
rect 36176 4437 36185 4471
rect 36185 4437 36219 4471
rect 36219 4437 36228 4471
rect 36176 4428 36228 4437
rect 36452 4428 36504 4480
rect 39028 4428 39080 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 2044 4224 2096 4276
rect 3240 4267 3292 4276
rect 3240 4233 3249 4267
rect 3249 4233 3283 4267
rect 3283 4233 3292 4267
rect 3240 4224 3292 4233
rect 3424 4224 3476 4276
rect 12256 4224 12308 4276
rect 14096 4224 14148 4276
rect 15568 4224 15620 4276
rect 18328 4224 18380 4276
rect 3700 4156 3752 4208
rect 3792 4156 3844 4208
rect 3240 4088 3292 4140
rect 5908 4156 5960 4208
rect 4620 4088 4672 4140
rect 4988 4088 5040 4140
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 6644 4131 6696 4140
rect 6644 4097 6653 4131
rect 6653 4097 6687 4131
rect 6687 4097 6696 4131
rect 6920 4131 6972 4140
rect 6644 4088 6696 4097
rect 6920 4097 6929 4131
rect 6929 4097 6963 4131
rect 6963 4097 6972 4131
rect 6920 4088 6972 4097
rect 10324 4156 10376 4208
rect 11244 4156 11296 4208
rect 3792 4020 3844 4072
rect 7196 4020 7248 4072
rect 5080 3952 5132 4004
rect 6828 3995 6880 4004
rect 6828 3961 6837 3995
rect 6837 3961 6871 3995
rect 6871 3961 6880 3995
rect 6828 3952 6880 3961
rect 5724 3884 5776 3936
rect 6644 3884 6696 3936
rect 8760 3927 8812 3936
rect 8760 3893 8769 3927
rect 8769 3893 8803 3927
rect 8803 3893 8812 3927
rect 8760 3884 8812 3893
rect 9496 4131 9548 4140
rect 9496 4097 9530 4131
rect 9530 4097 9548 4131
rect 9496 4088 9548 4097
rect 11428 4088 11480 4140
rect 10416 4020 10468 4072
rect 13544 4088 13596 4140
rect 14740 4156 14792 4208
rect 19432 4199 19484 4208
rect 19432 4165 19441 4199
rect 19441 4165 19475 4199
rect 19475 4165 19484 4199
rect 19432 4156 19484 4165
rect 19984 4224 20036 4276
rect 13912 4131 13964 4140
rect 13912 4097 13946 4131
rect 13946 4097 13964 4131
rect 13912 4088 13964 4097
rect 14280 4088 14332 4140
rect 14832 4088 14884 4140
rect 15292 4088 15344 4140
rect 15476 4131 15528 4140
rect 15476 4097 15485 4131
rect 15485 4097 15519 4131
rect 15519 4097 15528 4131
rect 15476 4088 15528 4097
rect 15752 4131 15804 4140
rect 15752 4097 15761 4131
rect 15761 4097 15795 4131
rect 15795 4097 15804 4131
rect 15752 4088 15804 4097
rect 11060 3952 11112 4004
rect 11612 3952 11664 4004
rect 9864 3884 9916 3936
rect 9956 3884 10008 3936
rect 13636 3952 13688 4004
rect 15660 3952 15712 4004
rect 15936 4088 15988 4140
rect 17040 4063 17092 4072
rect 13820 3884 13872 3936
rect 14740 3884 14792 3936
rect 17040 4029 17049 4063
rect 17049 4029 17083 4063
rect 17083 4029 17092 4063
rect 17040 4020 17092 4029
rect 19616 4131 19668 4140
rect 19616 4097 19625 4131
rect 19625 4097 19659 4131
rect 19659 4097 19668 4131
rect 19616 4088 19668 4097
rect 20352 4156 20404 4208
rect 20812 4156 20864 4208
rect 20536 4088 20588 4140
rect 20260 4063 20312 4072
rect 20260 4029 20269 4063
rect 20269 4029 20303 4063
rect 20303 4029 20312 4063
rect 20260 4020 20312 4029
rect 20352 4020 20404 4072
rect 22284 4156 22336 4208
rect 22100 4131 22152 4140
rect 22100 4097 22134 4131
rect 22134 4097 22152 4131
rect 22468 4224 22520 4276
rect 22652 4224 22704 4276
rect 33508 4267 33560 4276
rect 33508 4233 33517 4267
rect 33517 4233 33551 4267
rect 33551 4233 33560 4267
rect 33508 4224 33560 4233
rect 34796 4224 34848 4276
rect 35808 4267 35860 4276
rect 35808 4233 35817 4267
rect 35817 4233 35851 4267
rect 35851 4233 35860 4267
rect 35808 4224 35860 4233
rect 22100 4088 22152 4097
rect 24400 4020 24452 4072
rect 25688 4156 25740 4208
rect 25320 4088 25372 4140
rect 25780 4088 25832 4140
rect 26056 4131 26108 4140
rect 26056 4097 26065 4131
rect 26065 4097 26099 4131
rect 26099 4097 26108 4131
rect 26056 4088 26108 4097
rect 26148 4131 26200 4140
rect 26148 4097 26157 4131
rect 26157 4097 26191 4131
rect 26191 4097 26200 4131
rect 26332 4131 26384 4140
rect 26148 4088 26200 4097
rect 26332 4097 26341 4131
rect 26341 4097 26375 4131
rect 26375 4097 26384 4131
rect 26332 4088 26384 4097
rect 24952 4020 25004 4072
rect 16120 3884 16172 3936
rect 18052 3884 18104 3936
rect 19524 3952 19576 4004
rect 20168 3884 20220 3936
rect 21272 3952 21324 4004
rect 20812 3884 20864 3936
rect 22100 3884 22152 3936
rect 27620 4088 27672 4140
rect 30012 4156 30064 4208
rect 29460 4088 29512 4140
rect 29736 4088 29788 4140
rect 30288 4131 30340 4140
rect 30288 4097 30297 4131
rect 30297 4097 30331 4131
rect 30331 4097 30340 4131
rect 30288 4088 30340 4097
rect 30472 4131 30524 4140
rect 30472 4097 30481 4131
rect 30481 4097 30515 4131
rect 30515 4097 30524 4131
rect 30472 4088 30524 4097
rect 36084 4156 36136 4208
rect 36360 4156 36412 4208
rect 31392 4131 31444 4140
rect 26976 4063 27028 4072
rect 26976 4029 26985 4063
rect 26985 4029 27019 4063
rect 27019 4029 27028 4063
rect 26976 4020 27028 4029
rect 28080 4020 28132 4072
rect 28724 4020 28776 4072
rect 29000 4020 29052 4072
rect 30196 4020 30248 4072
rect 31392 4097 31401 4131
rect 31401 4097 31435 4131
rect 31435 4097 31444 4131
rect 31392 4088 31444 4097
rect 32680 4088 32732 4140
rect 37832 4131 37884 4140
rect 34428 4063 34480 4072
rect 23204 3927 23256 3936
rect 23204 3893 23213 3927
rect 23213 3893 23247 3927
rect 23247 3893 23256 3927
rect 23204 3884 23256 3893
rect 23296 3884 23348 3936
rect 25872 3884 25924 3936
rect 30656 3952 30708 4004
rect 34428 4029 34437 4063
rect 34437 4029 34471 4063
rect 34471 4029 34480 4063
rect 34428 4020 34480 4029
rect 37832 4097 37841 4131
rect 37841 4097 37875 4131
rect 37875 4097 37884 4131
rect 37832 4088 37884 4097
rect 37924 4020 37976 4072
rect 28356 3927 28408 3936
rect 28356 3893 28365 3927
rect 28365 3893 28399 3927
rect 28399 3893 28408 3927
rect 28356 3884 28408 3893
rect 30104 3927 30156 3936
rect 30104 3893 30113 3927
rect 30113 3893 30147 3927
rect 30147 3893 30156 3927
rect 30104 3884 30156 3893
rect 31024 3927 31076 3936
rect 31024 3893 31033 3927
rect 31033 3893 31067 3927
rect 31067 3893 31076 3927
rect 31024 3884 31076 3893
rect 32128 3884 32180 3936
rect 37740 3952 37792 4004
rect 36452 3927 36504 3936
rect 36452 3893 36461 3927
rect 36461 3893 36495 3927
rect 36495 3893 36504 3927
rect 36452 3884 36504 3893
rect 38292 3884 38344 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 3700 3680 3752 3732
rect 7104 3723 7156 3732
rect 1952 3519 2004 3528
rect 1952 3485 1961 3519
rect 1961 3485 1995 3519
rect 1995 3485 2004 3519
rect 1952 3476 2004 3485
rect 2964 3408 3016 3460
rect 5264 3612 5316 3664
rect 7104 3689 7113 3723
rect 7113 3689 7147 3723
rect 7147 3689 7156 3723
rect 7104 3680 7156 3689
rect 7196 3680 7248 3732
rect 8116 3680 8168 3732
rect 9496 3680 9548 3732
rect 9864 3680 9916 3732
rect 7380 3612 7432 3664
rect 9956 3612 10008 3664
rect 5080 3476 5132 3528
rect 4344 3408 4396 3460
rect 3976 3340 4028 3392
rect 4068 3340 4120 3392
rect 4896 3340 4948 3392
rect 7932 3544 7984 3596
rect 9036 3544 9088 3596
rect 10600 3680 10652 3732
rect 11336 3680 11388 3732
rect 11796 3612 11848 3664
rect 5908 3476 5960 3528
rect 7288 3519 7340 3528
rect 7288 3485 7297 3519
rect 7297 3485 7331 3519
rect 7331 3485 7340 3519
rect 7288 3476 7340 3485
rect 7380 3519 7432 3528
rect 7380 3485 7389 3519
rect 7389 3485 7423 3519
rect 7423 3485 7432 3519
rect 7380 3476 7432 3485
rect 5632 3408 5684 3460
rect 5724 3408 5776 3460
rect 6460 3408 6512 3460
rect 6644 3408 6696 3460
rect 8576 3476 8628 3528
rect 9404 3519 9456 3528
rect 9404 3485 9413 3519
rect 9413 3485 9447 3519
rect 9447 3485 9456 3519
rect 9404 3476 9456 3485
rect 10232 3476 10284 3528
rect 11336 3476 11388 3528
rect 11704 3519 11756 3528
rect 11704 3485 11713 3519
rect 11713 3485 11747 3519
rect 11747 3485 11756 3519
rect 11704 3476 11756 3485
rect 12164 3680 12216 3732
rect 13084 3680 13136 3732
rect 13636 3680 13688 3732
rect 15016 3680 15068 3732
rect 15476 3680 15528 3732
rect 17960 3680 18012 3732
rect 19616 3680 19668 3732
rect 18880 3612 18932 3664
rect 20628 3612 20680 3664
rect 21272 3680 21324 3732
rect 23204 3680 23256 3732
rect 25136 3680 25188 3732
rect 25504 3680 25556 3732
rect 27344 3680 27396 3732
rect 27528 3680 27580 3732
rect 30012 3680 30064 3732
rect 30472 3680 30524 3732
rect 10048 3408 10100 3460
rect 10600 3451 10652 3460
rect 10600 3417 10609 3451
rect 10609 3417 10643 3451
rect 10643 3417 10652 3451
rect 10600 3408 10652 3417
rect 11980 3408 12032 3460
rect 12164 3340 12216 3392
rect 12900 3340 12952 3392
rect 13084 3476 13136 3528
rect 14096 3544 14148 3596
rect 14464 3544 14516 3596
rect 14740 3544 14792 3596
rect 17040 3544 17092 3596
rect 20260 3544 20312 3596
rect 14280 3476 14332 3528
rect 16028 3476 16080 3528
rect 19432 3519 19484 3528
rect 13544 3408 13596 3460
rect 13728 3408 13780 3460
rect 15200 3408 15252 3460
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 20168 3476 20220 3528
rect 22192 3612 22244 3664
rect 21916 3544 21968 3596
rect 22284 3544 22336 3596
rect 21088 3476 21140 3528
rect 21732 3476 21784 3528
rect 22008 3476 22060 3528
rect 24400 3587 24452 3596
rect 24400 3553 24409 3587
rect 24409 3553 24443 3587
rect 24443 3553 24452 3587
rect 24400 3544 24452 3553
rect 25044 3544 25096 3596
rect 26056 3612 26108 3664
rect 32036 3680 32088 3732
rect 34520 3680 34572 3732
rect 36452 3680 36504 3732
rect 36912 3723 36964 3732
rect 36912 3689 36921 3723
rect 36921 3689 36955 3723
rect 36955 3689 36964 3723
rect 36912 3680 36964 3689
rect 32312 3612 32364 3664
rect 34612 3612 34664 3664
rect 26884 3544 26936 3596
rect 26976 3544 27028 3596
rect 24584 3519 24636 3528
rect 19800 3408 19852 3460
rect 20628 3408 20680 3460
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 26240 3476 26292 3528
rect 26424 3519 26476 3528
rect 26424 3485 26433 3519
rect 26433 3485 26467 3519
rect 26467 3485 26476 3519
rect 26424 3476 26476 3485
rect 30748 3544 30800 3596
rect 33416 3544 33468 3596
rect 34428 3544 34480 3596
rect 29736 3519 29788 3528
rect 29736 3485 29745 3519
rect 29745 3485 29779 3519
rect 29779 3485 29788 3519
rect 29736 3476 29788 3485
rect 32128 3476 32180 3528
rect 33508 3476 33560 3528
rect 35440 3476 35492 3528
rect 37464 3476 37516 3528
rect 22744 3451 22796 3460
rect 22744 3417 22778 3451
rect 22778 3417 22796 3451
rect 22744 3408 22796 3417
rect 23112 3408 23164 3460
rect 13820 3340 13872 3392
rect 15936 3340 15988 3392
rect 18604 3340 18656 3392
rect 19432 3340 19484 3392
rect 20904 3340 20956 3392
rect 21272 3340 21324 3392
rect 23664 3340 23716 3392
rect 23848 3383 23900 3392
rect 23848 3349 23857 3383
rect 23857 3349 23891 3383
rect 23891 3349 23900 3383
rect 23848 3340 23900 3349
rect 26332 3340 26384 3392
rect 28448 3408 28500 3460
rect 30104 3408 30156 3460
rect 30472 3408 30524 3460
rect 32404 3451 32456 3460
rect 32404 3417 32413 3451
rect 32413 3417 32447 3451
rect 32447 3417 32456 3451
rect 32404 3408 32456 3417
rect 35624 3408 35676 3460
rect 27528 3340 27580 3392
rect 28816 3340 28868 3392
rect 29368 3340 29420 3392
rect 31300 3340 31352 3392
rect 32220 3340 32272 3392
rect 33968 3340 34020 3392
rect 34336 3340 34388 3392
rect 35348 3340 35400 3392
rect 36360 3340 36412 3392
rect 37556 3340 37608 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2964 3136 3016 3188
rect 4252 3136 4304 3188
rect 4620 3136 4672 3188
rect 5632 3179 5684 3188
rect 5632 3145 5641 3179
rect 5641 3145 5675 3179
rect 5675 3145 5684 3179
rect 5632 3136 5684 3145
rect 8024 3179 8076 3188
rect 8024 3145 8033 3179
rect 8033 3145 8067 3179
rect 8067 3145 8076 3179
rect 8024 3136 8076 3145
rect 8116 3136 8168 3188
rect 3056 3000 3108 3052
rect 3792 3000 3844 3052
rect 4160 3000 4212 3052
rect 4896 3000 4948 3052
rect 5724 3000 5776 3052
rect 6000 3000 6052 3052
rect 9956 3068 10008 3120
rect 12900 3136 12952 3188
rect 15752 3136 15804 3188
rect 16580 3136 16632 3188
rect 18420 3136 18472 3188
rect 20536 3136 20588 3188
rect 20720 3179 20772 3188
rect 20720 3145 20729 3179
rect 20729 3145 20763 3179
rect 20763 3145 20772 3179
rect 20720 3136 20772 3145
rect 21732 3136 21784 3188
rect 23848 3136 23900 3188
rect 24492 3179 24544 3188
rect 24492 3145 24501 3179
rect 24501 3145 24535 3179
rect 24535 3145 24544 3179
rect 24492 3136 24544 3145
rect 25596 3136 25648 3188
rect 27804 3179 27856 3188
rect 27804 3145 27813 3179
rect 27813 3145 27847 3179
rect 27847 3145 27856 3179
rect 27804 3136 27856 3145
rect 28080 3136 28132 3188
rect 28908 3136 28960 3188
rect 30748 3136 30800 3188
rect 31392 3136 31444 3188
rect 10784 3068 10836 3120
rect 14740 3068 14792 3120
rect 15292 3068 15344 3120
rect 15568 3068 15620 3120
rect 18236 3111 18288 3120
rect 18236 3077 18245 3111
rect 18245 3077 18279 3111
rect 18279 3077 18288 3111
rect 18236 3068 18288 3077
rect 2964 2932 3016 2984
rect 5908 2932 5960 2984
rect 7380 3000 7432 3052
rect 6644 2864 6696 2916
rect 3424 2796 3476 2848
rect 4804 2796 4856 2848
rect 6920 2796 6972 2848
rect 7012 2796 7064 2848
rect 10048 3000 10100 3052
rect 8852 2975 8904 2984
rect 8852 2941 8861 2975
rect 8861 2941 8895 2975
rect 8895 2941 8904 2975
rect 8852 2932 8904 2941
rect 9036 2932 9088 2984
rect 10232 3000 10284 3052
rect 10508 3043 10560 3052
rect 10508 3009 10517 3043
rect 10517 3009 10551 3043
rect 10551 3009 10560 3043
rect 10508 3000 10560 3009
rect 11336 3000 11388 3052
rect 11428 3000 11480 3052
rect 11796 3043 11848 3052
rect 11796 3009 11830 3043
rect 11830 3009 11848 3043
rect 11796 3000 11848 3009
rect 12992 3000 13044 3052
rect 13544 3043 13596 3052
rect 13544 3009 13553 3043
rect 13553 3009 13587 3043
rect 13587 3009 13596 3043
rect 13544 3000 13596 3009
rect 11060 2932 11112 2984
rect 12716 2932 12768 2984
rect 14096 3000 14148 3052
rect 16120 3043 16172 3052
rect 14648 2975 14700 2984
rect 14648 2941 14657 2975
rect 14657 2941 14691 2975
rect 14691 2941 14700 2975
rect 14648 2932 14700 2941
rect 16120 3009 16129 3043
rect 16129 3009 16163 3043
rect 16163 3009 16172 3043
rect 16120 3000 16172 3009
rect 17960 3043 18012 3052
rect 17960 3009 17969 3043
rect 17969 3009 18003 3043
rect 18003 3009 18012 3043
rect 17960 3000 18012 3009
rect 18328 3043 18380 3052
rect 15752 2932 15804 2984
rect 16304 2932 16356 2984
rect 16948 2975 17000 2984
rect 16948 2941 16957 2975
rect 16957 2941 16991 2975
rect 16991 2941 17000 2975
rect 18328 3009 18337 3043
rect 18337 3009 18371 3043
rect 18371 3009 18380 3043
rect 18328 3000 18380 3009
rect 20628 3068 20680 3120
rect 20076 3000 20128 3052
rect 20260 3000 20312 3052
rect 20996 3000 21048 3052
rect 21732 3000 21784 3052
rect 16948 2932 17000 2941
rect 21916 2932 21968 2984
rect 22652 3068 22704 3120
rect 23480 3068 23532 3120
rect 23664 3068 23716 3120
rect 22192 3043 22244 3052
rect 22192 3009 22201 3043
rect 22201 3009 22235 3043
rect 22235 3009 22244 3043
rect 22192 3000 22244 3009
rect 22928 3000 22980 3052
rect 25964 3000 26016 3052
rect 27988 3068 28040 3120
rect 28540 3068 28592 3120
rect 28816 3068 28868 3120
rect 31024 3068 31076 3120
rect 33876 3136 33928 3188
rect 34152 3179 34204 3188
rect 34152 3145 34161 3179
rect 34161 3145 34195 3179
rect 34195 3145 34204 3179
rect 34152 3136 34204 3145
rect 35348 3111 35400 3120
rect 35348 3077 35357 3111
rect 35357 3077 35391 3111
rect 35391 3077 35400 3111
rect 35348 3068 35400 3077
rect 26884 3000 26936 3052
rect 29644 3000 29696 3052
rect 29736 3000 29788 3052
rect 30840 3000 30892 3052
rect 10232 2864 10284 2916
rect 10600 2864 10652 2916
rect 8300 2796 8352 2848
rect 9128 2796 9180 2848
rect 9312 2796 9364 2848
rect 9496 2796 9548 2848
rect 10140 2796 10192 2848
rect 10784 2796 10836 2848
rect 13728 2864 13780 2916
rect 21272 2864 21324 2916
rect 12992 2796 13044 2848
rect 13912 2839 13964 2848
rect 13912 2805 13921 2839
rect 13921 2805 13955 2839
rect 13955 2805 13964 2839
rect 13912 2796 13964 2805
rect 14556 2796 14608 2848
rect 16672 2796 16724 2848
rect 18052 2796 18104 2848
rect 21088 2796 21140 2848
rect 21180 2796 21232 2848
rect 22100 2796 22152 2848
rect 22284 2932 22336 2984
rect 24400 2932 24452 2984
rect 25136 2932 25188 2984
rect 22376 2907 22428 2916
rect 22376 2873 22385 2907
rect 22385 2873 22419 2907
rect 22419 2873 22428 2907
rect 22376 2864 22428 2873
rect 22928 2864 22980 2916
rect 23296 2864 23348 2916
rect 23848 2864 23900 2916
rect 29184 2932 29236 2984
rect 31300 3000 31352 3052
rect 31760 3000 31812 3052
rect 32864 3043 32916 3052
rect 32312 2932 32364 2984
rect 32864 3009 32873 3043
rect 32873 3009 32907 3043
rect 32907 3009 32916 3043
rect 32864 3000 32916 3009
rect 33324 2932 33376 2984
rect 25504 2864 25556 2916
rect 26056 2864 26108 2916
rect 28080 2864 28132 2916
rect 28540 2864 28592 2916
rect 23112 2796 23164 2848
rect 24308 2796 24360 2848
rect 24768 2796 24820 2848
rect 28632 2839 28684 2848
rect 28632 2805 28641 2839
rect 28641 2805 28675 2839
rect 28675 2805 28684 2839
rect 28632 2796 28684 2805
rect 28724 2796 28776 2848
rect 28908 2796 28960 2848
rect 29460 2839 29512 2848
rect 29460 2805 29469 2839
rect 29469 2805 29503 2839
rect 29503 2805 29512 2839
rect 29460 2796 29512 2805
rect 30748 2796 30800 2848
rect 31576 2796 31628 2848
rect 33784 2864 33836 2916
rect 36268 3136 36320 3188
rect 37096 3136 37148 3188
rect 35808 3068 35860 3120
rect 36360 3111 36412 3120
rect 36360 3077 36385 3111
rect 36385 3077 36412 3111
rect 36360 3068 36412 3077
rect 37372 3000 37424 3052
rect 36176 2864 36228 2916
rect 32312 2839 32364 2848
rect 32312 2805 32321 2839
rect 32321 2805 32355 2839
rect 32355 2805 32364 2839
rect 32312 2796 32364 2805
rect 36452 2796 36504 2848
rect 36820 2796 36872 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 572 2388 624 2440
rect 3240 2592 3292 2644
rect 3332 2592 3384 2644
rect 5356 2592 5408 2644
rect 6460 2592 6512 2644
rect 7380 2635 7432 2644
rect 7380 2601 7389 2635
rect 7389 2601 7423 2635
rect 7423 2601 7432 2635
rect 7380 2592 7432 2601
rect 8116 2592 8168 2644
rect 9220 2592 9272 2644
rect 10324 2635 10376 2644
rect 10324 2601 10333 2635
rect 10333 2601 10367 2635
rect 10367 2601 10376 2635
rect 10324 2592 10376 2601
rect 11244 2592 11296 2644
rect 11796 2592 11848 2644
rect 15844 2592 15896 2644
rect 16580 2592 16632 2644
rect 21548 2592 21600 2644
rect 23020 2592 23072 2644
rect 24952 2592 25004 2644
rect 27896 2592 27948 2644
rect 28632 2592 28684 2644
rect 28908 2592 28960 2644
rect 30748 2592 30800 2644
rect 6092 2524 6144 2576
rect 6920 2524 6972 2576
rect 8024 2524 8076 2576
rect 3884 2456 3936 2508
rect 3976 2456 4028 2508
rect 7380 2456 7432 2508
rect 3608 2388 3660 2440
rect 4620 2388 4672 2440
rect 4988 2431 5040 2440
rect 4988 2397 4997 2431
rect 4997 2397 5031 2431
rect 5031 2397 5040 2431
rect 4988 2388 5040 2397
rect 7472 2388 7524 2440
rect 8116 2431 8168 2440
rect 8116 2397 8125 2431
rect 8125 2397 8159 2431
rect 8159 2397 8168 2431
rect 8116 2388 8168 2397
rect 8208 2431 8260 2440
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 9220 2456 9272 2508
rect 8208 2388 8260 2397
rect 9036 2388 9088 2440
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 7840 2320 7892 2372
rect 9404 2388 9456 2440
rect 10140 2431 10192 2440
rect 10140 2397 10149 2431
rect 10149 2397 10183 2431
rect 10183 2397 10192 2431
rect 10140 2388 10192 2397
rect 13268 2524 13320 2576
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 16304 2524 16356 2576
rect 13912 2388 13964 2440
rect 3148 2252 3200 2304
rect 4712 2252 4764 2304
rect 7288 2252 7340 2304
rect 7380 2252 7432 2304
rect 9312 2252 9364 2304
rect 12348 2252 12400 2304
rect 14832 2456 14884 2508
rect 17408 2524 17460 2576
rect 24860 2524 24912 2576
rect 25596 2524 25648 2576
rect 27804 2524 27856 2576
rect 32312 2524 32364 2576
rect 34612 2524 34664 2576
rect 36084 2524 36136 2576
rect 17592 2456 17644 2508
rect 15752 2431 15804 2440
rect 15752 2397 15761 2431
rect 15761 2397 15795 2431
rect 15795 2397 15804 2431
rect 15752 2388 15804 2397
rect 16764 2431 16816 2440
rect 16764 2397 16773 2431
rect 16773 2397 16807 2431
rect 16807 2397 16816 2431
rect 16764 2388 16816 2397
rect 16948 2431 17000 2440
rect 16948 2397 16957 2431
rect 16957 2397 16991 2431
rect 16991 2397 17000 2431
rect 16948 2388 17000 2397
rect 17132 2388 17184 2440
rect 18328 2456 18380 2508
rect 17868 2431 17920 2440
rect 17868 2397 17877 2431
rect 17877 2397 17911 2431
rect 17911 2397 17920 2431
rect 17868 2388 17920 2397
rect 15660 2363 15712 2372
rect 15660 2329 15669 2363
rect 15669 2329 15703 2363
rect 15703 2329 15712 2363
rect 15660 2320 15712 2329
rect 16028 2320 16080 2372
rect 17040 2363 17092 2372
rect 16488 2252 16540 2304
rect 17040 2329 17049 2363
rect 17049 2329 17083 2363
rect 17083 2329 17092 2363
rect 17040 2320 17092 2329
rect 17592 2320 17644 2372
rect 18052 2388 18104 2440
rect 19340 2456 19392 2508
rect 22376 2499 22428 2508
rect 22376 2465 22385 2499
rect 22385 2465 22419 2499
rect 22419 2465 22428 2499
rect 22376 2456 22428 2465
rect 24216 2456 24268 2508
rect 18604 2388 18656 2440
rect 20812 2388 20864 2440
rect 21088 2431 21140 2440
rect 21088 2397 21097 2431
rect 21097 2397 21131 2431
rect 21131 2397 21140 2431
rect 21088 2388 21140 2397
rect 22560 2431 22612 2440
rect 22560 2397 22569 2431
rect 22569 2397 22603 2431
rect 22603 2397 22612 2431
rect 22560 2388 22612 2397
rect 24032 2388 24084 2440
rect 25228 2388 25280 2440
rect 25504 2431 25556 2440
rect 25504 2397 25513 2431
rect 25513 2397 25547 2431
rect 25547 2397 25556 2431
rect 25504 2388 25556 2397
rect 29276 2456 29328 2508
rect 29920 2456 29972 2508
rect 26240 2388 26292 2440
rect 26516 2388 26568 2440
rect 24308 2320 24360 2372
rect 28080 2388 28132 2440
rect 29552 2431 29604 2440
rect 28356 2363 28408 2372
rect 28356 2329 28365 2363
rect 28365 2329 28399 2363
rect 28399 2329 28408 2363
rect 28356 2320 28408 2329
rect 29552 2397 29561 2431
rect 29561 2397 29595 2431
rect 29595 2397 29604 2431
rect 29552 2388 29604 2397
rect 30380 2388 30432 2440
rect 35532 2456 35584 2508
rect 32036 2388 32088 2440
rect 33232 2388 33284 2440
rect 33416 2388 33468 2440
rect 34704 2431 34756 2440
rect 34704 2397 34713 2431
rect 34713 2397 34747 2431
rect 34747 2397 34756 2431
rect 34704 2388 34756 2397
rect 35900 2388 35952 2440
rect 37280 2431 37332 2440
rect 37280 2397 37289 2431
rect 37289 2397 37323 2431
rect 37323 2397 37332 2431
rect 37280 2388 37332 2397
rect 24124 2252 24176 2304
rect 29828 2320 29880 2372
rect 30104 2320 30156 2372
rect 28816 2252 28868 2304
rect 31760 2252 31812 2304
rect 35348 2320 35400 2372
rect 33140 2252 33192 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 3240 2048 3292 2100
rect 8392 2048 8444 2100
rect 8852 2048 8904 2100
rect 12348 2048 12400 2100
rect 7472 1980 7524 2032
rect 14004 1980 14056 2032
rect 1952 1912 2004 1964
rect 11336 1912 11388 1964
rect 1584 1844 1636 1896
rect 4988 1844 5040 1896
rect 11152 1844 11204 1896
rect 3056 1776 3108 1828
rect 17040 1776 17092 1828
rect 18972 1708 19024 1760
rect 2780 1640 2832 1692
rect 13268 1640 13320 1692
rect 1768 1572 1820 1624
rect 4988 1572 5040 1624
rect 5172 1572 5224 1624
rect 15660 1572 15712 1624
rect 3792 1368 3844 1420
rect 8024 1368 8076 1420
rect 27068 1368 27120 1420
rect 28816 1368 28868 1420
<< metal2 >>
rect 3974 49314 4030 50000
rect 11978 49314 12034 50000
rect 19982 49314 20038 50000
rect 27986 49314 28042 50000
rect 35990 49314 36046 50000
rect 3974 49286 4108 49314
rect 3974 49200 4030 49286
rect 4080 47138 4108 49286
rect 11978 49286 12296 49314
rect 11978 49200 12034 49286
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 12268 47258 12296 49286
rect 19982 49286 20300 49314
rect 19982 49200 20038 49286
rect 20272 47258 20300 49286
rect 27986 49286 28304 49314
rect 27986 49200 28042 49286
rect 28276 47258 28304 49286
rect 35990 49286 36216 49314
rect 35990 49200 36046 49286
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 12256 47252 12308 47258
rect 12256 47194 12308 47200
rect 20260 47252 20312 47258
rect 20260 47194 20312 47200
rect 28264 47252 28316 47258
rect 28264 47194 28316 47200
rect 4080 47110 4200 47138
rect 4172 47054 4200 47110
rect 36188 47054 36216 49286
rect 4160 47048 4212 47054
rect 4160 46990 4212 46996
rect 12440 47048 12492 47054
rect 12440 46990 12492 46996
rect 20352 47048 20404 47054
rect 20352 46990 20404 46996
rect 28080 47048 28132 47054
rect 28080 46990 28132 46996
rect 36176 47048 36228 47054
rect 36176 46990 36228 46996
rect 4620 46980 4672 46986
rect 4620 46922 4672 46928
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4632 29306 4660 46922
rect 12452 46714 12480 46990
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 12440 46708 12492 46714
rect 12440 46650 12492 46656
rect 12624 46572 12676 46578
rect 12624 46514 12676 46520
rect 15384 46572 15436 46578
rect 15384 46514 15436 46520
rect 12636 31754 12664 46514
rect 12544 31726 12664 31754
rect 4620 29300 4672 29306
rect 4620 29242 4672 29248
rect 12440 28960 12492 28966
rect 12440 28902 12492 28908
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 12452 28558 12480 28902
rect 9956 28552 10008 28558
rect 9956 28494 10008 28500
rect 11060 28552 11112 28558
rect 11060 28494 11112 28500
rect 11244 28552 11296 28558
rect 11244 28494 11296 28500
rect 12440 28552 12492 28558
rect 12440 28494 12492 28500
rect 8392 28484 8444 28490
rect 8392 28426 8444 28432
rect 9588 28484 9640 28490
rect 9588 28426 9640 28432
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 8404 27674 8432 28426
rect 8576 28076 8628 28082
rect 8576 28018 8628 28024
rect 8760 28076 8812 28082
rect 8760 28018 8812 28024
rect 8392 27668 8444 27674
rect 8392 27610 8444 27616
rect 8116 27532 8168 27538
rect 8116 27474 8168 27480
rect 8024 27464 8076 27470
rect 8024 27406 8076 27412
rect 8036 27130 8064 27406
rect 8024 27124 8076 27130
rect 8024 27066 8076 27072
rect 8024 26784 8076 26790
rect 8024 26726 8076 26732
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 8036 26586 8064 26726
rect 8024 26580 8076 26586
rect 8024 26522 8076 26528
rect 7748 26240 7800 26246
rect 7748 26182 7800 26188
rect 7760 25906 7788 26182
rect 8128 25906 8156 27474
rect 8392 26988 8444 26994
rect 8392 26930 8444 26936
rect 8300 26920 8352 26926
rect 8300 26862 8352 26868
rect 8312 26450 8340 26862
rect 8300 26444 8352 26450
rect 8300 26386 8352 26392
rect 8404 26330 8432 26930
rect 8588 26926 8616 28018
rect 8772 27334 8800 28018
rect 9128 27872 9180 27878
rect 9128 27814 9180 27820
rect 9140 27470 9168 27814
rect 8944 27464 8996 27470
rect 8944 27406 8996 27412
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 9220 27464 9272 27470
rect 9220 27406 9272 27412
rect 8760 27328 8812 27334
rect 8760 27270 8812 27276
rect 8772 26994 8800 27270
rect 8956 27062 8984 27406
rect 9232 27130 9260 27406
rect 9220 27124 9272 27130
rect 9220 27066 9272 27072
rect 8944 27056 8996 27062
rect 8944 26998 8996 27004
rect 8760 26988 8812 26994
rect 8760 26930 8812 26936
rect 8576 26920 8628 26926
rect 8576 26862 8628 26868
rect 8772 26586 8800 26930
rect 8944 26920 8996 26926
rect 8944 26862 8996 26868
rect 8852 26852 8904 26858
rect 8852 26794 8904 26800
rect 8760 26580 8812 26586
rect 8760 26522 8812 26528
rect 8668 26512 8720 26518
rect 8668 26454 8720 26460
rect 8312 26314 8432 26330
rect 8300 26308 8432 26314
rect 8352 26302 8432 26308
rect 8300 26250 8352 26256
rect 7748 25900 7800 25906
rect 7748 25842 7800 25848
rect 7932 25900 7984 25906
rect 7932 25842 7984 25848
rect 8116 25900 8168 25906
rect 8116 25842 8168 25848
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 7012 25288 7064 25294
rect 7012 25230 7064 25236
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 7024 23730 7052 25230
rect 7012 23724 7064 23730
rect 7012 23666 7064 23672
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 6932 22234 6960 22578
rect 6920 22228 6972 22234
rect 6920 22170 6972 22176
rect 7760 21554 7788 25842
rect 7944 24954 7972 25842
rect 8024 25832 8076 25838
rect 8024 25774 8076 25780
rect 8036 25498 8064 25774
rect 8024 25492 8076 25498
rect 8024 25434 8076 25440
rect 7932 24948 7984 24954
rect 7932 24890 7984 24896
rect 8128 23322 8156 25842
rect 8312 25242 8340 26250
rect 8392 25900 8444 25906
rect 8392 25842 8444 25848
rect 8404 25430 8432 25842
rect 8484 25696 8536 25702
rect 8484 25638 8536 25644
rect 8392 25424 8444 25430
rect 8392 25366 8444 25372
rect 8496 25294 8524 25638
rect 8680 25362 8708 26454
rect 8668 25356 8720 25362
rect 8668 25298 8720 25304
rect 8484 25288 8536 25294
rect 8312 25226 8432 25242
rect 8484 25230 8536 25236
rect 8312 25220 8444 25226
rect 8312 25214 8392 25220
rect 8392 25162 8444 25168
rect 8404 24818 8432 25162
rect 8680 24954 8708 25298
rect 8864 25158 8892 26794
rect 8956 26466 8984 26862
rect 9036 26512 9088 26518
rect 8956 26460 9036 26466
rect 8956 26454 9088 26460
rect 8956 26438 9076 26454
rect 9312 26444 9364 26450
rect 8956 26382 8984 26438
rect 9312 26386 9364 26392
rect 8944 26376 8996 26382
rect 8944 26318 8996 26324
rect 9128 26376 9180 26382
rect 9128 26318 9180 26324
rect 9140 26042 9168 26318
rect 9036 26036 9088 26042
rect 9036 25978 9088 25984
rect 9128 26036 9180 26042
rect 9128 25978 9180 25984
rect 9048 25702 9076 25978
rect 9036 25696 9088 25702
rect 9036 25638 9088 25644
rect 9128 25424 9180 25430
rect 9128 25366 9180 25372
rect 8852 25152 8904 25158
rect 8852 25094 8904 25100
rect 8668 24948 8720 24954
rect 8668 24890 8720 24896
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8116 23316 8168 23322
rect 8116 23258 8168 23264
rect 8128 22710 8156 23258
rect 8116 22704 8168 22710
rect 8116 22646 8168 22652
rect 8208 22636 8260 22642
rect 8208 22578 8260 22584
rect 8220 22166 8248 22578
rect 8404 22438 8432 24754
rect 8668 23520 8720 23526
rect 8668 23462 8720 23468
rect 8680 23118 8708 23462
rect 8668 23112 8720 23118
rect 8668 23054 8720 23060
rect 8864 23050 8892 25094
rect 9140 24954 9168 25366
rect 9128 24948 9180 24954
rect 9128 24890 9180 24896
rect 9324 24834 9352 26386
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 9140 24806 9352 24834
rect 8944 23724 8996 23730
rect 8944 23666 8996 23672
rect 8956 23322 8984 23666
rect 8944 23316 8996 23322
rect 8944 23258 8996 23264
rect 9140 23186 9168 24806
rect 9416 24750 9444 25842
rect 9220 24744 9272 24750
rect 9220 24686 9272 24692
rect 9404 24744 9456 24750
rect 9404 24686 9456 24692
rect 9232 24410 9260 24686
rect 9220 24404 9272 24410
rect 9220 24346 9272 24352
rect 9416 23322 9444 24686
rect 9496 23656 9548 23662
rect 9496 23598 9548 23604
rect 9404 23316 9456 23322
rect 9324 23276 9404 23304
rect 9220 23248 9272 23254
rect 9220 23190 9272 23196
rect 8944 23180 8996 23186
rect 8944 23122 8996 23128
rect 9128 23180 9180 23186
rect 9128 23122 9180 23128
rect 8852 23044 8904 23050
rect 8852 22986 8904 22992
rect 8668 22976 8720 22982
rect 8668 22918 8720 22924
rect 8576 22704 8628 22710
rect 8576 22646 8628 22652
rect 8300 22432 8352 22438
rect 8300 22374 8352 22380
rect 8392 22432 8444 22438
rect 8392 22374 8444 22380
rect 8208 22160 8260 22166
rect 8208 22102 8260 22108
rect 7932 21956 7984 21962
rect 7932 21898 7984 21904
rect 7944 21554 7972 21898
rect 8220 21894 8248 22102
rect 8312 22098 8340 22374
rect 8300 22092 8352 22098
rect 8300 22034 8352 22040
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 7748 21548 7800 21554
rect 7748 21490 7800 21496
rect 7932 21548 7984 21554
rect 7932 21490 7984 21496
rect 8024 21480 8076 21486
rect 8024 21422 8076 21428
rect 8312 21434 8340 22034
rect 8588 21962 8616 22646
rect 8576 21956 8628 21962
rect 8576 21898 8628 21904
rect 8484 21548 8536 21554
rect 8484 21490 8536 21496
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 8036 21146 8064 21422
rect 8312 21406 8432 21434
rect 8300 21344 8352 21350
rect 8300 21286 8352 21292
rect 8024 21140 8076 21146
rect 8024 21082 8076 21088
rect 8312 20466 8340 21286
rect 8404 20942 8432 21406
rect 8496 21146 8524 21490
rect 8484 21140 8536 21146
rect 8484 21082 8536 21088
rect 8392 20936 8444 20942
rect 8392 20878 8444 20884
rect 8588 20806 8616 21898
rect 8680 21010 8708 22918
rect 8956 22438 8984 23122
rect 9036 23044 9088 23050
rect 9036 22986 9088 22992
rect 8944 22432 8996 22438
rect 8944 22374 8996 22380
rect 9048 21350 9076 22986
rect 9232 22642 9260 23190
rect 9324 22982 9352 23276
rect 9404 23258 9456 23264
rect 9508 23186 9536 23598
rect 9496 23180 9548 23186
rect 9496 23122 9548 23128
rect 9404 23112 9456 23118
rect 9404 23054 9456 23060
rect 9312 22976 9364 22982
rect 9312 22918 9364 22924
rect 9416 22778 9444 23054
rect 9404 22772 9456 22778
rect 9404 22714 9456 22720
rect 9128 22636 9180 22642
rect 9128 22578 9180 22584
rect 9220 22636 9272 22642
rect 9220 22578 9272 22584
rect 9140 22234 9168 22578
rect 9508 22574 9536 23122
rect 9600 23118 9628 28426
rect 9772 28416 9824 28422
rect 9772 28358 9824 28364
rect 9680 28144 9732 28150
rect 9680 28086 9732 28092
rect 9692 27606 9720 28086
rect 9680 27600 9732 27606
rect 9680 27542 9732 27548
rect 9784 26994 9812 28358
rect 9968 27878 9996 28494
rect 10784 28416 10836 28422
rect 10784 28358 10836 28364
rect 9956 27872 10008 27878
rect 9956 27814 10008 27820
rect 10508 27872 10560 27878
rect 10508 27814 10560 27820
rect 10600 27872 10652 27878
rect 10600 27814 10652 27820
rect 10324 27532 10376 27538
rect 10324 27474 10376 27480
rect 9864 27396 9916 27402
rect 9864 27338 9916 27344
rect 9876 27130 9904 27338
rect 9864 27124 9916 27130
rect 9864 27066 9916 27072
rect 9772 26988 9824 26994
rect 9772 26930 9824 26936
rect 9784 25974 9812 26930
rect 10336 26382 10364 27474
rect 10520 27470 10548 27814
rect 10612 27538 10640 27814
rect 10600 27532 10652 27538
rect 10600 27474 10652 27480
rect 10796 27470 10824 28358
rect 10508 27464 10560 27470
rect 10508 27406 10560 27412
rect 10784 27464 10836 27470
rect 10784 27406 10836 27412
rect 10416 26784 10468 26790
rect 10416 26726 10468 26732
rect 10428 26450 10456 26726
rect 10416 26444 10468 26450
rect 10416 26386 10468 26392
rect 10324 26376 10376 26382
rect 10324 26318 10376 26324
rect 9772 25968 9824 25974
rect 9772 25910 9824 25916
rect 9680 25832 9732 25838
rect 9680 25774 9732 25780
rect 9692 25498 9720 25774
rect 9680 25492 9732 25498
rect 9680 25434 9732 25440
rect 9784 25362 9812 25910
rect 10048 25696 10100 25702
rect 10048 25638 10100 25644
rect 9772 25356 9824 25362
rect 9772 25298 9824 25304
rect 9956 25288 10008 25294
rect 9956 25230 10008 25236
rect 9968 24886 9996 25230
rect 9956 24880 10008 24886
rect 9956 24822 10008 24828
rect 9680 24200 9732 24206
rect 9680 24142 9732 24148
rect 9692 23594 9720 24142
rect 9680 23588 9732 23594
rect 9680 23530 9732 23536
rect 9588 23112 9640 23118
rect 9588 23054 9640 23060
rect 9588 22976 9640 22982
rect 9692 22964 9720 23530
rect 9968 23526 9996 24822
rect 10060 24750 10088 25638
rect 10336 25498 10364 26318
rect 10324 25492 10376 25498
rect 10324 25434 10376 25440
rect 10416 25356 10468 25362
rect 10416 25298 10468 25304
rect 10140 25220 10192 25226
rect 10140 25162 10192 25168
rect 10152 24818 10180 25162
rect 10428 24886 10456 25298
rect 10416 24880 10468 24886
rect 10416 24822 10468 24828
rect 10140 24812 10192 24818
rect 10140 24754 10192 24760
rect 10048 24744 10100 24750
rect 10048 24686 10100 24692
rect 10060 24206 10088 24686
rect 10048 24200 10100 24206
rect 10048 24142 10100 24148
rect 10152 23730 10180 24754
rect 10232 24336 10284 24342
rect 10232 24278 10284 24284
rect 10140 23724 10192 23730
rect 10140 23666 10192 23672
rect 9772 23520 9824 23526
rect 9772 23462 9824 23468
rect 9956 23520 10008 23526
rect 9956 23462 10008 23468
rect 9784 23118 9812 23462
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 9772 22976 9824 22982
rect 9692 22936 9772 22964
rect 9588 22918 9640 22924
rect 9772 22918 9824 22924
rect 9600 22624 9628 22918
rect 9600 22596 9720 22624
rect 9496 22568 9548 22574
rect 9548 22516 9628 22522
rect 9496 22510 9628 22516
rect 9312 22500 9364 22506
rect 9508 22494 9628 22510
rect 9312 22442 9364 22448
rect 9220 22432 9272 22438
rect 9220 22374 9272 22380
rect 9128 22228 9180 22234
rect 9128 22170 9180 22176
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 9036 21344 9088 21350
rect 9036 21286 9088 21292
rect 8668 21004 8720 21010
rect 8668 20946 8720 20952
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 8956 20534 8984 21286
rect 9140 21010 9168 21966
rect 9232 21690 9260 22374
rect 9324 22098 9352 22442
rect 9404 22432 9456 22438
rect 9404 22374 9456 22380
rect 9496 22432 9548 22438
rect 9496 22374 9548 22380
rect 9312 22092 9364 22098
rect 9312 22034 9364 22040
rect 9220 21684 9272 21690
rect 9220 21626 9272 21632
rect 9416 21554 9444 22374
rect 9508 22098 9536 22374
rect 9496 22092 9548 22098
rect 9496 22034 9548 22040
rect 9600 21962 9628 22494
rect 9692 22098 9720 22596
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 9588 21956 9640 21962
rect 9588 21898 9640 21904
rect 9496 21888 9548 21894
rect 9496 21830 9548 21836
rect 9508 21690 9536 21830
rect 9496 21684 9548 21690
rect 9496 21626 9548 21632
rect 9404 21548 9456 21554
rect 9404 21490 9456 21496
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 9600 21350 9628 21490
rect 9588 21344 9640 21350
rect 9588 21286 9640 21292
rect 9128 21004 9180 21010
rect 9128 20946 9180 20952
rect 9140 20602 9168 20946
rect 9128 20596 9180 20602
rect 9128 20538 9180 20544
rect 8944 20528 8996 20534
rect 8944 20470 8996 20476
rect 9404 20528 9456 20534
rect 9404 20470 9456 20476
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 8484 20460 8536 20466
rect 8484 20402 8536 20408
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 8496 19242 8524 20402
rect 9416 19938 9444 20470
rect 9496 20392 9548 20398
rect 9496 20334 9548 20340
rect 9508 20058 9536 20334
rect 9496 20052 9548 20058
rect 9496 19994 9548 20000
rect 9416 19910 9536 19938
rect 9508 19854 9536 19910
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 8484 19236 8536 19242
rect 8484 19178 8536 19184
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 8496 18290 8524 19178
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 8496 17746 8524 18226
rect 8484 17740 8536 17746
rect 8484 17682 8536 17688
rect 8496 17270 8524 17682
rect 8484 17264 8536 17270
rect 8484 17206 8536 17212
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 7748 16720 7800 16726
rect 7748 16662 7800 16668
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 7288 15428 7340 15434
rect 7288 15370 7340 15376
rect 7300 15162 7328 15370
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 7760 14414 7788 16662
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7852 15502 7880 15982
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7852 14958 7880 15438
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7852 13938 7880 14894
rect 7944 14618 7972 17138
rect 8496 16658 8524 17206
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 9232 16590 9260 16934
rect 9220 16584 9272 16590
rect 9220 16526 9272 16532
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 8220 16182 8248 16390
rect 8208 16176 8260 16182
rect 8208 16118 8260 16124
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 8852 15972 8904 15978
rect 8852 15914 8904 15920
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 8036 14090 8064 15846
rect 8864 15094 8892 15914
rect 9128 15428 9180 15434
rect 9128 15370 9180 15376
rect 9140 15162 9168 15370
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 8852 15088 8904 15094
rect 8852 15030 8904 15036
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 8128 14618 8156 14962
rect 9232 14618 9260 16050
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 9220 14612 9272 14618
rect 9220 14554 9272 14560
rect 9324 14414 9352 15302
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 8036 14062 8156 14090
rect 9232 14074 9260 14282
rect 8128 13938 8156 14062
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 7840 13932 7892 13938
rect 7840 13874 7892 13880
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8220 13818 8248 13942
rect 8220 13790 8340 13818
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 6000 12436 6052 12442
rect 8036 12434 8064 13126
rect 8312 12918 8340 13790
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9312 13252 9364 13258
rect 9312 13194 9364 13200
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 6000 12378 6052 12384
rect 7944 12406 8064 12434
rect 8680 12434 8708 12854
rect 9324 12850 9352 13194
rect 9416 12918 9444 13330
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9140 12442 9168 12786
rect 8852 12436 8904 12442
rect 8680 12406 8800 12434
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 4620 11008 4672 11014
rect 4620 10950 4672 10956
rect 204 10804 256 10810
rect 204 10746 256 10752
rect 216 800 244 10746
rect 1860 10600 1912 10606
rect 1860 10542 1912 10548
rect 1308 8492 1360 8498
rect 1308 8434 1360 8440
rect 940 7404 992 7410
rect 940 7346 992 7352
rect 572 2440 624 2446
rect 572 2382 624 2388
rect 584 800 612 2382
rect 952 800 980 7346
rect 1320 800 1348 8434
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1780 7546 1808 7822
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1872 6914 1900 10542
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 2136 8900 2188 8906
rect 2136 8842 2188 8848
rect 1952 8288 2004 8294
rect 1952 8230 2004 8236
rect 1964 7886 1992 8230
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 1780 6886 1900 6914
rect 1780 6458 1808 6886
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 1584 2304 1636 2310
rect 1584 2246 1636 2252
rect 1596 1902 1624 2246
rect 1584 1896 1636 1902
rect 1584 1838 1636 1844
rect 1780 1630 1808 5646
rect 2056 4282 2084 8026
rect 2148 7002 2176 8842
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 2332 7546 2360 7754
rect 2976 7546 3004 9930
rect 3988 9654 4016 9998
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 4632 9586 4660 10950
rect 5460 10606 5488 11018
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4724 10062 4752 10406
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 5276 8974 5304 9318
rect 5552 8974 5580 9998
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 2136 6996 2188 7002
rect 2136 6938 2188 6944
rect 2964 6996 3016 7002
rect 2964 6938 3016 6944
rect 2976 6905 3004 6938
rect 2962 6896 3018 6905
rect 2962 6831 3018 6840
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 2964 6792 3016 6798
rect 3068 6769 3096 6802
rect 2964 6734 3016 6740
rect 3054 6760 3110 6769
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2424 5409 2452 6054
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 2686 5672 2742 5681
rect 2410 5400 2466 5409
rect 2410 5335 2466 5344
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2332 4826 2360 4966
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2608 4457 2636 5646
rect 2686 5607 2742 5616
rect 2700 4690 2728 5607
rect 2792 5545 2820 6190
rect 2872 6180 2924 6186
rect 2872 6122 2924 6128
rect 2884 5681 2912 6122
rect 2976 5817 3004 6734
rect 3054 6695 3110 6704
rect 3054 6216 3110 6225
rect 3054 6151 3110 6160
rect 2962 5808 3018 5817
rect 2962 5743 3018 5752
rect 2870 5672 2926 5681
rect 2870 5607 2926 5616
rect 3068 5574 3096 6151
rect 3056 5568 3108 5574
rect 2778 5536 2834 5545
rect 3056 5510 3108 5516
rect 2778 5471 2834 5480
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 2872 5296 2924 5302
rect 2870 5264 2872 5273
rect 2924 5264 2926 5273
rect 2780 5228 2832 5234
rect 2870 5199 2926 5208
rect 2780 5170 2832 5176
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2594 4448 2650 4457
rect 2594 4383 2650 4392
rect 2044 4276 2096 4282
rect 2044 4218 2096 4224
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 1964 1970 1992 3470
rect 1952 1964 2004 1970
rect 1952 1906 2004 1912
rect 2792 1698 2820 5170
rect 3068 4758 3096 5306
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 2872 4548 2924 4554
rect 2872 4490 2924 4496
rect 2884 3233 2912 4490
rect 2964 3460 3016 3466
rect 2964 3402 3016 3408
rect 2976 3369 3004 3402
rect 2962 3360 3018 3369
rect 2962 3295 3018 3304
rect 2870 3224 2926 3233
rect 2870 3159 2926 3168
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 2976 2990 3004 3130
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 3068 2553 3096 2994
rect 3054 2544 3110 2553
rect 3054 2479 3110 2488
rect 3160 2394 3188 8774
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 3516 7880 3568 7886
rect 3238 7848 3294 7857
rect 3516 7822 3568 7828
rect 3238 7783 3294 7792
rect 3252 4282 3280 7783
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3252 3505 3280 4082
rect 3238 3496 3294 3505
rect 3238 3431 3294 3440
rect 3344 2650 3372 6054
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3436 4282 3464 5170
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3422 2952 3478 2961
rect 3422 2887 3478 2896
rect 3436 2854 3464 2887
rect 3424 2848 3476 2854
rect 3424 2790 3476 2796
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3068 2366 3188 2394
rect 3068 1834 3096 2366
rect 3148 2304 3200 2310
rect 3148 2246 3200 2252
rect 3056 1828 3108 1834
rect 3056 1770 3108 1776
rect 2780 1692 2832 1698
rect 2780 1634 2832 1640
rect 1768 1624 1820 1630
rect 1768 1566 1820 1572
rect 3160 800 3188 2246
rect 3252 2106 3280 2586
rect 3240 2100 3292 2106
rect 3240 2042 3292 2048
rect 3528 800 3556 7822
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3620 6866 3648 7278
rect 3608 6860 3660 6866
rect 3660 6820 3740 6848
rect 3608 6802 3660 6808
rect 3606 5672 3662 5681
rect 3606 5607 3662 5616
rect 3620 5098 3648 5607
rect 3712 5234 3740 6820
rect 3896 6458 3924 7346
rect 3988 6458 4016 8434
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4618 8120 4674 8129
rect 4618 8055 4674 8064
rect 4632 8022 4660 8055
rect 4620 8016 4672 8022
rect 4620 7958 4672 7964
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4080 6798 4108 7482
rect 4356 7478 4384 7686
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 4724 7313 4752 7890
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4816 7410 4844 7686
rect 4908 7449 4936 8434
rect 4894 7440 4950 7449
rect 4804 7404 4856 7410
rect 4894 7375 4950 7384
rect 4804 7346 4856 7352
rect 4710 7304 4766 7313
rect 4620 7268 4672 7274
rect 4710 7239 4766 7248
rect 4620 7210 4672 7216
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 4528 6724 4580 6730
rect 4528 6666 4580 6672
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 4436 6384 4488 6390
rect 4436 6326 4488 6332
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3896 5914 3924 6258
rect 4068 6112 4120 6118
rect 4448 6100 4476 6326
rect 4540 6322 4568 6666
rect 4632 6322 4660 7210
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4448 6072 4660 6100
rect 4068 6054 4120 6060
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 4080 5692 4108 6054
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4632 5914 4660 6072
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4160 5704 4212 5710
rect 4080 5664 4160 5692
rect 4160 5646 4212 5652
rect 4618 5400 4674 5409
rect 4618 5335 4620 5344
rect 4672 5335 4674 5344
rect 4620 5306 4672 5312
rect 3700 5228 3752 5234
rect 4620 5228 4672 5234
rect 3752 5188 3832 5216
rect 3700 5170 3752 5176
rect 3608 5092 3660 5098
rect 3608 5034 3660 5040
rect 3606 4312 3662 4321
rect 3606 4247 3662 4256
rect 3620 2446 3648 4247
rect 3804 4214 3832 5188
rect 4620 5170 4672 5176
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4160 4752 4212 4758
rect 4158 4720 4160 4729
rect 4212 4720 4214 4729
rect 4158 4655 4214 4664
rect 3884 4616 3936 4622
rect 3882 4584 3884 4593
rect 3936 4584 3938 4593
rect 4632 4554 4660 5170
rect 3882 4519 3938 4528
rect 4068 4548 4120 4554
rect 4068 4490 4120 4496
rect 4620 4548 4672 4554
rect 4620 4490 4672 4496
rect 3700 4208 3752 4214
rect 3698 4176 3700 4185
rect 3792 4208 3844 4214
rect 3752 4176 3754 4185
rect 3792 4150 3844 4156
rect 3698 4111 3754 4120
rect 3792 4072 3844 4078
rect 3790 4040 3792 4049
rect 3844 4040 3846 4049
rect 3790 3975 3846 3984
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 3712 3641 3740 3674
rect 3698 3632 3754 3641
rect 3698 3567 3754 3576
rect 4080 3398 4108 4490
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4344 3460 4396 3466
rect 4344 3402 4396 3408
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 3804 1426 3832 2994
rect 3988 2514 4016 3334
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4264 3097 4292 3130
rect 4250 3088 4306 3097
rect 4160 3052 4212 3058
rect 4356 3074 4384 3402
rect 4632 3194 4660 4082
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4356 3046 4660 3074
rect 4250 3023 4306 3032
rect 4160 2994 4212 3000
rect 4172 2938 4200 2994
rect 4080 2910 4200 2938
rect 4080 2530 4108 2910
rect 4632 2825 4660 3046
rect 4618 2816 4674 2825
rect 4214 2748 4522 2768
rect 4618 2751 4674 2760
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 3976 2508 4028 2514
rect 4080 2502 4292 2530
rect 3976 2450 4028 2456
rect 3792 1420 3844 1426
rect 3792 1362 3844 1368
rect 3896 800 3924 2450
rect 4264 800 4292 2502
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4632 800 4660 2382
rect 4724 2310 4752 6394
rect 4804 6316 4856 6322
rect 4804 6258 4856 6264
rect 4816 2854 4844 6258
rect 4908 4321 4936 7375
rect 5000 5030 5028 8774
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5080 8424 5132 8430
rect 5078 8392 5080 8401
rect 5132 8392 5134 8401
rect 5078 8327 5134 8336
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 5092 6361 5120 7754
rect 5078 6352 5134 6361
rect 5078 6287 5134 6296
rect 5092 5642 5120 6287
rect 5080 5636 5132 5642
rect 5080 5578 5132 5584
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 5092 4622 5120 5306
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 4894 4312 4950 4321
rect 4894 4247 4950 4256
rect 5000 4146 5028 4558
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5080 4004 5132 4010
rect 5080 3946 5132 3952
rect 5092 3534 5120 3946
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4908 3058 4936 3334
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 4712 2304 4764 2310
rect 4712 2246 4764 2252
rect 5000 1902 5028 2382
rect 4988 1896 5040 1902
rect 4988 1838 5040 1844
rect 5184 1630 5212 8570
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 5276 7274 5304 8366
rect 5264 7268 5316 7274
rect 5264 7210 5316 7216
rect 5262 5808 5318 5817
rect 5262 5743 5318 5752
rect 5276 5250 5304 5743
rect 5368 5370 5396 8910
rect 5644 8634 5672 9318
rect 5920 8974 5948 11834
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5724 8560 5776 8566
rect 5630 8528 5686 8537
rect 5724 8502 5776 8508
rect 5630 8463 5632 8472
rect 5684 8463 5686 8472
rect 5632 8434 5684 8440
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5460 7721 5488 7822
rect 5632 7812 5684 7818
rect 5632 7754 5684 7760
rect 5446 7712 5502 7721
rect 5446 7647 5502 7656
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5276 5222 5396 5250
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5276 4622 5304 4966
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5264 3664 5316 3670
rect 5262 3632 5264 3641
rect 5316 3632 5318 3641
rect 5262 3567 5318 3576
rect 5368 2774 5396 5222
rect 5460 3754 5488 7142
rect 5644 6866 5672 7754
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5538 6488 5594 6497
rect 5538 6423 5594 6432
rect 5552 6322 5580 6423
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5552 4758 5580 6054
rect 5644 5370 5672 6598
rect 5736 6236 5764 8502
rect 5828 7834 5856 8910
rect 5828 7806 5948 7834
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5828 7546 5856 7686
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5816 6248 5868 6254
rect 5736 6208 5816 6236
rect 5816 6190 5868 6196
rect 5920 5658 5948 7806
rect 6012 6866 6040 12378
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6472 10810 6500 11698
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 6920 11144 6972 11150
rect 7104 11144 7156 11150
rect 6972 11104 7104 11132
rect 6920 11086 6972 11092
rect 7104 11086 7156 11092
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6932 10674 6960 10746
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6380 10266 6408 10610
rect 7024 10266 7052 10950
rect 7116 10674 7144 10950
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 5998 6760 6054 6769
rect 5998 6695 6054 6704
rect 5736 5630 5948 5658
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5632 5212 5684 5218
rect 5632 5154 5684 5160
rect 5644 4826 5672 5154
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 5736 3942 5764 5630
rect 5908 5568 5960 5574
rect 5908 5510 5960 5516
rect 6012 5522 6040 6695
rect 6104 6458 6132 7822
rect 6196 7478 6224 7822
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 6196 5778 6224 6734
rect 6288 5930 6316 8978
rect 6380 7410 6408 9522
rect 6460 8288 6512 8294
rect 6458 8256 6460 8265
rect 6644 8288 6696 8294
rect 6512 8256 6514 8265
rect 6644 8230 6696 8236
rect 6458 8191 6514 8200
rect 6460 7744 6512 7750
rect 6460 7686 6512 7692
rect 6472 7410 6500 7686
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6656 7206 6684 8230
rect 6932 7936 6960 9930
rect 7116 9722 7144 9998
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7208 9178 7236 11154
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 7300 10810 7328 11018
rect 7288 10804 7340 10810
rect 7288 10746 7340 10752
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7300 10198 7328 10610
rect 7288 10192 7340 10198
rect 7288 10134 7340 10140
rect 7300 10062 7328 10134
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7300 8906 7328 9998
rect 7380 9716 7432 9722
rect 7380 9658 7432 9664
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 7392 8498 7420 9658
rect 7484 8974 7512 11494
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7852 10810 7880 11086
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7576 10062 7604 10610
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7576 9042 7604 9998
rect 7944 9058 7972 12406
rect 8772 11830 8800 12406
rect 8852 12378 8904 12384
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 8864 11937 8892 12378
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8850 11928 8906 11937
rect 8850 11863 8906 11872
rect 8760 11824 8812 11830
rect 8760 11766 8812 11772
rect 8300 11280 8352 11286
rect 8300 11222 8352 11228
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 8036 9178 8064 11154
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8128 10266 8156 11086
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8220 10130 8248 10406
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 7564 9036 7616 9042
rect 7944 9030 8064 9058
rect 7564 8978 7616 8984
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 6840 7908 6960 7936
rect 6736 7880 6788 7886
rect 6840 7868 6868 7908
rect 6788 7840 6868 7868
rect 6736 7822 6788 7828
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6564 6769 6592 7142
rect 6550 6760 6606 6769
rect 6550 6695 6606 6704
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6472 6497 6500 6598
rect 6458 6488 6514 6497
rect 6458 6423 6514 6432
rect 6288 5902 6408 5930
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6092 5636 6144 5642
rect 6288 5624 6316 5714
rect 6144 5596 6316 5624
rect 6092 5578 6144 5584
rect 5814 5264 5870 5273
rect 5814 5199 5870 5208
rect 5828 5166 5856 5199
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5920 4622 5948 5510
rect 6012 5494 6132 5522
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5828 4196 5856 4558
rect 5908 4208 5960 4214
rect 5828 4168 5908 4196
rect 5908 4150 5960 4156
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5460 3726 5856 3754
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5644 3194 5672 3402
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5736 3058 5764 3402
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5368 2746 5764 2774
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 4988 1624 5040 1630
rect 4988 1566 5040 1572
rect 5172 1624 5224 1630
rect 5172 1566 5224 1572
rect 5000 800 5028 1566
rect 5368 800 5396 2586
rect 5736 800 5764 2746
rect 202 0 258 800
rect 570 0 626 800
rect 938 0 994 800
rect 1306 0 1362 800
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 5828 762 5856 3726
rect 5920 3534 5948 4150
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 5920 2990 5948 3470
rect 6012 3058 6040 4966
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 6104 2582 6132 5494
rect 6092 2576 6144 2582
rect 6092 2518 6144 2524
rect 6380 1442 6408 5902
rect 6472 5642 6500 6423
rect 6656 6322 6684 7142
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6840 6118 6868 6734
rect 7024 6322 7052 8434
rect 7288 6384 7340 6390
rect 7380 6384 7432 6390
rect 7288 6326 7340 6332
rect 7378 6352 7380 6361
rect 7432 6352 7434 6361
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6460 5636 6512 5642
rect 6460 5578 6512 5584
rect 6472 5234 6500 5578
rect 6550 5264 6606 5273
rect 6460 5228 6512 5234
rect 6550 5199 6606 5208
rect 6460 5170 6512 5176
rect 6564 5114 6592 5199
rect 6472 5086 6592 5114
rect 6472 3466 6500 5086
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6564 4146 6592 4558
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6656 3942 6684 4082
rect 6840 4010 6868 6054
rect 7300 5574 7328 6326
rect 7378 6287 7434 6296
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6932 4146 6960 5306
rect 7024 4826 7052 5510
rect 7104 5296 7156 5302
rect 7104 5238 7156 5244
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6828 4004 6880 4010
rect 6828 3946 6880 3952
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 7116 3738 7144 5238
rect 7300 4622 7328 5510
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7208 3738 7236 4014
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7300 3534 7328 4558
rect 7392 3670 7420 5170
rect 7484 5166 7512 8910
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7576 6866 7604 8298
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7668 7886 7696 8230
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7668 6934 7696 7822
rect 7656 6928 7708 6934
rect 7656 6870 7708 6876
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7562 6760 7618 6769
rect 7562 6695 7618 6704
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7380 3664 7432 3670
rect 7380 3606 7432 3612
rect 7392 3534 7420 3606
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 6656 2922 6684 3402
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 6748 2910 7052 2938
rect 6748 2774 6776 2910
rect 7024 2854 7052 2910
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 6472 2746 6776 2774
rect 6472 2650 6500 2746
rect 6932 2689 6960 2790
rect 6918 2680 6974 2689
rect 6460 2644 6512 2650
rect 7392 2650 7420 2994
rect 7576 2774 7604 6695
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7760 5914 7788 6054
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7668 4690 7696 4966
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 7576 2746 7696 2774
rect 6918 2615 6974 2624
rect 7380 2644 7432 2650
rect 6460 2586 6512 2592
rect 7380 2586 7432 2592
rect 6920 2576 6972 2582
rect 6920 2518 6972 2524
rect 6380 1414 6592 1442
rect 6104 870 6224 898
rect 6104 762 6132 870
rect 6196 800 6224 870
rect 6564 800 6592 1414
rect 6932 800 6960 2518
rect 7380 2508 7432 2514
rect 7380 2450 7432 2456
rect 7392 2310 7420 2450
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7288 2304 7340 2310
rect 7288 2246 7340 2252
rect 7380 2304 7432 2310
rect 7380 2246 7432 2252
rect 7300 800 7328 2246
rect 7484 2038 7512 2382
rect 7472 2032 7524 2038
rect 7472 1974 7524 1980
rect 7668 800 7696 2746
rect 7852 2378 7880 8774
rect 7932 6724 7984 6730
rect 7932 6666 7984 6672
rect 7944 5370 7972 6666
rect 8036 5953 8064 9030
rect 8128 8362 8156 9522
rect 8312 8498 8340 11222
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 8404 10266 8432 10610
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8772 9518 8800 11766
rect 8956 10674 8984 12038
rect 9404 11280 9456 11286
rect 9404 11222 9456 11228
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8852 10056 8904 10062
rect 8904 10004 9168 10010
rect 8852 9998 9168 10004
rect 8864 9982 9168 9998
rect 9140 9722 9168 9982
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8496 8566 8524 8774
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 8404 8265 8432 8434
rect 8390 8256 8446 8265
rect 8390 8191 8446 8200
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8128 7342 8156 7822
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 8022 5944 8078 5953
rect 8022 5879 8078 5888
rect 8022 5400 8078 5409
rect 7932 5364 7984 5370
rect 8022 5335 8024 5344
rect 7932 5306 7984 5312
rect 8076 5335 8078 5344
rect 8024 5306 8076 5312
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 7944 3602 7972 4762
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 8036 3194 8064 5170
rect 8128 4826 8156 7278
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8220 6089 8248 6734
rect 8404 6254 8432 8191
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8496 7478 8524 7686
rect 8484 7472 8536 7478
rect 8484 7414 8536 7420
rect 8482 6488 8538 6497
rect 8482 6423 8538 6432
rect 8496 6390 8524 6423
rect 8484 6384 8536 6390
rect 8484 6326 8536 6332
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8206 6080 8262 6089
rect 8206 6015 8262 6024
rect 8220 5914 8248 6015
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8206 5672 8262 5681
rect 8206 5607 8262 5616
rect 8220 4826 8248 5607
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8128 3194 8156 3674
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 8036 2582 8064 3130
rect 8220 2961 8248 4558
rect 8298 3632 8354 3641
rect 8298 3567 8354 3576
rect 8206 2952 8262 2961
rect 8206 2887 8262 2896
rect 8312 2854 8340 3567
rect 8588 3534 8616 8910
rect 8772 6798 8800 9454
rect 9036 8900 9088 8906
rect 9036 8842 9088 8848
rect 8944 7856 8996 7862
rect 8852 7812 8904 7818
rect 8944 7798 8996 7804
rect 8852 7754 8904 7760
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8680 6361 8708 6734
rect 8666 6352 8722 6361
rect 8666 6287 8668 6296
rect 8720 6287 8722 6296
rect 8668 6258 8720 6264
rect 8680 6227 8708 6258
rect 8864 6254 8892 7754
rect 8956 6390 8984 7798
rect 9048 7041 9076 8842
rect 9034 7032 9090 7041
rect 9034 6967 9090 6976
rect 9036 6724 9088 6730
rect 9036 6666 9088 6672
rect 8944 6384 8996 6390
rect 8944 6326 8996 6332
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 8942 5808 8998 5817
rect 8942 5743 8998 5752
rect 8956 5710 8984 5743
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8956 4690 8984 4966
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 9048 4026 9076 6666
rect 9140 5234 9168 9658
rect 9416 8906 9444 11222
rect 9508 9586 9536 19790
rect 9600 19718 9628 21286
rect 9588 19712 9640 19718
rect 9588 19654 9640 19660
rect 9784 19514 9812 22918
rect 9968 19990 9996 23462
rect 10244 22778 10272 24278
rect 10428 24274 10456 24822
rect 10416 24268 10468 24274
rect 10416 24210 10468 24216
rect 10520 23798 10548 27406
rect 11072 27334 11100 28494
rect 11060 27328 11112 27334
rect 11060 27270 11112 27276
rect 11256 27130 11284 28494
rect 11336 28484 11388 28490
rect 11336 28426 11388 28432
rect 11244 27124 11296 27130
rect 11244 27066 11296 27072
rect 10600 26988 10652 26994
rect 10600 26930 10652 26936
rect 10612 24818 10640 26930
rect 10692 26920 10744 26926
rect 10692 26862 10744 26868
rect 11152 26920 11204 26926
rect 11152 26862 11204 26868
rect 10704 26586 10732 26862
rect 11164 26586 11192 26862
rect 10692 26580 10744 26586
rect 10692 26522 10744 26528
rect 11152 26580 11204 26586
rect 11152 26522 11204 26528
rect 11348 26518 11376 28426
rect 11980 28076 12032 28082
rect 11980 28018 12032 28024
rect 11612 27328 11664 27334
rect 11612 27270 11664 27276
rect 11336 26512 11388 26518
rect 11336 26454 11388 26460
rect 10784 26444 10836 26450
rect 10784 26386 10836 26392
rect 10796 25906 10824 26386
rect 11624 26382 11652 27270
rect 11992 26586 12020 28018
rect 12256 27396 12308 27402
rect 12256 27338 12308 27344
rect 12164 26920 12216 26926
rect 12164 26862 12216 26868
rect 11980 26580 12032 26586
rect 11980 26522 12032 26528
rect 11336 26376 11388 26382
rect 11336 26318 11388 26324
rect 11520 26376 11572 26382
rect 11520 26318 11572 26324
rect 11612 26376 11664 26382
rect 11612 26318 11664 26324
rect 11348 26042 11376 26318
rect 11336 26036 11388 26042
rect 11336 25978 11388 25984
rect 11532 25974 11560 26318
rect 11520 25968 11572 25974
rect 11520 25910 11572 25916
rect 10784 25900 10836 25906
rect 10784 25842 10836 25848
rect 10796 25770 10824 25842
rect 10784 25764 10836 25770
rect 10784 25706 10836 25712
rect 10692 25492 10744 25498
rect 10692 25434 10744 25440
rect 10704 24818 10732 25434
rect 11624 25226 11652 26318
rect 12176 25498 12204 26862
rect 12268 26042 12296 27338
rect 12440 26376 12492 26382
rect 12440 26318 12492 26324
rect 12348 26240 12400 26246
rect 12346 26208 12348 26217
rect 12400 26208 12402 26217
rect 12346 26143 12402 26152
rect 12452 26042 12480 26318
rect 12544 26246 12572 31726
rect 14740 30048 14792 30054
rect 14740 29990 14792 29996
rect 14752 29850 14780 29990
rect 14740 29844 14792 29850
rect 14740 29786 14792 29792
rect 14648 29708 14700 29714
rect 14648 29650 14700 29656
rect 14660 29238 14688 29650
rect 14740 29640 14792 29646
rect 14740 29582 14792 29588
rect 14648 29232 14700 29238
rect 14648 29174 14700 29180
rect 13084 29164 13136 29170
rect 13084 29106 13136 29112
rect 14464 29164 14516 29170
rect 14464 29106 14516 29112
rect 12624 29096 12676 29102
rect 12624 29038 12676 29044
rect 12532 26240 12584 26246
rect 12532 26182 12584 26188
rect 12256 26036 12308 26042
rect 12440 26036 12492 26042
rect 12308 25996 12388 26024
rect 12256 25978 12308 25984
rect 12360 25770 12388 25996
rect 12440 25978 12492 25984
rect 12348 25764 12400 25770
rect 12348 25706 12400 25712
rect 12164 25492 12216 25498
rect 12164 25434 12216 25440
rect 11796 25288 11848 25294
rect 12176 25242 12204 25434
rect 12360 25294 12388 25706
rect 11796 25230 11848 25236
rect 11612 25220 11664 25226
rect 11612 25162 11664 25168
rect 10600 24812 10652 24818
rect 10600 24754 10652 24760
rect 10692 24812 10744 24818
rect 10692 24754 10744 24760
rect 10612 24410 10640 24754
rect 10600 24404 10652 24410
rect 10600 24346 10652 24352
rect 10704 24290 10732 24754
rect 11520 24608 11572 24614
rect 11520 24550 11572 24556
rect 11612 24608 11664 24614
rect 11612 24550 11664 24556
rect 10968 24404 11020 24410
rect 10968 24346 11020 24352
rect 10612 24262 10732 24290
rect 10612 24206 10640 24262
rect 10600 24200 10652 24206
rect 10600 24142 10652 24148
rect 10600 24064 10652 24070
rect 10600 24006 10652 24012
rect 10508 23792 10560 23798
rect 10508 23734 10560 23740
rect 10416 23520 10468 23526
rect 10416 23462 10468 23468
rect 10232 22772 10284 22778
rect 10232 22714 10284 22720
rect 10428 22574 10456 23462
rect 10520 22778 10548 23734
rect 10508 22772 10560 22778
rect 10508 22714 10560 22720
rect 10508 22636 10560 22642
rect 10508 22578 10560 22584
rect 10416 22568 10468 22574
rect 10416 22510 10468 22516
rect 10520 22030 10548 22578
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 10416 21412 10468 21418
rect 10416 21354 10468 21360
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 9956 19984 10008 19990
rect 9956 19926 10008 19932
rect 10152 19854 10180 21286
rect 10428 21010 10456 21354
rect 10416 21004 10468 21010
rect 10416 20946 10468 20952
rect 10520 20942 10548 21966
rect 10508 20936 10560 20942
rect 10508 20878 10560 20884
rect 10520 20602 10548 20878
rect 10612 20602 10640 24006
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 10692 21480 10744 21486
rect 10692 21422 10744 21428
rect 10508 20596 10560 20602
rect 10508 20538 10560 20544
rect 10600 20596 10652 20602
rect 10600 20538 10652 20544
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 10244 19378 10272 20402
rect 10704 20058 10732 21422
rect 10796 21350 10824 21830
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10796 20058 10824 20402
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10508 19440 10560 19446
rect 10508 19382 10560 19388
rect 10232 19372 10284 19378
rect 10232 19314 10284 19320
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 9784 18970 9812 19110
rect 10244 18970 10272 19314
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 10232 18964 10284 18970
rect 10232 18906 10284 18912
rect 10520 18766 10548 19382
rect 10612 19378 10640 19790
rect 10692 19780 10744 19786
rect 10692 19722 10744 19728
rect 10704 19378 10732 19722
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10612 19174 10640 19314
rect 10600 19168 10652 19174
rect 10796 19122 10824 19994
rect 10888 19446 10916 20402
rect 10876 19440 10928 19446
rect 10876 19382 10928 19388
rect 10980 19310 11008 24346
rect 11532 24274 11560 24550
rect 11624 24274 11652 24550
rect 11808 24342 11836 25230
rect 11992 25214 12204 25242
rect 12348 25288 12400 25294
rect 12348 25230 12400 25236
rect 12256 25220 12308 25226
rect 11992 25158 12020 25214
rect 12256 25162 12308 25168
rect 11980 25152 12032 25158
rect 11980 25094 12032 25100
rect 11796 24336 11848 24342
rect 11796 24278 11848 24284
rect 11520 24268 11572 24274
rect 11520 24210 11572 24216
rect 11612 24268 11664 24274
rect 11612 24210 11664 24216
rect 11520 23724 11572 23730
rect 11624 23712 11652 24210
rect 12268 24206 12296 25162
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 12256 24200 12308 24206
rect 12256 24142 12308 24148
rect 11716 23730 11744 24142
rect 11888 24064 11940 24070
rect 11888 24006 11940 24012
rect 12348 24064 12400 24070
rect 12348 24006 12400 24012
rect 11900 23866 11928 24006
rect 11888 23860 11940 23866
rect 11888 23802 11940 23808
rect 11572 23684 11652 23712
rect 11704 23724 11756 23730
rect 11520 23666 11572 23672
rect 11704 23666 11756 23672
rect 11336 23656 11388 23662
rect 11336 23598 11388 23604
rect 11348 23322 11376 23598
rect 11612 23520 11664 23526
rect 11612 23462 11664 23468
rect 11152 23316 11204 23322
rect 11152 23258 11204 23264
rect 11336 23316 11388 23322
rect 11336 23258 11388 23264
rect 11164 22778 11192 23258
rect 11520 23248 11572 23254
rect 11520 23190 11572 23196
rect 11152 22772 11204 22778
rect 11152 22714 11204 22720
rect 11060 22500 11112 22506
rect 11060 22442 11112 22448
rect 11072 22166 11100 22442
rect 11060 22160 11112 22166
rect 11060 22102 11112 22108
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 11072 21554 11100 21966
rect 11060 21548 11112 21554
rect 11060 21490 11112 21496
rect 11072 21146 11100 21490
rect 11060 21140 11112 21146
rect 11060 21082 11112 21088
rect 11164 20942 11192 22714
rect 11336 22636 11388 22642
rect 11336 22578 11388 22584
rect 11348 21486 11376 22578
rect 11532 22030 11560 23190
rect 11624 23118 11652 23462
rect 11900 23118 11928 23802
rect 11978 23624 12034 23633
rect 11978 23559 12034 23568
rect 11612 23112 11664 23118
rect 11612 23054 11664 23060
rect 11888 23112 11940 23118
rect 11888 23054 11940 23060
rect 11796 22976 11848 22982
rect 11796 22918 11848 22924
rect 11428 22024 11480 22030
rect 11428 21966 11480 21972
rect 11520 22024 11572 22030
rect 11520 21966 11572 21972
rect 11440 21842 11468 21966
rect 11440 21814 11744 21842
rect 11716 21690 11744 21814
rect 11704 21684 11756 21690
rect 11704 21626 11756 21632
rect 11336 21480 11388 21486
rect 11336 21422 11388 21428
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 11060 20324 11112 20330
rect 11060 20266 11112 20272
rect 11072 19854 11100 20266
rect 11716 20058 11744 21626
rect 11808 20534 11836 22918
rect 11900 22030 11928 23054
rect 11992 22642 12020 23559
rect 12256 23248 12308 23254
rect 12256 23190 12308 23196
rect 11980 22636 12032 22642
rect 11980 22578 12032 22584
rect 11888 22024 11940 22030
rect 11888 21966 11940 21972
rect 11888 21548 11940 21554
rect 11888 21490 11940 21496
rect 11796 20528 11848 20534
rect 11796 20470 11848 20476
rect 11900 20466 11928 21490
rect 11992 21418 12020 22578
rect 12072 21956 12124 21962
rect 12072 21898 12124 21904
rect 12084 21554 12112 21898
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 12164 21480 12216 21486
rect 12164 21422 12216 21428
rect 11980 21412 12032 21418
rect 11980 21354 12032 21360
rect 12176 21350 12204 21422
rect 12164 21344 12216 21350
rect 12164 21286 12216 21292
rect 11980 20868 12032 20874
rect 11980 20810 12032 20816
rect 11888 20460 11940 20466
rect 11888 20402 11940 20408
rect 11992 20262 12020 20810
rect 11980 20256 12032 20262
rect 11980 20198 12032 20204
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11060 19848 11112 19854
rect 11060 19790 11112 19796
rect 11796 19848 11848 19854
rect 11796 19790 11848 19796
rect 11808 19446 11836 19790
rect 11992 19496 12020 20198
rect 11992 19468 12112 19496
rect 11796 19440 11848 19446
rect 11796 19382 11848 19388
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 10600 19110 10652 19116
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10508 18760 10560 18766
rect 10508 18702 10560 18708
rect 10428 17882 10456 18702
rect 10612 18698 10640 19110
rect 10704 19094 10824 19122
rect 10600 18692 10652 18698
rect 10600 18634 10652 18640
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10416 17876 10468 17882
rect 10416 17818 10468 17824
rect 10520 17202 10548 18362
rect 10612 17338 10640 18634
rect 10704 18426 10732 19094
rect 11532 18970 11560 19314
rect 10784 18964 10836 18970
rect 10784 18906 10836 18912
rect 11520 18964 11572 18970
rect 11520 18906 11572 18912
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 10796 17542 10824 18906
rect 10876 18692 10928 18698
rect 10876 18634 10928 18640
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 10600 17332 10652 17338
rect 10600 17274 10652 17280
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10048 16516 10100 16522
rect 10048 16458 10100 16464
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 9692 16114 9720 16390
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9692 15502 9720 16050
rect 9784 15706 9812 16050
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9692 15026 9720 15438
rect 9876 15094 9904 15846
rect 10060 15162 10088 16458
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10336 15570 10364 15982
rect 10888 15978 10916 18634
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10980 17882 11008 18226
rect 10968 17876 11020 17882
rect 10968 17818 11020 17824
rect 11796 17672 11848 17678
rect 11796 17614 11848 17620
rect 11808 17542 11836 17614
rect 11980 17604 12032 17610
rect 11980 17546 12032 17552
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 10876 15972 10928 15978
rect 10876 15914 10928 15920
rect 11072 15910 11100 16186
rect 11060 15904 11112 15910
rect 11808 15881 11836 17478
rect 11900 16590 11928 17478
rect 11992 16794 12020 17546
rect 12084 17202 12112 19468
rect 12176 18970 12204 21286
rect 12268 20602 12296 23190
rect 12360 22982 12388 24006
rect 12532 23860 12584 23866
rect 12532 23802 12584 23808
rect 12440 23520 12492 23526
rect 12440 23462 12492 23468
rect 12452 23186 12480 23462
rect 12544 23322 12572 23802
rect 12532 23316 12584 23322
rect 12532 23258 12584 23264
rect 12636 23254 12664 29038
rect 12716 28144 12768 28150
rect 12716 28086 12768 28092
rect 12728 27538 12756 28086
rect 12716 27532 12768 27538
rect 12716 27474 12768 27480
rect 12992 27464 13044 27470
rect 12992 27406 13044 27412
rect 12808 27056 12860 27062
rect 12808 26998 12860 27004
rect 12820 24614 12848 26998
rect 13004 26382 13032 27406
rect 13096 27130 13124 29106
rect 13544 28416 13596 28422
rect 13544 28358 13596 28364
rect 13556 28014 13584 28358
rect 14188 28144 14240 28150
rect 14188 28086 14240 28092
rect 13544 28008 13596 28014
rect 13544 27950 13596 27956
rect 13556 27538 13584 27950
rect 14004 27872 14056 27878
rect 14004 27814 14056 27820
rect 13544 27532 13596 27538
rect 13544 27474 13596 27480
rect 13084 27124 13136 27130
rect 13084 27066 13136 27072
rect 13268 26988 13320 26994
rect 13268 26930 13320 26936
rect 13280 26858 13308 26930
rect 13268 26852 13320 26858
rect 13268 26794 13320 26800
rect 13280 26382 13308 26794
rect 12992 26376 13044 26382
rect 12992 26318 13044 26324
rect 13268 26376 13320 26382
rect 13268 26318 13320 26324
rect 13004 25838 13032 26318
rect 13280 25906 13308 26318
rect 13268 25900 13320 25906
rect 13268 25842 13320 25848
rect 12992 25832 13044 25838
rect 13176 25832 13228 25838
rect 13044 25792 13124 25820
rect 12992 25774 13044 25780
rect 12900 25356 12952 25362
rect 12900 25298 12952 25304
rect 12808 24608 12860 24614
rect 12808 24550 12860 24556
rect 12716 23588 12768 23594
rect 12716 23530 12768 23536
rect 12624 23248 12676 23254
rect 12624 23190 12676 23196
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12624 23112 12676 23118
rect 12624 23054 12676 23060
rect 12532 23044 12584 23050
rect 12532 22986 12584 22992
rect 12348 22976 12400 22982
rect 12348 22918 12400 22924
rect 12544 22794 12572 22986
rect 12452 22766 12572 22794
rect 12636 22778 12664 23054
rect 12728 22778 12756 23530
rect 12820 23089 12848 24550
rect 12912 24206 12940 25298
rect 12900 24200 12952 24206
rect 12900 24142 12952 24148
rect 13096 23730 13124 25792
rect 13176 25774 13228 25780
rect 13188 24342 13216 25774
rect 13360 25764 13412 25770
rect 13360 25706 13412 25712
rect 13268 25696 13320 25702
rect 13268 25638 13320 25644
rect 13280 25158 13308 25638
rect 13372 25158 13400 25706
rect 13268 25152 13320 25158
rect 13268 25094 13320 25100
rect 13360 25152 13412 25158
rect 13360 25094 13412 25100
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 13176 24336 13228 24342
rect 13176 24278 13228 24284
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 13176 23860 13228 23866
rect 13176 23802 13228 23808
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 13004 23633 13032 23666
rect 12990 23624 13046 23633
rect 12990 23559 13046 23568
rect 12900 23112 12952 23118
rect 12806 23080 12862 23089
rect 12900 23054 12952 23060
rect 12806 23015 12862 23024
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12624 22772 12676 22778
rect 12452 22094 12480 22766
rect 12624 22714 12676 22720
rect 12716 22772 12768 22778
rect 12716 22714 12768 22720
rect 12728 22624 12756 22714
rect 12820 22642 12848 22918
rect 12636 22596 12756 22624
rect 12808 22636 12860 22642
rect 12452 22066 12572 22094
rect 12544 22030 12572 22066
rect 12348 22024 12400 22030
rect 12348 21966 12400 21972
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12360 21622 12388 21966
rect 12348 21616 12400 21622
rect 12348 21558 12400 21564
rect 12348 21412 12400 21418
rect 12348 21354 12400 21360
rect 12360 21010 12388 21354
rect 12348 21004 12400 21010
rect 12348 20946 12400 20952
rect 12360 20602 12388 20946
rect 12256 20596 12308 20602
rect 12256 20538 12308 20544
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 12348 20256 12400 20262
rect 12348 20198 12400 20204
rect 12256 19780 12308 19786
rect 12256 19722 12308 19728
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12268 17678 12296 19722
rect 12360 18086 12388 20198
rect 12544 19514 12572 21966
rect 12636 21894 12664 22596
rect 12808 22578 12860 22584
rect 12714 22536 12770 22545
rect 12714 22471 12770 22480
rect 12728 22030 12756 22471
rect 12808 22228 12860 22234
rect 12808 22170 12860 22176
rect 12820 22030 12848 22170
rect 12912 22098 12940 23054
rect 13096 22964 13124 23666
rect 13188 23118 13216 23802
rect 13268 23588 13320 23594
rect 13268 23530 13320 23536
rect 13176 23112 13228 23118
rect 13176 23054 13228 23060
rect 13280 23050 13308 23530
rect 13268 23044 13320 23050
rect 13268 22986 13320 22992
rect 13096 22936 13216 22964
rect 13084 22704 13136 22710
rect 13084 22646 13136 22652
rect 12900 22092 12952 22098
rect 12900 22034 12952 22040
rect 12716 22024 12768 22030
rect 12716 21966 12768 21972
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 12624 21888 12676 21894
rect 12624 21830 12676 21836
rect 12900 21344 12952 21350
rect 12900 21286 12952 21292
rect 12912 20942 12940 21286
rect 12900 20936 12952 20942
rect 12900 20878 12952 20884
rect 12624 20868 12676 20874
rect 12624 20810 12676 20816
rect 12532 19508 12584 19514
rect 12532 19450 12584 19456
rect 12348 18080 12400 18086
rect 12348 18022 12400 18028
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 12072 17196 12124 17202
rect 12072 17138 12124 17144
rect 12256 17128 12308 17134
rect 12256 17070 12308 17076
rect 11980 16788 12032 16794
rect 11980 16730 12032 16736
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 12268 15910 12296 17070
rect 12256 15904 12308 15910
rect 11060 15846 11112 15852
rect 11794 15872 11850 15881
rect 12256 15846 12308 15852
rect 11794 15807 11850 15816
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 9864 15088 9916 15094
rect 9864 15030 9916 15036
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 10336 14482 10364 15506
rect 10784 15428 10836 15434
rect 10784 15370 10836 15376
rect 10796 15162 10824 15370
rect 12268 15366 12296 15846
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 11520 15088 11572 15094
rect 11520 15030 11572 15036
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10336 14074 10364 14418
rect 10520 14346 10548 14962
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10508 14340 10560 14346
rect 10508 14282 10560 14288
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10336 13394 10364 14010
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9692 12238 9720 13126
rect 9876 12986 9904 13194
rect 10520 12986 10548 14282
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10612 12434 10640 14214
rect 10704 12850 10732 14554
rect 10876 14340 10928 14346
rect 10876 14282 10928 14288
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10612 12406 10732 12434
rect 10140 12368 10192 12374
rect 10140 12310 10192 12316
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9784 11762 9812 12038
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9600 11014 9628 11494
rect 9968 11354 9996 12174
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9692 9654 9720 11018
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 9494 8664 9550 8673
rect 9494 8599 9550 8608
rect 9508 8498 9536 8599
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9324 8362 9352 8434
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9324 8090 9527 8106
rect 9324 8084 9548 8090
rect 9324 8078 9496 8084
rect 9324 8022 9352 8078
rect 9496 8026 9548 8032
rect 9312 8016 9364 8022
rect 9312 7958 9364 7964
rect 9404 8016 9456 8022
rect 9456 7964 9536 7970
rect 9404 7958 9536 7964
rect 9416 7942 9536 7958
rect 9312 7880 9364 7886
rect 9404 7880 9456 7886
rect 9312 7822 9364 7828
rect 9402 7848 9404 7857
rect 9456 7848 9458 7857
rect 9220 7200 9272 7206
rect 9324 7188 9352 7822
rect 9402 7783 9458 7792
rect 9508 7546 9536 7942
rect 9588 7744 9640 7750
rect 9586 7712 9588 7721
rect 9640 7712 9642 7721
rect 9586 7647 9642 7656
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9508 7410 9536 7482
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9402 7304 9458 7313
rect 9402 7239 9404 7248
rect 9456 7239 9458 7248
rect 9404 7210 9456 7216
rect 9272 7160 9352 7188
rect 9220 7142 9272 7148
rect 9232 7002 9260 7142
rect 9402 7032 9458 7041
rect 9220 6996 9272 7002
rect 9402 6967 9404 6976
rect 9220 6938 9272 6944
rect 9456 6967 9458 6976
rect 9404 6938 9456 6944
rect 9402 6896 9458 6905
rect 9402 6831 9458 6840
rect 9416 6798 9444 6831
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9588 6656 9640 6662
rect 9494 6624 9550 6633
rect 9588 6598 9640 6604
rect 9494 6559 9550 6568
rect 9508 6458 9536 6559
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9600 6118 9628 6598
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9692 5692 9720 9590
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 9876 9194 9904 9454
rect 9784 9166 9904 9194
rect 9784 8430 9812 9166
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9876 8090 9904 8502
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9784 7936 9812 8026
rect 9864 7948 9916 7954
rect 9784 7908 9864 7936
rect 9864 7890 9916 7896
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9784 7342 9812 7754
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9784 5817 9812 7278
rect 9968 6322 9996 10406
rect 10046 9480 10102 9489
rect 10046 9415 10102 9424
rect 10060 8974 10088 9415
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 10152 8906 10180 12310
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 10244 9654 10272 12242
rect 10704 12238 10732 12406
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 10138 8664 10194 8673
rect 10138 8599 10194 8608
rect 10152 8498 10180 8599
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10152 8362 10180 8434
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10244 7886 10272 9318
rect 10336 8634 10364 12106
rect 10428 11626 10456 12174
rect 10796 11898 10824 13194
rect 10888 11898 10916 14282
rect 11532 14006 11560 15030
rect 11716 14822 11744 15302
rect 12268 15162 12296 15302
rect 12360 15162 12388 18022
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12452 16182 12480 16390
rect 12440 16176 12492 16182
rect 12440 16118 12492 16124
rect 12636 16114 12664 20810
rect 13096 20602 13124 22646
rect 13188 22574 13216 22936
rect 13176 22568 13228 22574
rect 13176 22510 13228 22516
rect 13176 22432 13228 22438
rect 13176 22374 13228 22380
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 12716 20528 12768 20534
rect 12716 20470 12768 20476
rect 12728 19718 12756 20470
rect 12992 20460 13044 20466
rect 12992 20402 13044 20408
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12728 17202 12756 19654
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12820 17746 12848 18566
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12636 15706 12664 15846
rect 12820 15706 12848 16526
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12532 15496 12584 15502
rect 12438 15464 12494 15473
rect 12532 15438 12584 15444
rect 12438 15399 12440 15408
rect 12492 15399 12494 15408
rect 12440 15370 12492 15376
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 12544 14414 12572 15438
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 11520 14000 11572 14006
rect 11520 13942 11572 13948
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 10980 12238 11008 13874
rect 11428 13456 11480 13462
rect 11428 13398 11480 13404
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10416 11620 10468 11626
rect 10416 11562 10468 11568
rect 10428 10538 10456 11562
rect 10980 11150 11008 12174
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 11072 11014 11100 12854
rect 11440 11762 11468 13398
rect 11532 13258 11560 13942
rect 11520 13252 11572 13258
rect 11520 13194 11572 13200
rect 11532 12918 11560 13194
rect 11624 12986 11652 14350
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11716 13734 11744 14214
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11520 12912 11572 12918
rect 11520 12854 11572 12860
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11716 12442 11744 12582
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11900 11762 11928 13670
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 11348 10538 11376 11222
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11808 10810 11836 11018
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11808 10674 11836 10746
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 10416 10532 10468 10538
rect 10416 10474 10468 10480
rect 10968 10532 11020 10538
rect 10968 10474 11020 10480
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 10980 9994 11008 10474
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10612 8090 10640 9522
rect 10796 8673 10824 9522
rect 10980 8974 11008 9930
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11256 9586 11284 9862
rect 12084 9722 12112 10610
rect 12176 10198 12204 13262
rect 12452 13258 12480 13942
rect 12544 13530 12572 14350
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12440 13252 12492 13258
rect 12440 13194 12492 13200
rect 12268 13161 12296 13194
rect 12254 13152 12310 13161
rect 12254 13087 12310 13096
rect 12452 12918 12480 13194
rect 12636 12918 12664 13874
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12624 12912 12676 12918
rect 12624 12854 12676 12860
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 12346 11928 12402 11937
rect 12346 11863 12402 11872
rect 12360 11830 12388 11863
rect 12256 11824 12308 11830
rect 12256 11766 12308 11772
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 12268 11257 12296 11766
rect 12360 11354 12388 11766
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12254 11248 12310 11257
rect 12254 11183 12310 11192
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 12164 10192 12216 10198
rect 12164 10134 12216 10140
rect 12360 9926 12388 11154
rect 12452 11150 12480 12106
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12544 11898 12572 12038
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12530 11248 12586 11257
rect 12530 11183 12532 11192
rect 12584 11183 12586 11192
rect 12532 11154 12584 11160
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12636 11014 12664 12854
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 10130 12480 10406
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 11796 9648 11848 9654
rect 11794 9616 11796 9625
rect 11848 9616 11850 9625
rect 11244 9580 11296 9586
rect 11794 9551 11850 9560
rect 11244 9522 11296 9528
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10782 8664 10838 8673
rect 10782 8599 10838 8608
rect 10876 8560 10928 8566
rect 10796 8520 10876 8548
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10152 7750 10180 7822
rect 10048 7744 10100 7750
rect 10046 7712 10048 7721
rect 10140 7744 10192 7750
rect 10100 7712 10102 7721
rect 10140 7686 10192 7692
rect 10046 7647 10102 7656
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9770 5808 9826 5817
rect 9770 5743 9826 5752
rect 9968 5710 9996 6258
rect 10060 6118 10088 7482
rect 10152 7410 10180 7686
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10152 6458 10180 7346
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10244 6390 10272 7822
rect 10428 7546 10456 8026
rect 10508 7880 10560 7886
rect 10506 7848 10508 7857
rect 10560 7848 10562 7857
rect 10704 7818 10732 8298
rect 10506 7783 10562 7792
rect 10692 7812 10744 7818
rect 10692 7754 10744 7760
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10704 7206 10732 7754
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10600 6724 10652 6730
rect 10600 6666 10652 6672
rect 10612 6458 10640 6666
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10704 6458 10732 6598
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10232 6384 10284 6390
rect 10232 6326 10284 6332
rect 10796 6322 10824 8520
rect 10876 8502 10928 8508
rect 10980 7410 11008 8910
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10876 6724 10928 6730
rect 10876 6666 10928 6672
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10232 6180 10284 6186
rect 10152 6140 10232 6168
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 9772 5704 9824 5710
rect 9692 5664 9772 5692
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9600 5030 9628 5170
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9588 5024 9640 5030
rect 9692 5001 9720 5664
rect 9956 5704 10008 5710
rect 9772 5646 9824 5652
rect 9862 5672 9918 5681
rect 9956 5646 10008 5652
rect 9862 5607 9918 5616
rect 9770 5400 9826 5409
rect 9770 5335 9772 5344
rect 9824 5335 9826 5344
rect 9772 5306 9824 5312
rect 9876 5250 9904 5607
rect 10152 5556 10180 6140
rect 10232 6122 10284 6128
rect 10232 5840 10284 5846
rect 10232 5782 10284 5788
rect 10322 5808 10378 5817
rect 9784 5222 9904 5250
rect 9968 5528 10180 5556
rect 9784 5098 9812 5222
rect 9772 5092 9824 5098
rect 9772 5034 9824 5040
rect 9588 4966 9640 4972
rect 9678 4992 9734 5001
rect 8772 3998 9076 4026
rect 8772 3942 8800 3998
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 9048 3602 9076 3998
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 8024 2576 8076 2582
rect 8024 2518 8076 2524
rect 8128 2446 8156 2586
rect 8758 2544 8814 2553
rect 8758 2479 8814 2488
rect 8116 2440 8168 2446
rect 8208 2440 8260 2446
rect 8116 2382 8168 2388
rect 8206 2408 8208 2417
rect 8260 2408 8262 2417
rect 7840 2372 7892 2378
rect 8206 2343 8262 2352
rect 7840 2314 7892 2320
rect 8392 2100 8444 2106
rect 8392 2042 8444 2048
rect 8024 1420 8076 1426
rect 8024 1362 8076 1368
rect 8036 800 8064 1362
rect 8404 800 8432 2042
rect 8772 800 8800 2479
rect 8864 2106 8892 2926
rect 9048 2446 9076 2926
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 8852 2100 8904 2106
rect 8852 2042 8904 2048
rect 9140 800 9168 2790
rect 9232 2650 9260 4966
rect 9678 4927 9734 4936
rect 9968 4865 9996 5528
rect 10048 5296 10100 5302
rect 10048 5238 10100 5244
rect 10060 4978 10088 5238
rect 10244 5234 10272 5782
rect 10322 5743 10378 5752
rect 10336 5370 10364 5743
rect 10414 5536 10470 5545
rect 10414 5471 10470 5480
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10322 4992 10378 5001
rect 10060 4950 10272 4978
rect 10244 4865 10272 4950
rect 10322 4927 10378 4936
rect 9494 4856 9550 4865
rect 9312 4820 9364 4826
rect 9494 4791 9550 4800
rect 9954 4856 10010 4865
rect 9954 4791 10010 4800
rect 10230 4856 10286 4865
rect 10230 4791 10286 4800
rect 9312 4762 9364 4768
rect 9324 4321 9352 4762
rect 9508 4758 9536 4791
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 9772 4752 9824 4758
rect 9824 4712 9996 4740
rect 9772 4694 9824 4700
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9310 4312 9366 4321
rect 9310 4247 9366 4256
rect 9310 4040 9366 4049
rect 9310 3975 9366 3984
rect 9324 2854 9352 3975
rect 9416 3641 9444 4422
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 9508 3738 9536 4082
rect 9968 4026 9996 4712
rect 10336 4690 10364 4927
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10336 4214 10364 4626
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10428 4078 10456 5471
rect 10520 5409 10548 6258
rect 10888 6225 10916 6666
rect 10874 6216 10930 6225
rect 10874 6151 10930 6160
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10506 5400 10562 5409
rect 10506 5335 10562 5344
rect 10690 5400 10746 5409
rect 10690 5335 10746 5344
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10520 4570 10548 5170
rect 10704 5114 10732 5335
rect 10888 5234 10916 5510
rect 10966 5400 11022 5409
rect 10966 5335 10968 5344
rect 11020 5335 11022 5344
rect 10968 5306 11020 5312
rect 11060 5296 11112 5302
rect 11060 5238 11112 5244
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 10612 5098 10732 5114
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10600 5092 10732 5098
rect 10652 5086 10732 5092
rect 10600 5034 10652 5040
rect 10692 5024 10744 5030
rect 10980 5012 11008 5102
rect 10744 4984 11008 5012
rect 10692 4966 10744 4972
rect 10874 4584 10930 4593
rect 10520 4542 10732 4570
rect 10600 4480 10652 4486
rect 10600 4422 10652 4428
rect 9876 3998 9996 4026
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 9876 3942 9904 3998
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9402 3632 9458 3641
rect 9402 3567 9458 3576
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 9232 2514 9260 2586
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 9416 2446 9444 3470
rect 9876 3210 9904 3674
rect 9968 3670 9996 3878
rect 10612 3738 10640 4422
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 10336 3556 10548 3584
rect 10232 3528 10284 3534
rect 10336 3516 10364 3556
rect 10284 3488 10364 3516
rect 10414 3496 10470 3505
rect 10232 3470 10284 3476
rect 10048 3460 10100 3466
rect 10414 3431 10470 3440
rect 10048 3402 10100 3408
rect 10060 3210 10088 3402
rect 9876 3182 9996 3210
rect 10060 3182 10364 3210
rect 9968 3126 9996 3182
rect 9956 3120 10008 3126
rect 9586 3088 9642 3097
rect 9642 3046 9904 3074
rect 9956 3062 10008 3068
rect 10046 3088 10102 3097
rect 9586 3023 9642 3032
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9404 2440 9456 2446
rect 9310 2408 9366 2417
rect 9404 2382 9456 2388
rect 9310 2343 9366 2352
rect 9324 2310 9352 2343
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9508 800 9536 2790
rect 9876 800 9904 3046
rect 10046 3023 10048 3032
rect 10100 3023 10102 3032
rect 10232 3052 10284 3058
rect 10048 2994 10100 3000
rect 10232 2994 10284 3000
rect 10244 2922 10272 2994
rect 10232 2916 10284 2922
rect 10232 2858 10284 2864
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 10230 2816 10286 2825
rect 10152 2446 10180 2790
rect 10230 2751 10286 2760
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10244 800 10272 2751
rect 10336 2650 10364 3182
rect 10428 2774 10456 3431
rect 10520 3058 10548 3556
rect 10600 3460 10652 3466
rect 10704 3448 10732 4542
rect 10874 4519 10930 4528
rect 10782 4448 10838 4457
rect 10782 4383 10838 4392
rect 10652 3420 10732 3448
rect 10600 3402 10652 3408
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10612 2922 10640 3402
rect 10796 3126 10824 4383
rect 10784 3120 10836 3126
rect 10784 3062 10836 3068
rect 10600 2916 10652 2922
rect 10600 2858 10652 2864
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 10428 2746 10640 2774
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 10612 800 10640 2746
rect 10796 2689 10824 2790
rect 10888 2774 10916 4519
rect 11072 4128 11100 5238
rect 10980 4100 11100 4128
rect 10980 3369 11008 4100
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 10966 3360 11022 3369
rect 10966 3295 11022 3304
rect 11072 2990 11100 3946
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 10888 2746 11008 2774
rect 10782 2680 10838 2689
rect 10782 2615 10838 2624
rect 10980 800 11008 2746
rect 11164 1902 11192 9454
rect 11796 9444 11848 9450
rect 11796 9386 11848 9392
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11256 8498 11284 9318
rect 11808 8838 11836 9386
rect 12544 8906 12572 10950
rect 12728 10606 12756 14894
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12820 13394 12848 13874
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12820 11762 12848 12174
rect 13004 12170 13032 20402
rect 13096 19446 13124 20538
rect 13188 20058 13216 22374
rect 13372 22030 13400 24006
rect 13464 23798 13492 24754
rect 13452 23792 13504 23798
rect 13452 23734 13504 23740
rect 13464 22438 13492 23734
rect 13556 23730 13584 27474
rect 13728 26240 13780 26246
rect 13728 26182 13780 26188
rect 13740 25838 13768 26182
rect 13728 25832 13780 25838
rect 13728 25774 13780 25780
rect 14016 25430 14044 27814
rect 14096 27328 14148 27334
rect 14096 27270 14148 27276
rect 14108 26994 14136 27270
rect 14096 26988 14148 26994
rect 14096 26930 14148 26936
rect 14096 26512 14148 26518
rect 14096 26454 14148 26460
rect 14108 25906 14136 26454
rect 14200 25974 14228 28086
rect 14476 27130 14504 29106
rect 14660 28558 14688 29174
rect 14648 28552 14700 28558
rect 14648 28494 14700 28500
rect 14556 27872 14608 27878
rect 14556 27814 14608 27820
rect 14464 27124 14516 27130
rect 14464 27066 14516 27072
rect 14280 26784 14332 26790
rect 14280 26726 14332 26732
rect 14188 25968 14240 25974
rect 14188 25910 14240 25916
rect 14096 25900 14148 25906
rect 14096 25842 14148 25848
rect 14004 25424 14056 25430
rect 14004 25366 14056 25372
rect 14016 24750 14044 25366
rect 13728 24744 13780 24750
rect 13728 24686 13780 24692
rect 14004 24744 14056 24750
rect 14004 24686 14056 24692
rect 13636 24336 13688 24342
rect 13636 24278 13688 24284
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 13544 23520 13596 23526
rect 13544 23462 13596 23468
rect 13452 22432 13504 22438
rect 13452 22374 13504 22380
rect 13556 22234 13584 23462
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13542 22128 13598 22137
rect 13542 22063 13544 22072
rect 13596 22063 13598 22072
rect 13544 22034 13596 22040
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13268 21548 13320 21554
rect 13372 21536 13400 21966
rect 13452 21888 13504 21894
rect 13452 21830 13504 21836
rect 13320 21508 13400 21536
rect 13268 21490 13320 21496
rect 13360 20936 13412 20942
rect 13360 20878 13412 20884
rect 13176 20052 13228 20058
rect 13176 19994 13228 20000
rect 13372 19990 13400 20878
rect 13464 20262 13492 21830
rect 13556 21554 13584 22034
rect 13544 21548 13596 21554
rect 13544 21490 13596 21496
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13360 19984 13412 19990
rect 13360 19926 13412 19932
rect 13464 19854 13492 20198
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13084 19440 13136 19446
rect 13084 19382 13136 19388
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13084 18760 13136 18766
rect 13084 18702 13136 18708
rect 13096 18426 13124 18702
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 13556 18290 13584 19110
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 13268 18284 13320 18290
rect 13268 18226 13320 18232
rect 13544 18284 13596 18290
rect 13544 18226 13596 18232
rect 13096 16998 13124 18226
rect 13174 17776 13230 17785
rect 13174 17711 13230 17720
rect 13188 17678 13216 17711
rect 13176 17672 13228 17678
rect 13176 17614 13228 17620
rect 13280 17270 13308 18226
rect 13556 17678 13584 18226
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13372 17338 13400 17614
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13268 17264 13320 17270
rect 13268 17206 13320 17212
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 13372 16046 13400 17070
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 13096 15094 13124 15846
rect 13372 15502 13400 15982
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13358 15328 13414 15337
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 13176 14544 13228 14550
rect 13176 14486 13228 14492
rect 13188 13326 13216 14486
rect 13280 14414 13308 15302
rect 13358 15263 13414 15272
rect 13372 14414 13400 15263
rect 13556 14618 13584 16186
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13280 14006 13308 14350
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 13176 13320 13228 13326
rect 13176 13262 13228 13268
rect 13188 12986 13216 13262
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 13096 11762 13124 12242
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12728 10470 12756 10542
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12636 9450 12664 9998
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12728 9489 12756 9522
rect 12714 9480 12770 9489
rect 12624 9444 12676 9450
rect 12714 9415 12770 9424
rect 12624 9386 12676 9392
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11348 7886 11376 8774
rect 11702 8664 11758 8673
rect 11702 8599 11758 8608
rect 11716 8566 11744 8599
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 11532 7936 11560 8434
rect 12254 8120 12310 8129
rect 12254 8055 12310 8064
rect 12440 8084 12492 8090
rect 12268 8022 12296 8055
rect 12440 8026 12492 8032
rect 12256 8016 12308 8022
rect 12256 7958 12308 7964
rect 12452 7954 12480 8026
rect 11612 7948 11664 7954
rect 11532 7908 11612 7936
rect 11612 7890 11664 7896
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 11242 5808 11298 5817
rect 11242 5743 11298 5752
rect 11256 5710 11284 5743
rect 11348 5710 11376 7822
rect 12268 7002 12296 7822
rect 12348 7472 12400 7478
rect 12346 7440 12348 7449
rect 12400 7440 12402 7449
rect 12346 7375 12402 7384
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11440 5409 11468 6054
rect 11532 5778 11560 6054
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 11426 5400 11482 5409
rect 11336 5364 11388 5370
rect 11426 5335 11482 5344
rect 11336 5306 11388 5312
rect 11348 5273 11376 5306
rect 11334 5264 11390 5273
rect 11334 5199 11390 5208
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11244 4208 11296 4214
rect 11244 4150 11296 4156
rect 11256 2650 11284 4150
rect 11348 3738 11376 4966
rect 11518 4176 11574 4185
rect 11428 4140 11480 4146
rect 11518 4111 11574 4120
rect 11428 4082 11480 4088
rect 11336 3732 11388 3738
rect 11336 3674 11388 3680
rect 11348 3534 11376 3674
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11348 3058 11376 3470
rect 11440 3058 11468 4082
rect 11336 3052 11388 3058
rect 11336 2994 11388 3000
rect 11428 3052 11480 3058
rect 11428 2994 11480 3000
rect 11532 2774 11560 4111
rect 11624 4010 11652 6190
rect 11716 5846 11744 6258
rect 11992 6186 12020 6734
rect 12164 6724 12216 6730
rect 12164 6666 12216 6672
rect 11980 6180 12032 6186
rect 11980 6122 12032 6128
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11704 5840 11756 5846
rect 11704 5782 11756 5788
rect 11796 5772 11848 5778
rect 11796 5714 11848 5720
rect 11808 4826 11836 5714
rect 11900 5545 11928 5850
rect 12176 5846 12204 6666
rect 12268 5914 12296 6938
rect 12348 6928 12400 6934
rect 12346 6896 12348 6905
rect 12400 6896 12402 6905
rect 12346 6831 12402 6840
rect 12346 6352 12402 6361
rect 12346 6287 12348 6296
rect 12400 6287 12402 6296
rect 12348 6258 12400 6264
rect 12452 6225 12480 7346
rect 12438 6216 12494 6225
rect 12438 6151 12494 6160
rect 12346 6080 12402 6089
rect 12346 6015 12402 6024
rect 12360 5914 12388 6015
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 12544 5681 12572 7822
rect 12728 6458 12756 8434
rect 12820 6934 12848 11698
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12912 11218 12940 11494
rect 13096 11286 13124 11698
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 13280 10690 13308 13194
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13464 12442 13492 12582
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 12912 10674 13308 10690
rect 12900 10668 13308 10674
rect 12952 10662 13308 10668
rect 12900 10610 12952 10616
rect 12808 6928 12860 6934
rect 12808 6870 12860 6876
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12912 5846 12940 10610
rect 13648 10282 13676 24278
rect 13740 21010 13768 24686
rect 14016 24274 14044 24686
rect 14004 24268 14056 24274
rect 14004 24210 14056 24216
rect 14200 24138 14228 25910
rect 14292 24410 14320 26726
rect 14370 26208 14426 26217
rect 14370 26143 14426 26152
rect 14280 24404 14332 24410
rect 14280 24346 14332 24352
rect 14188 24132 14240 24138
rect 14188 24074 14240 24080
rect 14200 23730 14228 24074
rect 14188 23724 14240 23730
rect 14188 23666 14240 23672
rect 13820 23588 13872 23594
rect 13820 23530 13872 23536
rect 13832 21554 13860 23530
rect 13912 23248 13964 23254
rect 13912 23190 13964 23196
rect 13924 22438 13952 23190
rect 14004 22976 14056 22982
rect 14004 22918 14056 22924
rect 14016 22574 14044 22918
rect 14096 22704 14148 22710
rect 14096 22646 14148 22652
rect 14004 22568 14056 22574
rect 14004 22510 14056 22516
rect 13912 22432 13964 22438
rect 13912 22374 13964 22380
rect 13912 22160 13964 22166
rect 13912 22102 13964 22108
rect 13924 21690 13952 22102
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13728 21004 13780 21010
rect 13728 20946 13780 20952
rect 14108 20482 14136 22646
rect 14200 22166 14228 23666
rect 14280 23520 14332 23526
rect 14280 23462 14332 23468
rect 14292 22778 14320 23462
rect 14280 22772 14332 22778
rect 14280 22714 14332 22720
rect 14188 22160 14240 22166
rect 14188 22102 14240 22108
rect 14188 21888 14240 21894
rect 14188 21830 14240 21836
rect 14200 20874 14228 21830
rect 14188 20868 14240 20874
rect 14188 20810 14240 20816
rect 14016 20454 14136 20482
rect 13728 19984 13780 19990
rect 13728 19926 13780 19932
rect 13740 14346 13768 19926
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13832 18222 13860 18770
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 13832 17610 13860 18158
rect 13820 17604 13872 17610
rect 13820 17546 13872 17552
rect 13832 17134 13860 17546
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13832 16590 13860 17070
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 14016 16114 14044 20454
rect 14096 20392 14148 20398
rect 14096 20334 14148 20340
rect 14108 19242 14136 20334
rect 14384 19514 14412 26143
rect 14568 25362 14596 27814
rect 14660 26518 14688 28494
rect 14648 26512 14700 26518
rect 14648 26454 14700 26460
rect 14648 26376 14700 26382
rect 14648 26318 14700 26324
rect 14556 25356 14608 25362
rect 14556 25298 14608 25304
rect 14464 24948 14516 24954
rect 14464 24890 14516 24896
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14096 19236 14148 19242
rect 14096 19178 14148 19184
rect 14108 17678 14136 19178
rect 14384 18970 14412 19450
rect 14476 19174 14504 24890
rect 14556 24812 14608 24818
rect 14556 24754 14608 24760
rect 14568 24614 14596 24754
rect 14660 24750 14688 26318
rect 14648 24744 14700 24750
rect 14648 24686 14700 24692
rect 14556 24608 14608 24614
rect 14556 24550 14608 24556
rect 14568 22137 14596 24550
rect 14554 22128 14610 22137
rect 14554 22063 14610 22072
rect 14464 19168 14516 19174
rect 14516 19128 14596 19156
rect 14464 19110 14516 19116
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14384 18766 14412 18906
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14200 18193 14228 18226
rect 14186 18184 14242 18193
rect 14186 18119 14242 18128
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 14200 17678 14228 18022
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14004 16108 14056 16114
rect 14004 16050 14056 16056
rect 14016 14890 14044 16050
rect 14004 14884 14056 14890
rect 14004 14826 14056 14832
rect 14108 14482 14136 17614
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14292 14958 14320 15302
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 14384 14414 14412 18566
rect 14568 18290 14596 19128
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14476 16454 14504 18226
rect 14568 16590 14596 18226
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14752 16130 14780 29582
rect 15292 29572 15344 29578
rect 15292 29514 15344 29520
rect 14924 29504 14976 29510
rect 14924 29446 14976 29452
rect 14832 27328 14884 27334
rect 14832 27270 14884 27276
rect 14844 24886 14872 27270
rect 14936 26994 14964 29446
rect 15108 28484 15160 28490
rect 15108 28426 15160 28432
rect 15120 28218 15148 28426
rect 15108 28212 15160 28218
rect 15108 28154 15160 28160
rect 15304 28082 15332 29514
rect 15292 28076 15344 28082
rect 15292 28018 15344 28024
rect 15304 27538 15332 28018
rect 15292 27532 15344 27538
rect 15292 27474 15344 27480
rect 15200 27124 15252 27130
rect 15200 27066 15252 27072
rect 15016 27056 15068 27062
rect 15016 26998 15068 27004
rect 15108 27012 15160 27018
rect 14924 26988 14976 26994
rect 14924 26930 14976 26936
rect 14936 26790 14964 26930
rect 14924 26784 14976 26790
rect 14924 26726 14976 26732
rect 14924 26444 14976 26450
rect 14924 26386 14976 26392
rect 14936 25498 14964 26386
rect 14924 25492 14976 25498
rect 14924 25434 14976 25440
rect 15028 25430 15056 26998
rect 15212 26994 15240 27066
rect 15108 26954 15160 26960
rect 15200 26988 15252 26994
rect 15120 25498 15148 26954
rect 15200 26930 15252 26936
rect 15200 26852 15252 26858
rect 15200 26794 15252 26800
rect 15212 26518 15240 26794
rect 15200 26512 15252 26518
rect 15200 26454 15252 26460
rect 15304 26450 15332 27474
rect 15292 26444 15344 26450
rect 15292 26386 15344 26392
rect 15292 26308 15344 26314
rect 15292 26250 15344 26256
rect 15200 25764 15252 25770
rect 15200 25706 15252 25712
rect 15108 25492 15160 25498
rect 15108 25434 15160 25440
rect 15016 25424 15068 25430
rect 15016 25366 15068 25372
rect 15108 25356 15160 25362
rect 15108 25298 15160 25304
rect 14924 25152 14976 25158
rect 14924 25094 14976 25100
rect 14832 24880 14884 24886
rect 14832 24822 14884 24828
rect 14936 24138 14964 25094
rect 15120 24682 15148 25298
rect 15212 25294 15240 25706
rect 15200 25288 15252 25294
rect 15200 25230 15252 25236
rect 15212 24818 15240 25230
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15108 24676 15160 24682
rect 15108 24618 15160 24624
rect 15108 24336 15160 24342
rect 15108 24278 15160 24284
rect 14832 24132 14884 24138
rect 14832 24074 14884 24080
rect 14924 24132 14976 24138
rect 14924 24074 14976 24080
rect 14844 23322 14872 24074
rect 15120 23866 15148 24278
rect 15108 23860 15160 23866
rect 15108 23802 15160 23808
rect 15200 23792 15252 23798
rect 15200 23734 15252 23740
rect 14924 23724 14976 23730
rect 14924 23666 14976 23672
rect 14832 23316 14884 23322
rect 14832 23258 14884 23264
rect 14832 22976 14884 22982
rect 14936 22964 14964 23666
rect 15016 23656 15068 23662
rect 15068 23616 15148 23644
rect 15016 23598 15068 23604
rect 15120 23118 15148 23616
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 15016 22976 15068 22982
rect 14936 22936 15016 22964
rect 14832 22918 14884 22924
rect 15016 22918 15068 22924
rect 14844 22506 14872 22918
rect 14832 22500 14884 22506
rect 14832 22442 14884 22448
rect 14832 22228 14884 22234
rect 14832 22170 14884 22176
rect 14844 21690 14872 22170
rect 14924 22024 14976 22030
rect 14924 21966 14976 21972
rect 14832 21684 14884 21690
rect 14832 21626 14884 21632
rect 14844 21554 14872 21626
rect 14832 21548 14884 21554
rect 14832 21490 14884 21496
rect 14936 21350 14964 21966
rect 14924 21344 14976 21350
rect 14924 21286 14976 21292
rect 14832 20868 14884 20874
rect 14832 20810 14884 20816
rect 14844 20058 14872 20810
rect 14832 20052 14884 20058
rect 14832 19994 14884 20000
rect 15028 19990 15056 22918
rect 15120 22778 15148 23054
rect 15108 22772 15160 22778
rect 15108 22714 15160 22720
rect 15108 22636 15160 22642
rect 15108 22578 15160 22584
rect 15016 19984 15068 19990
rect 15016 19926 15068 19932
rect 14924 19440 14976 19446
rect 14922 19408 14924 19417
rect 14976 19408 14978 19417
rect 14922 19343 14978 19352
rect 15120 19292 15148 22578
rect 15212 21690 15240 23734
rect 15304 22778 15332 26250
rect 15396 24410 15424 46514
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 17960 33992 18012 33998
rect 17960 33934 18012 33940
rect 16948 33448 17000 33454
rect 16948 33390 17000 33396
rect 16856 32768 16908 32774
rect 16856 32710 16908 32716
rect 16868 32502 16896 32710
rect 16856 32496 16908 32502
rect 16856 32438 16908 32444
rect 16960 32434 16988 33390
rect 17972 33114 18000 33934
rect 20260 33924 20312 33930
rect 20260 33866 20312 33872
rect 19432 33856 19484 33862
rect 19432 33798 19484 33804
rect 18420 33516 18472 33522
rect 18420 33458 18472 33464
rect 18432 33114 18460 33458
rect 17960 33108 18012 33114
rect 17960 33050 18012 33056
rect 18420 33108 18472 33114
rect 18420 33050 18472 33056
rect 17408 32972 17460 32978
rect 17408 32914 17460 32920
rect 17040 32904 17092 32910
rect 17040 32846 17092 32852
rect 16672 32428 16724 32434
rect 16672 32370 16724 32376
rect 16948 32428 17000 32434
rect 16948 32370 17000 32376
rect 16580 31136 16632 31142
rect 16580 31078 16632 31084
rect 15568 29776 15620 29782
rect 15568 29718 15620 29724
rect 16592 29730 16620 31078
rect 16684 30190 16712 32370
rect 17052 32026 17080 32846
rect 17040 32020 17092 32026
rect 17040 31962 17092 31968
rect 17420 31822 17448 32914
rect 17684 32904 17736 32910
rect 17684 32846 17736 32852
rect 18512 32904 18564 32910
rect 18512 32846 18564 32852
rect 17696 32570 17724 32846
rect 17684 32564 17736 32570
rect 17684 32506 17736 32512
rect 18420 32224 18472 32230
rect 18420 32166 18472 32172
rect 17408 31816 17460 31822
rect 17408 31758 17460 31764
rect 16856 31340 16908 31346
rect 16856 31282 16908 31288
rect 16764 31136 16816 31142
rect 16764 31078 16816 31084
rect 16776 30394 16804 31078
rect 16868 30394 16896 31282
rect 17420 30870 17448 31758
rect 18432 31754 18460 32166
rect 18524 32026 18552 32846
rect 19444 32842 19472 33798
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 20272 33658 20300 33866
rect 20260 33652 20312 33658
rect 20260 33594 20312 33600
rect 19984 33312 20036 33318
rect 19984 33254 20036 33260
rect 19432 32836 19484 32842
rect 19432 32778 19484 32784
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19340 32428 19392 32434
rect 19340 32370 19392 32376
rect 19616 32428 19668 32434
rect 19616 32370 19668 32376
rect 19248 32360 19300 32366
rect 19248 32302 19300 32308
rect 18880 32224 18932 32230
rect 18880 32166 18932 32172
rect 18512 32020 18564 32026
rect 18512 31962 18564 31968
rect 18512 31816 18564 31822
rect 18512 31758 18564 31764
rect 18328 31748 18380 31754
rect 18328 31690 18380 31696
rect 18420 31748 18472 31754
rect 18420 31690 18472 31696
rect 17960 31680 18012 31686
rect 17960 31622 18012 31628
rect 17972 31346 18000 31622
rect 18340 31482 18368 31690
rect 18328 31476 18380 31482
rect 18328 31418 18380 31424
rect 18052 31408 18104 31414
rect 18052 31350 18104 31356
rect 17960 31340 18012 31346
rect 17960 31282 18012 31288
rect 17408 30864 17460 30870
rect 17408 30806 17460 30812
rect 16948 30592 17000 30598
rect 16948 30534 17000 30540
rect 16764 30388 16816 30394
rect 16764 30330 16816 30336
rect 16856 30388 16908 30394
rect 16856 30330 16908 30336
rect 16764 30252 16816 30258
rect 16764 30194 16816 30200
rect 16672 30184 16724 30190
rect 16672 30126 16724 30132
rect 16684 29850 16712 30126
rect 16672 29844 16724 29850
rect 16672 29786 16724 29792
rect 15580 28082 15608 29718
rect 16592 29702 16712 29730
rect 16684 29646 16712 29702
rect 16672 29640 16724 29646
rect 16672 29582 16724 29588
rect 16580 29572 16632 29578
rect 16580 29514 16632 29520
rect 15660 28960 15712 28966
rect 15660 28902 15712 28908
rect 15672 28082 15700 28902
rect 16592 28762 16620 29514
rect 16776 29306 16804 30194
rect 16764 29300 16816 29306
rect 16764 29242 16816 29248
rect 16960 29170 16988 30534
rect 17420 30054 17448 30806
rect 17408 30048 17460 30054
rect 17408 29990 17460 29996
rect 18064 29510 18092 31350
rect 18524 31346 18552 31758
rect 18892 31346 18920 32166
rect 19260 31822 19288 32302
rect 19248 31816 19300 31822
rect 19248 31758 19300 31764
rect 19260 31686 19288 31758
rect 19248 31680 19300 31686
rect 19248 31622 19300 31628
rect 18144 31340 18196 31346
rect 18144 31282 18196 31288
rect 18512 31340 18564 31346
rect 18512 31282 18564 31288
rect 18788 31340 18840 31346
rect 18788 31282 18840 31288
rect 18880 31340 18932 31346
rect 18880 31282 18932 31288
rect 18052 29504 18104 29510
rect 18052 29446 18104 29452
rect 18064 29170 18092 29446
rect 18156 29306 18184 31282
rect 18800 30734 18828 31282
rect 18236 30728 18288 30734
rect 18236 30670 18288 30676
rect 18788 30728 18840 30734
rect 18788 30670 18840 30676
rect 18248 30054 18276 30670
rect 18328 30660 18380 30666
rect 18328 30602 18380 30608
rect 18236 30048 18288 30054
rect 18236 29990 18288 29996
rect 18248 29510 18276 29990
rect 18340 29850 18368 30602
rect 18800 30258 18828 30670
rect 18788 30252 18840 30258
rect 18788 30194 18840 30200
rect 18512 30184 18564 30190
rect 18512 30126 18564 30132
rect 18328 29844 18380 29850
rect 18328 29786 18380 29792
rect 18236 29504 18288 29510
rect 18236 29446 18288 29452
rect 18144 29300 18196 29306
rect 18144 29242 18196 29248
rect 16948 29164 17000 29170
rect 16948 29106 17000 29112
rect 18052 29164 18104 29170
rect 18052 29106 18104 29112
rect 16672 29028 16724 29034
rect 16672 28970 16724 28976
rect 16580 28756 16632 28762
rect 16580 28698 16632 28704
rect 15844 28620 15896 28626
rect 15844 28562 15896 28568
rect 15568 28076 15620 28082
rect 15568 28018 15620 28024
rect 15660 28076 15712 28082
rect 15660 28018 15712 28024
rect 15568 27940 15620 27946
rect 15568 27882 15620 27888
rect 15476 26988 15528 26994
rect 15476 26930 15528 26936
rect 15488 25888 15516 26930
rect 15580 26926 15608 27882
rect 15856 27674 15884 28562
rect 16580 28552 16632 28558
rect 16684 28540 16712 28970
rect 16632 28512 16712 28540
rect 16580 28494 16632 28500
rect 16028 28416 16080 28422
rect 16028 28358 16080 28364
rect 16040 28150 16068 28358
rect 16028 28144 16080 28150
rect 16028 28086 16080 28092
rect 15936 28076 15988 28082
rect 15936 28018 15988 28024
rect 15844 27668 15896 27674
rect 15844 27610 15896 27616
rect 15856 27130 15884 27610
rect 15844 27124 15896 27130
rect 15844 27066 15896 27072
rect 15948 26994 15976 28018
rect 16488 27464 16540 27470
rect 16488 27406 16540 27412
rect 16120 27396 16172 27402
rect 16120 27338 16172 27344
rect 15936 26988 15988 26994
rect 15936 26930 15988 26936
rect 15568 26920 15620 26926
rect 15568 26862 15620 26868
rect 16028 26920 16080 26926
rect 16028 26862 16080 26868
rect 15580 26353 15608 26862
rect 15844 26580 15896 26586
rect 15844 26522 15896 26528
rect 15856 26489 15884 26522
rect 15842 26480 15898 26489
rect 15842 26415 15898 26424
rect 15844 26376 15896 26382
rect 15566 26344 15622 26353
rect 15844 26318 15896 26324
rect 15934 26344 15990 26353
rect 15566 26279 15622 26288
rect 15856 26042 15884 26318
rect 15934 26279 15990 26288
rect 15844 26036 15896 26042
rect 15844 25978 15896 25984
rect 15488 25860 15608 25888
rect 15580 25498 15608 25860
rect 15568 25492 15620 25498
rect 15568 25434 15620 25440
rect 15476 25220 15528 25226
rect 15476 25162 15528 25168
rect 15752 25220 15804 25226
rect 15752 25162 15804 25168
rect 15384 24404 15436 24410
rect 15384 24346 15436 24352
rect 15384 24132 15436 24138
rect 15384 24074 15436 24080
rect 15396 23662 15424 24074
rect 15488 23798 15516 25162
rect 15764 24886 15792 25162
rect 15752 24880 15804 24886
rect 15752 24822 15804 24828
rect 15844 24812 15896 24818
rect 15844 24754 15896 24760
rect 15752 24200 15804 24206
rect 15752 24142 15804 24148
rect 15476 23792 15528 23798
rect 15476 23734 15528 23740
rect 15568 23792 15620 23798
rect 15568 23734 15620 23740
rect 15384 23656 15436 23662
rect 15384 23598 15436 23604
rect 15292 22772 15344 22778
rect 15292 22714 15344 22720
rect 15200 21684 15252 21690
rect 15200 21626 15252 21632
rect 14936 19264 15148 19292
rect 14936 18902 14964 19264
rect 15108 19168 15160 19174
rect 15028 19128 15108 19156
rect 14924 18896 14976 18902
rect 14924 18838 14976 18844
rect 14924 18760 14976 18766
rect 14922 18728 14924 18737
rect 14976 18728 14978 18737
rect 14922 18663 14978 18672
rect 14936 17610 14964 18663
rect 14924 17604 14976 17610
rect 14924 17546 14976 17552
rect 14832 16516 14884 16522
rect 14884 16476 14964 16504
rect 14832 16458 14884 16464
rect 14660 16102 14780 16130
rect 14462 15600 14518 15609
rect 14462 15535 14518 15544
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 13924 12986 13952 13670
rect 14096 13320 14148 13326
rect 14096 13262 14148 13268
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 13912 12708 13964 12714
rect 13912 12650 13964 12656
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13740 11830 13768 12310
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13832 12102 13860 12242
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 13832 11558 13860 12038
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13464 10254 13676 10282
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 13004 7392 13032 7822
rect 13096 7721 13124 8230
rect 13372 7886 13400 8774
rect 13464 8294 13492 10254
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13544 9988 13596 9994
rect 13544 9930 13596 9936
rect 13556 9625 13584 9930
rect 13542 9616 13598 9625
rect 13542 9551 13598 9560
rect 13648 9500 13676 10066
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13740 9654 13768 9862
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13728 9512 13780 9518
rect 13648 9472 13728 9500
rect 13728 9454 13780 9460
rect 13740 9178 13768 9454
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13634 8528 13690 8537
rect 13544 8492 13596 8498
rect 13740 8498 13768 8910
rect 13924 8634 13952 12650
rect 14108 12186 14136 13262
rect 14200 12434 14228 14350
rect 14476 13938 14504 15535
rect 14660 15450 14688 16102
rect 14740 15972 14792 15978
rect 14740 15914 14792 15920
rect 14568 15422 14688 15450
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14280 13728 14332 13734
rect 14280 13670 14332 13676
rect 14292 13530 14320 13670
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14292 12850 14320 13466
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14384 12646 14412 13806
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14200 12406 14412 12434
rect 14108 12170 14228 12186
rect 14108 12164 14240 12170
rect 14108 12158 14188 12164
rect 14188 12106 14240 12112
rect 14200 11354 14228 12106
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14108 9586 14136 9862
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13634 8463 13690 8472
rect 13728 8492 13780 8498
rect 13544 8434 13596 8440
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13082 7712 13138 7721
rect 13082 7647 13138 7656
rect 13084 7404 13136 7410
rect 13004 7364 13084 7392
rect 13084 7346 13136 7352
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 13004 6458 13032 6734
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 12992 6316 13044 6322
rect 13096 6304 13124 7346
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13188 6390 13216 6734
rect 13176 6384 13228 6390
rect 13176 6326 13228 6332
rect 13280 6322 13308 7142
rect 13044 6276 13124 6304
rect 13268 6316 13320 6322
rect 12992 6258 13044 6264
rect 13268 6258 13320 6264
rect 13372 6118 13400 7822
rect 13464 7342 13492 8230
rect 13556 8090 13584 8434
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13464 6905 13492 7142
rect 13450 6896 13506 6905
rect 13450 6831 13506 6840
rect 13556 6798 13584 7822
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 12900 5840 12952 5846
rect 12900 5782 12952 5788
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 12530 5672 12586 5681
rect 12820 5658 12848 5714
rect 13648 5710 13676 8463
rect 13728 8434 13780 8440
rect 13740 7750 13768 8434
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13636 5704 13688 5710
rect 12820 5630 13032 5658
rect 13636 5646 13688 5652
rect 12530 5607 12586 5616
rect 12900 5568 12952 5574
rect 11886 5536 11942 5545
rect 11886 5471 11942 5480
rect 12714 5536 12770 5545
rect 12900 5510 12952 5516
rect 12714 5471 12770 5480
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 11978 5128 12034 5137
rect 11978 5063 12034 5072
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11702 4720 11758 4729
rect 11702 4655 11758 4664
rect 11612 4004 11664 4010
rect 11612 3946 11664 3952
rect 11716 3534 11744 4655
rect 11808 3670 11836 4762
rect 11796 3664 11848 3670
rect 11796 3606 11848 3612
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 11992 3466 12020 5063
rect 12176 3738 12204 5170
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12254 4856 12310 4865
rect 12254 4791 12310 4800
rect 12268 4282 12296 4791
rect 12452 4622 12480 4966
rect 12530 4856 12586 4865
rect 12530 4791 12586 4800
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 11980 3460 12032 3466
rect 11980 3402 12032 3408
rect 12164 3392 12216 3398
rect 12162 3360 12164 3369
rect 12216 3360 12218 3369
rect 12162 3295 12218 3304
rect 12162 3224 12218 3233
rect 12162 3159 12218 3168
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11532 2746 11744 2774
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11336 1964 11388 1970
rect 11336 1906 11388 1912
rect 11152 1896 11204 1902
rect 11152 1838 11204 1844
rect 11348 800 11376 1906
rect 11716 1442 11744 2746
rect 11808 2650 11836 2994
rect 11796 2644 11848 2650
rect 11796 2586 11848 2592
rect 11716 1414 11836 1442
rect 11808 800 11836 1414
rect 12176 800 12204 3159
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 12360 2106 12388 2246
rect 12348 2100 12400 2106
rect 12348 2042 12400 2048
rect 12544 800 12572 4791
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12636 2514 12664 4558
rect 12728 2990 12756 5471
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12820 2774 12848 5102
rect 12912 4622 12940 5510
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12912 3194 12940 3334
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 13004 3058 13032 5630
rect 13740 5574 13768 7686
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13280 5234 13308 5510
rect 13358 5400 13414 5409
rect 13358 5335 13414 5344
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 13096 3738 13124 4558
rect 13268 4480 13320 4486
rect 13268 4422 13320 4428
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 13082 3632 13138 3641
rect 13082 3567 13138 3576
rect 13096 3534 13124 3567
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 13004 2854 13032 2994
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 12820 2746 12940 2774
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 12912 800 12940 2746
rect 13280 2582 13308 4422
rect 13372 2774 13400 5335
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13556 3890 13584 4082
rect 13648 4010 13676 4422
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 13832 3942 13860 6190
rect 13924 6118 13952 7822
rect 14004 6996 14056 7002
rect 14004 6938 14056 6944
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 14016 5846 14044 6938
rect 14186 6352 14242 6361
rect 14096 6316 14148 6322
rect 14186 6287 14242 6296
rect 14096 6258 14148 6264
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 14002 5672 14058 5681
rect 14002 5607 14004 5616
rect 14056 5607 14058 5616
rect 14004 5578 14056 5584
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 13912 4684 13964 4690
rect 13912 4626 13964 4632
rect 13924 4321 13952 4626
rect 13910 4312 13966 4321
rect 13910 4247 13966 4256
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 13820 3936 13872 3942
rect 13556 3862 13676 3890
rect 13820 3878 13872 3884
rect 13648 3738 13676 3862
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13544 3460 13596 3466
rect 13544 3402 13596 3408
rect 13728 3460 13780 3466
rect 13728 3402 13780 3408
rect 13556 3058 13584 3402
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13740 2922 13768 3402
rect 13832 3398 13860 3878
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13924 3097 13952 4082
rect 13910 3088 13966 3097
rect 13910 3023 13966 3032
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 13372 2746 13676 2774
rect 13268 2576 13320 2582
rect 13268 2518 13320 2524
rect 13268 1692 13320 1698
rect 13268 1634 13320 1640
rect 13280 800 13308 1634
rect 13648 800 13676 2746
rect 13924 2446 13952 2790
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 14016 2038 14044 4966
rect 14108 4622 14136 6258
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14108 4282 14136 4558
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 14108 3058 14136 3538
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 14200 2774 14228 6287
rect 14292 5030 14320 8978
rect 14280 5024 14332 5030
rect 14384 5012 14412 12406
rect 14476 11830 14504 13262
rect 14568 13258 14596 15422
rect 14752 15366 14780 15914
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14844 14074 14872 15438
rect 14936 14074 14964 16476
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 14648 14000 14700 14006
rect 14648 13942 14700 13948
rect 14660 13530 14688 13942
rect 14648 13524 14700 13530
rect 14648 13466 14700 13472
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14924 13252 14976 13258
rect 14924 13194 14976 13200
rect 14556 12368 14608 12374
rect 14556 12310 14608 12316
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14476 10062 14504 11086
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14464 8560 14516 8566
rect 14464 8502 14516 8508
rect 14476 7954 14504 8502
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 14568 6730 14596 12310
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14844 11558 14872 11698
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 14844 11082 14872 11494
rect 14936 11354 14964 13194
rect 15028 12442 15056 19128
rect 15108 19110 15160 19116
rect 15212 18850 15240 21626
rect 15304 21622 15332 22714
rect 15396 22642 15424 23598
rect 15476 23520 15528 23526
rect 15476 23462 15528 23468
rect 15488 22982 15516 23462
rect 15580 23186 15608 23734
rect 15764 23662 15792 24142
rect 15856 23798 15884 24754
rect 15844 23792 15896 23798
rect 15844 23734 15896 23740
rect 15752 23656 15804 23662
rect 15752 23598 15804 23604
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15568 23180 15620 23186
rect 15568 23122 15620 23128
rect 15476 22976 15528 22982
rect 15476 22918 15528 22924
rect 15568 22976 15620 22982
rect 15568 22918 15620 22924
rect 15580 22642 15608 22918
rect 15384 22636 15436 22642
rect 15384 22578 15436 22584
rect 15568 22636 15620 22642
rect 15568 22578 15620 22584
rect 15384 22500 15436 22506
rect 15384 22442 15436 22448
rect 15396 22234 15424 22442
rect 15384 22228 15436 22234
rect 15384 22170 15436 22176
rect 15580 22094 15608 22578
rect 15488 22066 15608 22094
rect 15384 21888 15436 21894
rect 15384 21830 15436 21836
rect 15396 21690 15424 21830
rect 15384 21684 15436 21690
rect 15384 21626 15436 21632
rect 15292 21616 15344 21622
rect 15292 21558 15344 21564
rect 15384 21480 15436 21486
rect 15384 21422 15436 21428
rect 15212 18822 15332 18850
rect 15304 18766 15332 18822
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 15200 18692 15252 18698
rect 15200 18634 15252 18640
rect 15108 17264 15160 17270
rect 15108 17206 15160 17212
rect 15120 16794 15148 17206
rect 15212 17202 15240 18634
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15108 16788 15160 16794
rect 15108 16730 15160 16736
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 15120 15434 15148 16390
rect 15108 15428 15160 15434
rect 15108 15370 15160 15376
rect 15108 14340 15160 14346
rect 15108 14282 15160 14288
rect 15120 13462 15148 14282
rect 15212 13802 15240 17138
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15304 16114 15332 16458
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 15304 15502 15332 16050
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 15108 13456 15160 13462
rect 15108 13398 15160 13404
rect 15396 13326 15424 21422
rect 15488 20534 15516 22066
rect 15568 21412 15620 21418
rect 15568 21354 15620 21360
rect 15580 20602 15608 21354
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15476 20528 15528 20534
rect 15476 20470 15528 20476
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15488 19854 15516 20198
rect 15476 19848 15528 19854
rect 15476 19790 15528 19796
rect 15476 19440 15528 19446
rect 15476 19382 15528 19388
rect 15488 18834 15516 19382
rect 15476 18828 15528 18834
rect 15476 18770 15528 18776
rect 15488 18290 15516 18770
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 15476 17876 15528 17882
rect 15476 17818 15528 17824
rect 15488 17134 15516 17818
rect 15580 17814 15608 20538
rect 15672 19446 15700 23258
rect 15948 22234 15976 26279
rect 16040 26042 16068 26862
rect 16132 26382 16160 27338
rect 16396 27328 16448 27334
rect 16396 27270 16448 27276
rect 16212 26988 16264 26994
rect 16212 26930 16264 26936
rect 16120 26376 16172 26382
rect 16120 26318 16172 26324
rect 16028 26036 16080 26042
rect 16028 25978 16080 25984
rect 16120 25832 16172 25838
rect 16120 25774 16172 25780
rect 16028 25492 16080 25498
rect 16028 25434 16080 25440
rect 16040 24138 16068 25434
rect 16132 25430 16160 25774
rect 16120 25424 16172 25430
rect 16120 25366 16172 25372
rect 16224 25158 16252 26930
rect 16302 26480 16358 26489
rect 16302 26415 16358 26424
rect 16316 25974 16344 26415
rect 16408 26382 16436 27270
rect 16500 26858 16528 27406
rect 16488 26852 16540 26858
rect 16488 26794 16540 26800
rect 16396 26376 16448 26382
rect 16396 26318 16448 26324
rect 16304 25968 16356 25974
rect 16304 25910 16356 25916
rect 16212 25152 16264 25158
rect 16212 25094 16264 25100
rect 16224 24818 16252 25094
rect 16212 24812 16264 24818
rect 16212 24754 16264 24760
rect 16120 24404 16172 24410
rect 16120 24346 16172 24352
rect 16132 24206 16160 24346
rect 16120 24200 16172 24206
rect 16120 24142 16172 24148
rect 16028 24132 16080 24138
rect 16028 24074 16080 24080
rect 15936 22228 15988 22234
rect 15936 22170 15988 22176
rect 16040 22094 16068 24074
rect 16120 23724 16172 23730
rect 16120 23666 16172 23672
rect 16132 23186 16160 23666
rect 16120 23180 16172 23186
rect 16120 23122 16172 23128
rect 15948 22066 16068 22094
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 15660 19440 15712 19446
rect 15660 19382 15712 19388
rect 15764 19378 15792 19654
rect 15856 19378 15884 21490
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 15856 19122 15884 19314
rect 15672 19094 15884 19122
rect 15568 17808 15620 17814
rect 15568 17750 15620 17756
rect 15672 17660 15700 19094
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 15580 17632 15700 17660
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15488 16046 15516 17070
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15488 15094 15516 15438
rect 15476 15088 15528 15094
rect 15476 15030 15528 15036
rect 15580 14346 15608 17632
rect 15658 17504 15714 17513
rect 15658 17439 15714 17448
rect 15672 17338 15700 17439
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15660 16992 15712 16998
rect 15660 16934 15712 16940
rect 15672 16794 15700 16934
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15764 16658 15792 18226
rect 15856 17746 15884 18702
rect 15844 17740 15896 17746
rect 15844 17682 15896 17688
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15660 16516 15712 16522
rect 15660 16458 15712 16464
rect 15672 16182 15700 16458
rect 15764 16250 15792 16594
rect 15856 16454 15884 17478
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 15660 16176 15712 16182
rect 15856 16130 15884 16390
rect 15660 16118 15712 16124
rect 15672 15706 15700 16118
rect 15764 16114 15884 16130
rect 15752 16108 15884 16114
rect 15804 16102 15884 16108
rect 15752 16050 15804 16056
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15488 13870 15516 14214
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 14936 11150 14964 11290
rect 14924 11144 14976 11150
rect 14924 11086 14976 11092
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14844 10538 14872 11018
rect 14832 10532 14884 10538
rect 14832 10474 14884 10480
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 14832 10056 14884 10062
rect 14832 9998 14884 10004
rect 14648 9988 14700 9994
rect 14648 9930 14700 9936
rect 14660 8430 14688 9930
rect 14844 9654 14872 9998
rect 14832 9648 14884 9654
rect 14832 9590 14884 9596
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 14936 8566 14964 8774
rect 14924 8560 14976 8566
rect 14924 8502 14976 8508
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 14924 8356 14976 8362
rect 14924 8298 14976 8304
rect 14936 7274 14964 8298
rect 15120 7886 15148 8910
rect 15212 8362 15240 10066
rect 15304 9586 15332 12378
rect 15396 11898 15424 13262
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15488 12850 15516 13126
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15672 12646 15700 13874
rect 15764 12918 15792 16050
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 15752 12912 15804 12918
rect 15752 12854 15804 12860
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15488 11626 15516 12174
rect 15672 11762 15700 12242
rect 15856 12238 15884 13466
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 15660 11620 15712 11626
rect 15660 11562 15712 11568
rect 15488 11150 15516 11562
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15672 10674 15700 11562
rect 15856 11286 15884 12174
rect 15948 11898 15976 22066
rect 16028 21616 16080 21622
rect 16028 21558 16080 21564
rect 16040 20618 16068 21558
rect 16040 20590 16160 20618
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 16040 18766 16068 19246
rect 16028 18760 16080 18766
rect 16028 18702 16080 18708
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 16040 17678 16068 18158
rect 16028 17672 16080 17678
rect 16028 17614 16080 17620
rect 16040 16182 16068 17614
rect 16132 17513 16160 20590
rect 16118 17504 16174 17513
rect 16118 17439 16174 17448
rect 16120 17060 16172 17066
rect 16224 17048 16252 24754
rect 16304 24404 16356 24410
rect 16304 24346 16356 24352
rect 16316 23322 16344 24346
rect 16396 24064 16448 24070
rect 16396 24006 16448 24012
rect 16304 23316 16356 23322
rect 16304 23258 16356 23264
rect 16408 23118 16436 24006
rect 16500 23730 16528 26794
rect 16592 25294 16620 28494
rect 17500 28484 17552 28490
rect 17500 28426 17552 28432
rect 16856 28076 16908 28082
rect 16856 28018 16908 28024
rect 17132 28076 17184 28082
rect 17132 28018 17184 28024
rect 16868 27402 16896 28018
rect 16856 27396 16908 27402
rect 16856 27338 16908 27344
rect 16868 26858 16896 27338
rect 16856 26852 16908 26858
rect 16856 26794 16908 26800
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16684 26217 16712 26318
rect 16868 26314 16896 26794
rect 16948 26784 17000 26790
rect 16948 26726 17000 26732
rect 16960 26450 16988 26726
rect 16948 26444 17000 26450
rect 16948 26386 17000 26392
rect 17038 26344 17094 26353
rect 16856 26308 16908 26314
rect 17038 26279 17040 26288
rect 16856 26250 16908 26256
rect 17092 26279 17094 26288
rect 17040 26250 17092 26256
rect 16670 26208 16726 26217
rect 16670 26143 16726 26152
rect 16764 25832 16816 25838
rect 16764 25774 16816 25780
rect 16580 25288 16632 25294
rect 16580 25230 16632 25236
rect 16488 23724 16540 23730
rect 16488 23666 16540 23672
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 16488 21684 16540 21690
rect 16488 21626 16540 21632
rect 16304 20800 16356 20806
rect 16304 20742 16356 20748
rect 16316 19990 16344 20742
rect 16304 19984 16356 19990
rect 16304 19926 16356 19932
rect 16172 17020 16252 17048
rect 16120 17002 16172 17008
rect 16316 16810 16344 19926
rect 16396 19848 16448 19854
rect 16396 19790 16448 19796
rect 16408 19378 16436 19790
rect 16396 19372 16448 19378
rect 16396 19314 16448 19320
rect 16408 17882 16436 19314
rect 16500 17898 16528 21626
rect 16580 21412 16632 21418
rect 16580 21354 16632 21360
rect 16592 20942 16620 21354
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16776 20466 16804 25774
rect 16948 24812 17000 24818
rect 16948 24754 17000 24760
rect 16960 24410 16988 24754
rect 17144 24614 17172 28018
rect 17316 27464 17368 27470
rect 17316 27406 17368 27412
rect 17224 26988 17276 26994
rect 17224 26930 17276 26936
rect 17236 26382 17264 26930
rect 17224 26376 17276 26382
rect 17224 26318 17276 26324
rect 17236 26246 17264 26318
rect 17224 26240 17276 26246
rect 17224 26182 17276 26188
rect 17224 25220 17276 25226
rect 17224 25162 17276 25168
rect 17132 24608 17184 24614
rect 17132 24550 17184 24556
rect 16948 24404 17000 24410
rect 16948 24346 17000 24352
rect 17040 24268 17092 24274
rect 17040 24210 17092 24216
rect 16948 24200 17000 24206
rect 16948 24142 17000 24148
rect 16856 24064 16908 24070
rect 16856 24006 16908 24012
rect 16868 23866 16896 24006
rect 16856 23860 16908 23866
rect 16856 23802 16908 23808
rect 16960 23526 16988 24142
rect 16948 23520 17000 23526
rect 16948 23462 17000 23468
rect 16856 23112 16908 23118
rect 16856 23054 16908 23060
rect 16868 22642 16896 23054
rect 16960 22778 16988 23462
rect 16948 22772 17000 22778
rect 16948 22714 17000 22720
rect 17052 22642 17080 24210
rect 17144 24070 17172 24550
rect 17236 24274 17264 25162
rect 17224 24268 17276 24274
rect 17224 24210 17276 24216
rect 17132 24064 17184 24070
rect 17132 24006 17184 24012
rect 17132 23656 17184 23662
rect 17132 23598 17184 23604
rect 17144 22982 17172 23598
rect 17236 23322 17264 24210
rect 17224 23316 17276 23322
rect 17224 23258 17276 23264
rect 17132 22976 17184 22982
rect 17132 22918 17184 22924
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 17040 22636 17092 22642
rect 17040 22578 17092 22584
rect 17144 22094 17172 22918
rect 17328 22438 17356 27406
rect 17408 26580 17460 26586
rect 17408 26522 17460 26528
rect 17420 25770 17448 26522
rect 17512 25838 17540 28426
rect 17776 28008 17828 28014
rect 17776 27950 17828 27956
rect 17788 27470 17816 27950
rect 17960 27872 18012 27878
rect 17960 27814 18012 27820
rect 17972 27674 18000 27814
rect 17960 27668 18012 27674
rect 17960 27610 18012 27616
rect 17776 27464 17828 27470
rect 17776 27406 17828 27412
rect 17960 27328 18012 27334
rect 17960 27270 18012 27276
rect 17972 27062 18000 27270
rect 17960 27056 18012 27062
rect 17960 26998 18012 27004
rect 17868 26988 17920 26994
rect 17868 26930 17920 26936
rect 17880 26586 17908 26930
rect 17868 26580 17920 26586
rect 17868 26522 17920 26528
rect 17972 26314 18000 26998
rect 17960 26308 18012 26314
rect 17960 26250 18012 26256
rect 17592 26240 17644 26246
rect 17592 26182 17644 26188
rect 17500 25832 17552 25838
rect 17500 25774 17552 25780
rect 17408 25764 17460 25770
rect 17408 25706 17460 25712
rect 17408 25492 17460 25498
rect 17512 25480 17540 25774
rect 17604 25498 17632 26182
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 17684 25764 17736 25770
rect 17684 25706 17736 25712
rect 17460 25452 17540 25480
rect 17592 25492 17644 25498
rect 17408 25434 17460 25440
rect 17592 25434 17644 25440
rect 17696 24818 17724 25706
rect 17776 25356 17828 25362
rect 17776 25298 17828 25304
rect 17684 24812 17736 24818
rect 17684 24754 17736 24760
rect 17788 24750 17816 25298
rect 17972 24954 18000 25842
rect 17960 24948 18012 24954
rect 17960 24890 18012 24896
rect 17776 24744 17828 24750
rect 17776 24686 17828 24692
rect 17788 24274 17816 24686
rect 18064 24410 18092 29106
rect 18524 28218 18552 30126
rect 18512 28212 18564 28218
rect 18512 28154 18564 28160
rect 18604 28076 18656 28082
rect 18604 28018 18656 28024
rect 18616 27130 18644 28018
rect 18604 27124 18656 27130
rect 18604 27066 18656 27072
rect 18328 26240 18380 26246
rect 18248 26200 18328 26228
rect 18052 24404 18104 24410
rect 18052 24346 18104 24352
rect 17776 24268 17828 24274
rect 17776 24210 17828 24216
rect 17684 23792 17736 23798
rect 17684 23734 17736 23740
rect 17592 22636 17644 22642
rect 17592 22578 17644 22584
rect 17316 22432 17368 22438
rect 17316 22374 17368 22380
rect 17500 22432 17552 22438
rect 17500 22374 17552 22380
rect 16868 22066 17172 22094
rect 16868 21554 16896 22066
rect 17512 22030 17540 22374
rect 17224 22024 17276 22030
rect 17224 21966 17276 21972
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 16856 21548 16908 21554
rect 16856 21490 16908 21496
rect 17236 20874 17264 21966
rect 17316 21956 17368 21962
rect 17316 21898 17368 21904
rect 17328 21690 17356 21898
rect 17604 21690 17632 22578
rect 17316 21684 17368 21690
rect 17316 21626 17368 21632
rect 17592 21684 17644 21690
rect 17592 21626 17644 21632
rect 17316 21548 17368 21554
rect 17316 21490 17368 21496
rect 17132 20868 17184 20874
rect 17132 20810 17184 20816
rect 17224 20868 17276 20874
rect 17224 20810 17276 20816
rect 17144 20602 17172 20810
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 16578 19000 16634 19009
rect 16578 18935 16634 18944
rect 16592 18834 16620 18935
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16580 18624 16632 18630
rect 16580 18566 16632 18572
rect 16592 18358 16620 18566
rect 16580 18352 16632 18358
rect 16580 18294 16632 18300
rect 16868 18086 16896 18702
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16856 18080 16908 18086
rect 16856 18022 16908 18028
rect 16396 17876 16448 17882
rect 16500 17870 16804 17898
rect 16396 17818 16448 17824
rect 16488 17808 16540 17814
rect 16488 17750 16540 17756
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16224 16782 16344 16810
rect 16120 16516 16172 16522
rect 16120 16458 16172 16464
rect 16028 16176 16080 16182
rect 16028 16118 16080 16124
rect 16040 15434 16068 16118
rect 16028 15428 16080 15434
rect 16028 15370 16080 15376
rect 16040 14890 16068 15370
rect 16028 14884 16080 14890
rect 16028 14826 16080 14832
rect 16028 14272 16080 14278
rect 16028 14214 16080 14220
rect 16040 12306 16068 14214
rect 16132 13938 16160 16458
rect 16224 14482 16252 16782
rect 16408 16726 16436 17682
rect 16396 16720 16448 16726
rect 16396 16662 16448 16668
rect 16500 16658 16528 17750
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16488 16652 16540 16658
rect 16488 16594 16540 16600
rect 16212 14476 16264 14482
rect 16212 14418 16264 14424
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 16316 13870 16344 16594
rect 16684 16522 16712 17070
rect 16776 16590 16804 17870
rect 16960 17134 16988 18566
rect 16948 17128 17000 17134
rect 16948 17070 17000 17076
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16488 16516 16540 16522
rect 16488 16458 16540 16464
rect 16672 16516 16724 16522
rect 16672 16458 16724 16464
rect 16856 16516 16908 16522
rect 16856 16458 16908 16464
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16316 13394 16344 13806
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16028 12300 16080 12306
rect 16028 12242 16080 12248
rect 15936 11892 15988 11898
rect 15936 11834 15988 11840
rect 15844 11280 15896 11286
rect 15844 11222 15896 11228
rect 15856 11150 15884 11222
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15856 10674 15884 11086
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15304 8974 15332 9522
rect 15672 9382 15700 10610
rect 16408 9994 16436 15846
rect 16500 12442 16528 16458
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16592 15366 16620 16050
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16580 14816 16632 14822
rect 16580 14758 16632 14764
rect 16592 14414 16620 14758
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16578 14104 16634 14113
rect 16578 14039 16580 14048
rect 16632 14039 16634 14048
rect 16580 14010 16632 14016
rect 16684 13530 16712 16458
rect 16764 16108 16816 16114
rect 16764 16050 16816 16056
rect 16672 13524 16724 13530
rect 16672 13466 16724 13472
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 16592 13190 16620 13330
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 16592 11150 16620 11766
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16684 11218 16712 11494
rect 16776 11354 16804 16050
rect 16868 15978 16896 16458
rect 16856 15972 16908 15978
rect 16856 15914 16908 15920
rect 16854 15872 16910 15881
rect 16854 15807 16910 15816
rect 16868 14482 16896 15807
rect 16948 15632 17000 15638
rect 16948 15574 17000 15580
rect 16960 15473 16988 15574
rect 16946 15464 17002 15473
rect 16946 15399 17002 15408
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 17052 13938 17080 20402
rect 17132 18828 17184 18834
rect 17132 18770 17184 18776
rect 17144 18698 17172 18770
rect 17132 18692 17184 18698
rect 17132 18634 17184 18640
rect 17236 18222 17264 20810
rect 17328 19530 17356 21490
rect 17408 20800 17460 20806
rect 17408 20742 17460 20748
rect 17420 20466 17448 20742
rect 17408 20460 17460 20466
rect 17408 20402 17460 20408
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 17500 20324 17552 20330
rect 17500 20266 17552 20272
rect 17408 20052 17460 20058
rect 17512 20040 17540 20266
rect 17604 20058 17632 20402
rect 17460 20012 17540 20040
rect 17408 19994 17460 20000
rect 17328 19502 17448 19530
rect 17316 19440 17368 19446
rect 17316 19382 17368 19388
rect 17328 18630 17356 19382
rect 17420 19009 17448 19502
rect 17406 19000 17462 19009
rect 17406 18935 17462 18944
rect 17512 18873 17540 20012
rect 17592 20052 17644 20058
rect 17592 19994 17644 20000
rect 17592 19780 17644 19786
rect 17592 19722 17644 19728
rect 17604 19446 17632 19722
rect 17592 19440 17644 19446
rect 17592 19382 17644 19388
rect 17696 18970 17724 23734
rect 17788 23662 17816 24210
rect 17776 23656 17828 23662
rect 17776 23598 17828 23604
rect 17776 23112 17828 23118
rect 17776 23054 17828 23060
rect 17788 22642 17816 23054
rect 17868 22976 17920 22982
rect 17868 22918 17920 22924
rect 17776 22636 17828 22642
rect 17776 22578 17828 22584
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 17498 18864 17554 18873
rect 17498 18799 17554 18808
rect 17316 18624 17368 18630
rect 17316 18566 17368 18572
rect 17224 18216 17276 18222
rect 17130 18184 17186 18193
rect 17224 18158 17276 18164
rect 17130 18119 17186 18128
rect 17144 17066 17172 18119
rect 17132 17060 17184 17066
rect 17132 17002 17184 17008
rect 17236 16658 17264 18158
rect 17512 17954 17540 18799
rect 17788 18612 17816 22578
rect 17880 22574 17908 22918
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 18156 22148 18184 22510
rect 18248 22506 18276 26200
rect 18328 26182 18380 26188
rect 18788 25832 18840 25838
rect 18788 25774 18840 25780
rect 18420 25220 18472 25226
rect 18420 25162 18472 25168
rect 18432 24682 18460 25162
rect 18800 24818 18828 25774
rect 18788 24812 18840 24818
rect 18788 24754 18840 24760
rect 18420 24676 18472 24682
rect 18420 24618 18472 24624
rect 18328 23860 18380 23866
rect 18432 23848 18460 24618
rect 18512 24404 18564 24410
rect 18512 24346 18564 24352
rect 18696 24404 18748 24410
rect 18696 24346 18748 24352
rect 18380 23820 18460 23848
rect 18328 23802 18380 23808
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 18340 22710 18368 23054
rect 18328 22704 18380 22710
rect 18328 22646 18380 22652
rect 18340 22574 18368 22646
rect 18328 22568 18380 22574
rect 18328 22510 18380 22516
rect 18236 22500 18288 22506
rect 18236 22442 18288 22448
rect 18236 22160 18288 22166
rect 18156 22120 18236 22148
rect 18236 22102 18288 22108
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 18156 19938 18184 20198
rect 18064 19910 18184 19938
rect 17868 19780 17920 19786
rect 17868 19722 17920 19728
rect 17880 19417 17908 19722
rect 17866 19408 17922 19417
rect 17866 19343 17868 19352
rect 17920 19343 17922 19352
rect 17868 19314 17920 19320
rect 17866 19000 17922 19009
rect 17866 18935 17868 18944
rect 17920 18935 17922 18944
rect 17868 18906 17920 18912
rect 17328 17926 17540 17954
rect 17604 18584 17816 18612
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17236 15502 17264 16594
rect 17328 16522 17356 17926
rect 17500 17196 17552 17202
rect 17604 17184 17632 18584
rect 17958 17912 18014 17921
rect 17958 17847 17960 17856
rect 18012 17847 18014 17856
rect 17960 17818 18012 17824
rect 18064 17762 18092 19910
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 18156 19446 18184 19790
rect 18144 19440 18196 19446
rect 18144 19382 18196 19388
rect 18340 19334 18368 22510
rect 18248 19306 18368 19334
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 18156 18766 18184 19110
rect 18144 18760 18196 18766
rect 18144 18702 18196 18708
rect 18248 18086 18276 19306
rect 18328 18760 18380 18766
rect 18326 18728 18328 18737
rect 18380 18728 18382 18737
rect 18326 18663 18382 18672
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 18340 17898 18368 18663
rect 17880 17746 18092 17762
rect 17868 17740 18092 17746
rect 17920 17734 18092 17740
rect 18156 17870 18368 17898
rect 17868 17682 17920 17688
rect 17776 17672 17828 17678
rect 17776 17614 17828 17620
rect 17552 17156 17632 17184
rect 17500 17138 17552 17144
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17420 16590 17448 16934
rect 17408 16584 17460 16590
rect 17408 16526 17460 16532
rect 17316 16516 17368 16522
rect 17316 16458 17368 16464
rect 17604 16454 17632 17156
rect 17684 17196 17736 17202
rect 17684 17138 17736 17144
rect 17500 16448 17552 16454
rect 17500 16390 17552 16396
rect 17592 16448 17644 16454
rect 17592 16390 17644 16396
rect 17512 16114 17540 16390
rect 17696 16266 17724 17138
rect 17788 16998 17816 17614
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 17696 16250 17816 16266
rect 17696 16244 17828 16250
rect 17696 16238 17776 16244
rect 17776 16186 17828 16192
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 17512 16017 17540 16050
rect 17880 16046 17908 17682
rect 17960 17672 18012 17678
rect 17958 17640 17960 17649
rect 18012 17640 18014 17649
rect 17958 17575 18014 17584
rect 18156 17202 18184 17870
rect 18234 17776 18290 17785
rect 18234 17711 18290 17720
rect 18328 17740 18380 17746
rect 18248 17678 18276 17711
rect 18328 17682 18380 17688
rect 18236 17672 18288 17678
rect 18236 17614 18288 17620
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18340 17134 18368 17682
rect 18328 17128 18380 17134
rect 18328 17070 18380 17076
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 17868 16040 17920 16046
rect 17498 16008 17554 16017
rect 17868 15982 17920 15988
rect 17498 15943 17554 15952
rect 17684 15972 17736 15978
rect 17684 15914 17736 15920
rect 17696 15706 17724 15914
rect 17500 15700 17552 15706
rect 17684 15700 17736 15706
rect 17552 15660 17632 15688
rect 17500 15642 17552 15648
rect 17316 15564 17368 15570
rect 17316 15506 17368 15512
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 17224 15020 17276 15026
rect 17328 15008 17356 15506
rect 17408 15156 17460 15162
rect 17460 15116 17540 15144
rect 17408 15098 17460 15104
rect 17276 14980 17356 15008
rect 17224 14962 17276 14968
rect 17222 14920 17278 14929
rect 17222 14855 17224 14864
rect 17276 14855 17278 14864
rect 17224 14826 17276 14832
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 17052 13530 17080 13670
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 16960 12918 16988 13126
rect 16948 12912 17000 12918
rect 16948 12854 17000 12860
rect 16856 12776 16908 12782
rect 16856 12718 16908 12724
rect 16868 11762 16896 12718
rect 16960 12306 16988 12854
rect 17052 12646 17080 13466
rect 17144 13394 17172 14350
rect 17236 14346 17264 14826
rect 17314 14648 17370 14657
rect 17314 14583 17316 14592
rect 17368 14583 17370 14592
rect 17408 14612 17460 14618
rect 17316 14554 17368 14560
rect 17408 14554 17460 14560
rect 17224 14340 17276 14346
rect 17224 14282 17276 14288
rect 17132 13388 17184 13394
rect 17132 13330 17184 13336
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 17144 12306 17172 13330
rect 17236 12918 17264 14282
rect 17420 13852 17448 14554
rect 17512 14006 17540 15116
rect 17500 14000 17552 14006
rect 17500 13942 17552 13948
rect 17500 13864 17552 13870
rect 17420 13824 17500 13852
rect 17500 13806 17552 13812
rect 17512 13734 17540 13806
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17236 12186 17264 12854
rect 17512 12782 17540 13670
rect 17604 13530 17632 15660
rect 17684 15642 17736 15648
rect 17684 15360 17736 15366
rect 17684 15302 17736 15308
rect 17696 15026 17724 15302
rect 17684 15020 17736 15026
rect 17684 14962 17736 14968
rect 17868 14884 17920 14890
rect 17868 14826 17920 14832
rect 17776 14408 17828 14414
rect 17696 14368 17776 14396
rect 17592 13524 17644 13530
rect 17592 13466 17644 13472
rect 17696 12850 17724 14368
rect 17776 14350 17828 14356
rect 17880 14346 17908 14826
rect 17868 14340 17920 14346
rect 17868 14282 17920 14288
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 17880 13462 17908 13670
rect 17868 13456 17920 13462
rect 17868 13398 17920 13404
rect 17972 13258 18000 16390
rect 18432 15162 18460 23820
rect 18524 19854 18552 24346
rect 18708 22438 18736 24346
rect 18800 24206 18828 24754
rect 18788 24200 18840 24206
rect 18788 24142 18840 24148
rect 18800 23866 18828 24142
rect 18788 23860 18840 23866
rect 18788 23802 18840 23808
rect 18604 22432 18656 22438
rect 18604 22374 18656 22380
rect 18696 22432 18748 22438
rect 18696 22374 18748 22380
rect 18616 22098 18644 22374
rect 18604 22092 18656 22098
rect 18604 22034 18656 22040
rect 18708 21622 18736 22374
rect 18696 21616 18748 21622
rect 18696 21558 18748 21564
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18708 20058 18736 20402
rect 18696 20052 18748 20058
rect 18696 19994 18748 20000
rect 18512 19848 18564 19854
rect 18512 19790 18564 19796
rect 18696 19304 18748 19310
rect 18696 19246 18748 19252
rect 18510 18864 18566 18873
rect 18510 18799 18512 18808
rect 18564 18799 18566 18808
rect 18512 18770 18564 18776
rect 18512 18692 18564 18698
rect 18512 18634 18564 18640
rect 18524 16250 18552 18634
rect 18708 18154 18736 19246
rect 18696 18148 18748 18154
rect 18696 18090 18748 18096
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18616 17202 18644 17478
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 18708 15706 18736 18090
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18696 15700 18748 15706
rect 18696 15642 18748 15648
rect 18708 15434 18736 15642
rect 18696 15428 18748 15434
rect 18696 15370 18748 15376
rect 18800 15314 18828 18022
rect 18892 17678 18920 31282
rect 19156 30728 19208 30734
rect 19156 30670 19208 30676
rect 19168 27538 19196 30670
rect 19260 30598 19288 31622
rect 19352 31482 19380 32370
rect 19628 31822 19656 32370
rect 19996 31822 20024 33254
rect 19432 31816 19484 31822
rect 19432 31758 19484 31764
rect 19616 31816 19668 31822
rect 19616 31758 19668 31764
rect 19984 31816 20036 31822
rect 19984 31758 20036 31764
rect 19340 31476 19392 31482
rect 19340 31418 19392 31424
rect 19248 30592 19300 30598
rect 19248 30534 19300 30540
rect 19444 30122 19472 31758
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 20260 31340 20312 31346
rect 20260 31282 20312 31288
rect 20076 30592 20128 30598
rect 20076 30534 20128 30540
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19432 30116 19484 30122
rect 19432 30058 19484 30064
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19248 28620 19300 28626
rect 19248 28562 19300 28568
rect 19260 28014 19288 28562
rect 19984 28484 20036 28490
rect 19984 28426 20036 28432
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19340 28076 19392 28082
rect 19340 28018 19392 28024
rect 19248 28008 19300 28014
rect 19248 27950 19300 27956
rect 19156 27532 19208 27538
rect 19156 27474 19208 27480
rect 18972 27464 19024 27470
rect 18972 27406 19024 27412
rect 18984 26926 19012 27406
rect 19352 27062 19380 28018
rect 19432 27600 19484 27606
rect 19432 27542 19484 27548
rect 19444 27112 19472 27542
rect 19996 27538 20024 28426
rect 20088 27962 20116 30534
rect 20272 30394 20300 31282
rect 20260 30388 20312 30394
rect 20260 30330 20312 30336
rect 20272 29646 20300 30330
rect 20260 29640 20312 29646
rect 20260 29582 20312 29588
rect 20272 29306 20300 29582
rect 20260 29300 20312 29306
rect 20260 29242 20312 29248
rect 20168 28416 20220 28422
rect 20168 28358 20220 28364
rect 20260 28416 20312 28422
rect 20260 28358 20312 28364
rect 20180 28082 20208 28358
rect 20168 28076 20220 28082
rect 20168 28018 20220 28024
rect 20088 27934 20208 27962
rect 20076 27872 20128 27878
rect 20074 27840 20076 27849
rect 20128 27840 20130 27849
rect 20074 27775 20130 27784
rect 20076 27668 20128 27674
rect 20076 27610 20128 27616
rect 19984 27532 20036 27538
rect 19984 27474 20036 27480
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19444 27084 19564 27112
rect 19340 27056 19392 27062
rect 19340 26998 19392 27004
rect 18972 26920 19024 26926
rect 18972 26862 19024 26868
rect 19352 26586 19380 26998
rect 19432 26852 19484 26858
rect 19432 26794 19484 26800
rect 19340 26580 19392 26586
rect 19340 26522 19392 26528
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 19340 26376 19392 26382
rect 19340 26318 19392 26324
rect 19260 25498 19288 26318
rect 19352 25786 19380 26318
rect 19444 26296 19472 26794
rect 19536 26790 19564 27084
rect 19996 26994 20024 27474
rect 20088 27130 20116 27610
rect 20076 27124 20128 27130
rect 20076 27066 20128 27072
rect 19984 26988 20036 26994
rect 19984 26930 20036 26936
rect 19524 26784 19576 26790
rect 19524 26726 19576 26732
rect 19984 26784 20036 26790
rect 19984 26726 20036 26732
rect 19524 26308 19576 26314
rect 19444 26268 19524 26296
rect 19444 25906 19472 26268
rect 19524 26250 19576 26256
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19432 25900 19484 25906
rect 19432 25842 19484 25848
rect 19352 25758 19472 25786
rect 19340 25696 19392 25702
rect 19340 25638 19392 25644
rect 19248 25492 19300 25498
rect 19248 25434 19300 25440
rect 18972 25152 19024 25158
rect 18972 25094 19024 25100
rect 18984 24818 19012 25094
rect 18972 24812 19024 24818
rect 18972 24754 19024 24760
rect 19260 24410 19288 25434
rect 19352 25226 19380 25638
rect 19340 25220 19392 25226
rect 19340 25162 19392 25168
rect 19444 24750 19472 25758
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19432 24744 19484 24750
rect 19432 24686 19484 24692
rect 19248 24404 19300 24410
rect 19248 24346 19300 24352
rect 19444 24138 19472 24686
rect 19432 24132 19484 24138
rect 19432 24074 19484 24080
rect 19996 24070 20024 26726
rect 20076 25220 20128 25226
rect 20076 25162 20128 25168
rect 20088 24274 20116 25162
rect 20076 24268 20128 24274
rect 20076 24210 20128 24216
rect 19984 24064 20036 24070
rect 19984 24006 20036 24012
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 20088 23322 20116 24210
rect 20076 23316 20128 23322
rect 20076 23258 20128 23264
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19432 22432 19484 22438
rect 19432 22374 19484 22380
rect 19444 21672 19472 22374
rect 20180 22094 20208 27934
rect 20272 26586 20300 28358
rect 20260 26580 20312 26586
rect 20260 26522 20312 26528
rect 20260 26240 20312 26246
rect 20260 26182 20312 26188
rect 20088 22066 20208 22094
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19260 21644 19472 21672
rect 19260 20516 19288 21644
rect 19340 21548 19392 21554
rect 19340 21490 19392 21496
rect 19352 21146 19380 21490
rect 19984 21344 20036 21350
rect 19984 21286 20036 21292
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19340 21004 19392 21010
rect 19340 20946 19392 20952
rect 19168 20488 19288 20516
rect 19168 20398 19196 20488
rect 19156 20392 19208 20398
rect 19156 20334 19208 20340
rect 19248 20256 19300 20262
rect 19352 20244 19380 20946
rect 19996 20942 20024 21286
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19984 20936 20036 20942
rect 19984 20878 20036 20884
rect 19300 20216 19380 20244
rect 19248 20198 19300 20204
rect 19444 20058 19472 20878
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19996 20534 20024 20878
rect 19984 20528 20036 20534
rect 19984 20470 20036 20476
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 18972 19984 19024 19990
rect 18972 19926 19024 19932
rect 19616 19984 19668 19990
rect 19616 19926 19668 19932
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 18708 15286 18828 15314
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 18604 15020 18656 15026
rect 18604 14962 18656 14968
rect 18156 14006 18184 14962
rect 18144 14000 18196 14006
rect 18144 13942 18196 13948
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 18064 13326 18092 13874
rect 18156 13734 18184 13942
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 18156 13258 18184 13670
rect 17960 13252 18012 13258
rect 17960 13194 18012 13200
rect 18144 13252 18196 13258
rect 18144 13194 18196 13200
rect 18052 13184 18104 13190
rect 18248 13138 18276 14962
rect 18616 14929 18644 14962
rect 18602 14920 18658 14929
rect 18602 14855 18658 14864
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18420 13864 18472 13870
rect 18420 13806 18472 13812
rect 18432 13734 18460 13806
rect 18420 13728 18472 13734
rect 18420 13670 18472 13676
rect 18524 13530 18552 14214
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18052 13126 18104 13132
rect 17684 12844 17736 12850
rect 17684 12786 17736 12792
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17512 12238 17540 12718
rect 17144 12158 17264 12186
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16764 11348 16816 11354
rect 16764 11290 16816 11296
rect 16672 11212 16724 11218
rect 16672 11154 16724 11160
rect 16868 11150 16896 11698
rect 17144 11218 17172 12158
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17144 10674 17172 10950
rect 17132 10668 17184 10674
rect 16960 10628 17132 10656
rect 16396 9988 16448 9994
rect 16396 9930 16448 9936
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 16212 9104 16264 9110
rect 16212 9046 16264 9052
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15200 8356 15252 8362
rect 15200 8298 15252 8304
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 15120 7546 15148 7822
rect 15476 7812 15528 7818
rect 15476 7754 15528 7760
rect 15488 7546 15516 7754
rect 16040 7750 16068 8230
rect 16132 8090 16160 8230
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 14924 7268 14976 7274
rect 14924 7210 14976 7216
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 14556 6724 14608 6730
rect 14556 6666 14608 6672
rect 14740 6724 14792 6730
rect 14740 6666 14792 6672
rect 14752 6322 14780 6666
rect 15212 6662 15240 6802
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 15120 6458 15148 6598
rect 15108 6452 15160 6458
rect 15108 6394 15160 6400
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 14384 4984 14596 5012
rect 14280 4966 14332 4972
rect 14370 4720 14426 4729
rect 14370 4655 14426 4664
rect 14280 4548 14332 4554
rect 14280 4490 14332 4496
rect 14292 4146 14320 4490
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14292 3534 14320 4082
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14108 2746 14228 2774
rect 14004 2032 14056 2038
rect 14004 1974 14056 1980
rect 14108 1442 14136 2746
rect 14016 1414 14136 1442
rect 14016 800 14044 1414
rect 14384 800 14412 4655
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14476 3602 14504 4558
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14568 2854 14596 4984
rect 14660 4826 14688 5170
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14752 4690 14780 6258
rect 15028 6225 15056 6258
rect 15014 6216 15070 6225
rect 15014 6151 15070 6160
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15120 5574 15148 5714
rect 15212 5642 15240 6598
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 15304 5914 15332 6326
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 15200 5636 15252 5642
rect 15200 5578 15252 5584
rect 15108 5568 15160 5574
rect 15108 5510 15160 5516
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 14660 2990 14688 4558
rect 14752 4214 14780 4626
rect 14740 4208 14792 4214
rect 14740 4150 14792 4156
rect 14752 3942 14780 4150
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14752 3602 14780 3878
rect 14740 3596 14792 3602
rect 14740 3538 14792 3544
rect 14740 3120 14792 3126
rect 14740 3062 14792 3068
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 14752 800 14780 3062
rect 14844 2514 14872 4082
rect 15016 3732 15068 3738
rect 15016 3674 15068 3680
rect 15028 2774 15056 3674
rect 15120 3482 15148 5306
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15212 4026 15240 4966
rect 15304 4146 15332 5714
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15212 3998 15332 4026
rect 15120 3466 15240 3482
rect 15120 3460 15252 3466
rect 15120 3454 15200 3460
rect 15200 3402 15252 3408
rect 15304 3126 15332 3998
rect 15396 3369 15424 4966
rect 15580 4282 15608 5170
rect 15568 4276 15620 4282
rect 15568 4218 15620 4224
rect 15672 4162 15700 7142
rect 15764 5914 15792 7346
rect 16040 7002 16068 7346
rect 16120 7336 16172 7342
rect 16120 7278 16172 7284
rect 16028 6996 16080 7002
rect 16028 6938 16080 6944
rect 16132 6798 16160 7278
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15948 5681 15976 6598
rect 16132 6254 16160 6734
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 16132 5914 16160 6054
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 15934 5672 15990 5681
rect 15934 5607 15990 5616
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15580 4134 15700 4162
rect 15752 4140 15804 4146
rect 15488 3738 15516 4082
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15580 3618 15608 4134
rect 15752 4082 15804 4088
rect 15660 4004 15712 4010
rect 15660 3946 15712 3952
rect 15488 3590 15608 3618
rect 15382 3360 15438 3369
rect 15382 3295 15438 3304
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 15028 2746 15148 2774
rect 14832 2508 14884 2514
rect 14832 2450 14884 2456
rect 15120 800 15148 2746
rect 15488 800 15516 3590
rect 15568 3120 15620 3126
rect 15568 3062 15620 3068
rect 5828 734 6132 762
rect 6182 0 6238 800
rect 6550 0 6606 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8390 0 8446 800
rect 8758 0 8814 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9862 0 9918 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15580 762 15608 3062
rect 15672 2972 15700 3946
rect 15764 3194 15792 4082
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 15752 2984 15804 2990
rect 15672 2944 15752 2972
rect 15752 2926 15804 2932
rect 15764 2446 15792 2926
rect 15856 2650 15884 5170
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 15948 3398 15976 4082
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 16040 2378 16068 3470
rect 16132 3058 16160 3878
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 15660 2372 15712 2378
rect 15660 2314 15712 2320
rect 16028 2372 16080 2378
rect 16028 2314 16080 2320
rect 15672 1630 15700 2314
rect 15660 1624 15712 1630
rect 15660 1566 15712 1572
rect 15764 870 15884 898
rect 15764 762 15792 870
rect 15856 800 15884 870
rect 16224 800 16252 9046
rect 16408 8906 16436 9522
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16684 9042 16712 9454
rect 16960 9450 16988 10628
rect 17132 10610 17184 10616
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 16948 9444 17000 9450
rect 16948 9386 17000 9392
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16396 8900 16448 8906
rect 16396 8842 16448 8848
rect 16592 8634 16620 8910
rect 16672 8900 16724 8906
rect 16672 8842 16724 8848
rect 16684 8634 16712 8842
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16396 8356 16448 8362
rect 16396 8298 16448 8304
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16316 7002 16344 7890
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 16316 5642 16344 6598
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 16304 2984 16356 2990
rect 16408 2972 16436 8298
rect 16592 8090 16620 8434
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16488 8016 16540 8022
rect 16684 7970 16712 8570
rect 16540 7964 16712 7970
rect 16488 7958 16712 7964
rect 16500 7942 16712 7958
rect 16960 7886 16988 9386
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16592 7410 16620 7686
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 16500 6458 16528 6734
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 16592 5914 16620 7346
rect 17052 7290 17080 10202
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 17144 8974 17172 10066
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17144 8498 17172 8910
rect 17236 8498 17264 11290
rect 17696 11218 17724 12786
rect 18064 11354 18092 13126
rect 18156 13110 18276 13138
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 17316 11212 17368 11218
rect 17316 11154 17368 11160
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17328 9110 17356 11154
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17880 10606 17908 11018
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 18156 10538 18184 13110
rect 18708 12918 18736 15286
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18788 14544 18840 14550
rect 18788 14486 18840 14492
rect 18696 12912 18748 12918
rect 18696 12854 18748 12860
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18248 12442 18276 12786
rect 18236 12436 18288 12442
rect 18236 12378 18288 12384
rect 18248 11064 18276 12378
rect 18524 11898 18552 12786
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18420 11076 18472 11082
rect 18248 11036 18420 11064
rect 18420 11018 18472 11024
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 18144 10532 18196 10538
rect 18144 10474 18196 10480
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17776 10056 17828 10062
rect 17880 10044 17908 10406
rect 18524 10266 18552 10610
rect 18604 10464 18656 10470
rect 18604 10406 18656 10412
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 17828 10016 17908 10044
rect 17776 9998 17828 10004
rect 17684 9648 17736 9654
rect 17684 9590 17736 9596
rect 17498 9480 17554 9489
rect 17498 9415 17554 9424
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17144 7410 17172 8434
rect 17512 8090 17540 9415
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17604 8906 17632 9318
rect 17696 8906 17724 9590
rect 17880 8974 17908 10016
rect 18616 9994 18644 10406
rect 18604 9988 18656 9994
rect 18604 9930 18656 9936
rect 18694 9752 18750 9761
rect 18694 9687 18750 9696
rect 17960 9580 18012 9586
rect 18236 9580 18288 9586
rect 18012 9540 18092 9568
rect 17960 9522 18012 9528
rect 17960 9444 18012 9450
rect 17960 9386 18012 9392
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17592 8900 17644 8906
rect 17592 8842 17644 8848
rect 17684 8900 17736 8906
rect 17684 8842 17736 8848
rect 17880 8498 17908 8910
rect 17972 8838 18000 9386
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17500 8084 17552 8090
rect 17552 8044 17632 8072
rect 17500 8026 17552 8032
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 17420 7342 17448 7686
rect 17408 7336 17460 7342
rect 17052 7262 17356 7290
rect 17408 7278 17460 7284
rect 16672 6996 16724 7002
rect 16672 6938 16724 6944
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16684 5778 16712 6938
rect 17222 6488 17278 6497
rect 17222 6423 17278 6432
rect 17236 6322 17264 6423
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 17130 5944 17186 5953
rect 17130 5879 17186 5888
rect 17144 5846 17172 5879
rect 17132 5840 17184 5846
rect 17132 5782 17184 5788
rect 16672 5772 16724 5778
rect 16672 5714 16724 5720
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16500 4486 16528 5646
rect 16948 5568 17000 5574
rect 16948 5510 17000 5516
rect 16960 5302 16988 5510
rect 16948 5296 17000 5302
rect 16948 5238 17000 5244
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 16580 4548 16632 4554
rect 16580 4490 16632 4496
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 16356 2944 16436 2972
rect 16304 2926 16356 2932
rect 16316 2582 16344 2926
rect 16304 2576 16356 2582
rect 16304 2518 16356 2524
rect 16500 2310 16528 4422
rect 16592 3194 16620 4490
rect 17040 4072 17092 4078
rect 17040 4014 17092 4020
rect 17052 3602 17080 4014
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 16672 2848 16724 2854
rect 16724 2796 16804 2802
rect 16672 2790 16804 2796
rect 16684 2774 16804 2790
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 16592 800 16620 2586
rect 16776 2446 16804 2774
rect 16960 2446 16988 2926
rect 17144 2446 17172 4626
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 17040 2372 17092 2378
rect 17040 2314 17092 2320
rect 17052 1834 17080 2314
rect 17040 1828 17092 1834
rect 17040 1770 17092 1776
rect 16960 870 17080 898
rect 16960 800 16988 870
rect 15580 734 15792 762
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17052 762 17080 870
rect 17328 762 17356 7262
rect 17420 5234 17448 7278
rect 17512 5370 17540 7890
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17604 4622 17632 8044
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 17696 5710 17724 6190
rect 17788 5953 17816 8366
rect 17880 6798 17908 8434
rect 17972 7818 18000 8774
rect 18064 7886 18092 9540
rect 18236 9522 18288 9528
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 18156 8090 18184 8434
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18248 7886 18276 9522
rect 18616 8634 18644 9522
rect 18708 9450 18736 9687
rect 18800 9586 18828 14486
rect 18892 12850 18920 14826
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18984 12434 19012 19926
rect 19628 19854 19656 19926
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19616 19848 19668 19854
rect 19720 19825 19748 19858
rect 19616 19790 19668 19796
rect 19706 19816 19762 19825
rect 19352 19378 19380 19790
rect 19706 19751 19762 19760
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19444 19417 19472 19654
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19430 19408 19486 19417
rect 19340 19372 19392 19378
rect 19430 19343 19486 19352
rect 19340 19314 19392 19320
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 19064 19168 19116 19174
rect 19064 19110 19116 19116
rect 19076 18358 19104 19110
rect 19168 18766 19196 19246
rect 19156 18760 19208 18766
rect 19156 18702 19208 18708
rect 19064 18352 19116 18358
rect 19064 18294 19116 18300
rect 19352 17954 19380 19314
rect 19996 18834 20024 20470
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 19432 18692 19484 18698
rect 19432 18634 19484 18640
rect 19444 18034 19472 18634
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19892 18284 19944 18290
rect 19996 18272 20024 18770
rect 19944 18244 20024 18272
rect 19892 18226 19944 18232
rect 19444 18006 19840 18034
rect 19352 17926 19472 17954
rect 19444 17814 19472 17926
rect 19432 17808 19484 17814
rect 19154 17776 19210 17785
rect 19432 17750 19484 17756
rect 19524 17808 19576 17814
rect 19524 17750 19576 17756
rect 19154 17711 19210 17720
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 19076 12714 19104 15438
rect 19064 12708 19116 12714
rect 19064 12650 19116 12656
rect 18892 12406 19012 12434
rect 18788 9580 18840 9586
rect 18788 9522 18840 9528
rect 18696 9444 18748 9450
rect 18696 9386 18748 9392
rect 18708 9178 18736 9386
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18892 8480 18920 12406
rect 18972 12164 19024 12170
rect 18972 12106 19024 12112
rect 18984 9382 19012 12106
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 18800 8452 18920 8480
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 17960 7812 18012 7818
rect 17960 7754 18012 7760
rect 18248 7546 18276 7822
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18052 6928 18104 6934
rect 18052 6870 18104 6876
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17774 5944 17830 5953
rect 18064 5914 18092 6870
rect 17774 5879 17830 5888
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 18432 5710 18460 5850
rect 18616 5778 18644 7482
rect 18800 6934 18828 8452
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 18880 8356 18932 8362
rect 18880 8298 18932 8304
rect 18788 6928 18840 6934
rect 18788 6870 18840 6876
rect 18892 6390 18920 8298
rect 18880 6384 18932 6390
rect 18880 6326 18932 6332
rect 18604 5772 18656 5778
rect 18604 5714 18656 5720
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 18420 5704 18472 5710
rect 18420 5646 18472 5652
rect 18616 5574 18644 5714
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18604 5568 18656 5574
rect 18604 5510 18656 5516
rect 18156 5302 18184 5510
rect 18984 5370 19012 8366
rect 19076 6798 19104 12650
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 18972 5364 19024 5370
rect 18972 5306 19024 5312
rect 18144 5296 18196 5302
rect 17774 5264 17830 5273
rect 18144 5238 18196 5244
rect 17774 5199 17830 5208
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17408 2576 17460 2582
rect 17408 2518 17460 2524
rect 17420 800 17448 2518
rect 17592 2508 17644 2514
rect 17592 2450 17644 2456
rect 17604 2378 17632 2450
rect 17592 2372 17644 2378
rect 17592 2314 17644 2320
rect 17788 800 17816 5199
rect 18604 5092 18656 5098
rect 18604 5034 18656 5040
rect 18510 4856 18566 4865
rect 18616 4826 18644 5034
rect 18510 4791 18566 4800
rect 18604 4820 18656 4826
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 18144 4480 18196 4486
rect 18144 4422 18196 4428
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 17972 3097 18000 3674
rect 17958 3088 18014 3097
rect 17958 3023 17960 3032
rect 18012 3023 18014 3032
rect 17960 2994 18012 3000
rect 18064 2854 18092 3878
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 17868 2440 17920 2446
rect 18052 2440 18104 2446
rect 17920 2400 18052 2428
rect 17868 2382 17920 2388
rect 18052 2382 18104 2388
rect 18156 800 18184 4422
rect 18328 4276 18380 4282
rect 18328 4218 18380 4224
rect 18236 3120 18288 3126
rect 18234 3088 18236 3097
rect 18288 3088 18290 3097
rect 18340 3058 18368 4218
rect 18432 3194 18460 4558
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 18234 3023 18290 3032
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 18340 2514 18368 2994
rect 18328 2508 18380 2514
rect 18328 2450 18380 2456
rect 18524 800 18552 4791
rect 18604 4762 18656 4768
rect 18880 3664 18932 3670
rect 18880 3606 18932 3612
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18616 2446 18644 3334
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 18892 800 18920 3606
rect 19076 2774 19104 6734
rect 19168 6186 19196 17711
rect 19260 17678 19288 17709
rect 19248 17672 19300 17678
rect 19246 17640 19248 17649
rect 19300 17640 19302 17649
rect 19536 17626 19564 17750
rect 19708 17672 19760 17678
rect 19302 17598 19564 17626
rect 19706 17640 19708 17649
rect 19760 17640 19762 17649
rect 19246 17575 19302 17584
rect 19706 17575 19762 17584
rect 19248 17536 19300 17542
rect 19248 17478 19300 17484
rect 19340 17536 19392 17542
rect 19812 17524 19840 18006
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 19340 17478 19392 17484
rect 19444 17496 19840 17524
rect 19260 16114 19288 17478
rect 19352 16590 19380 17478
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19340 16176 19392 16182
rect 19340 16118 19392 16124
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19248 14952 19300 14958
rect 19246 14920 19248 14929
rect 19300 14920 19302 14929
rect 19246 14855 19302 14864
rect 19248 14816 19300 14822
rect 19248 14758 19300 14764
rect 19260 13938 19288 14758
rect 19352 14113 19380 16118
rect 19338 14104 19394 14113
rect 19338 14039 19394 14048
rect 19248 13932 19300 13938
rect 19248 13874 19300 13880
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19352 13258 19380 13806
rect 19248 13252 19300 13258
rect 19248 13194 19300 13200
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19260 13161 19288 13194
rect 19246 13152 19302 13161
rect 19246 13087 19302 13096
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 19352 10010 19380 12038
rect 19444 10742 19472 17496
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19798 17232 19854 17241
rect 19616 17196 19668 17202
rect 19798 17167 19854 17176
rect 19616 17138 19668 17144
rect 19628 17105 19656 17138
rect 19614 17096 19670 17105
rect 19614 17031 19670 17040
rect 19706 16960 19762 16969
rect 19706 16895 19762 16904
rect 19720 16794 19748 16895
rect 19708 16788 19760 16794
rect 19708 16730 19760 16736
rect 19812 16522 19840 17167
rect 19996 17134 20024 17682
rect 20088 17649 20116 22066
rect 20168 22024 20220 22030
rect 20168 21966 20220 21972
rect 20180 19174 20208 21966
rect 20272 19990 20300 26182
rect 20364 22030 20392 46990
rect 28092 46374 28120 46990
rect 36268 46912 36320 46918
rect 36268 46854 36320 46860
rect 28080 46368 28132 46374
rect 28080 46310 28132 46316
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 22008 34604 22060 34610
rect 22008 34546 22060 34552
rect 21824 34400 21876 34406
rect 21824 34342 21876 34348
rect 21180 33992 21232 33998
rect 21180 33934 21232 33940
rect 20812 33516 20864 33522
rect 20812 33458 20864 33464
rect 21088 33516 21140 33522
rect 21088 33458 21140 33464
rect 20824 33114 20852 33458
rect 20812 33108 20864 33114
rect 20812 33050 20864 33056
rect 20628 32768 20680 32774
rect 20628 32710 20680 32716
rect 20996 32768 21048 32774
rect 20996 32710 21048 32716
rect 20536 32496 20588 32502
rect 20536 32438 20588 32444
rect 20444 31816 20496 31822
rect 20444 31758 20496 31764
rect 20456 30326 20484 31758
rect 20444 30320 20496 30326
rect 20444 30262 20496 30268
rect 20456 29594 20484 30262
rect 20548 29850 20576 32438
rect 20640 32366 20668 32710
rect 21008 32434 21036 32710
rect 21100 32570 21128 33458
rect 21192 33454 21220 33934
rect 21180 33448 21232 33454
rect 21180 33390 21232 33396
rect 21192 32910 21220 33390
rect 21836 32910 21864 34342
rect 21916 33856 21968 33862
rect 21916 33798 21968 33804
rect 21180 32904 21232 32910
rect 21180 32846 21232 32852
rect 21824 32904 21876 32910
rect 21824 32846 21876 32852
rect 21088 32564 21140 32570
rect 21088 32506 21140 32512
rect 20720 32428 20772 32434
rect 20720 32370 20772 32376
rect 20996 32428 21048 32434
rect 20996 32370 21048 32376
rect 20628 32360 20680 32366
rect 20628 32302 20680 32308
rect 20640 31346 20668 32302
rect 20732 31890 20760 32370
rect 20720 31884 20772 31890
rect 20720 31826 20772 31832
rect 20628 31340 20680 31346
rect 20628 31282 20680 31288
rect 20640 30598 20668 31282
rect 20720 31272 20772 31278
rect 20720 31214 20772 31220
rect 20904 31272 20956 31278
rect 20904 31214 20956 31220
rect 20628 30592 20680 30598
rect 20628 30534 20680 30540
rect 20536 29844 20588 29850
rect 20536 29786 20588 29792
rect 20628 29708 20680 29714
rect 20628 29650 20680 29656
rect 20456 29566 20576 29594
rect 20444 29504 20496 29510
rect 20444 29446 20496 29452
rect 20456 26246 20484 29446
rect 20444 26240 20496 26246
rect 20444 26182 20496 26188
rect 20444 25696 20496 25702
rect 20444 25638 20496 25644
rect 20456 25226 20484 25638
rect 20444 25220 20496 25226
rect 20444 25162 20496 25168
rect 20548 22094 20576 29566
rect 20640 28218 20668 29650
rect 20732 28762 20760 31214
rect 20916 29306 20944 31214
rect 21008 29832 21036 32370
rect 21088 31748 21140 31754
rect 21088 31690 21140 31696
rect 21100 31482 21128 31690
rect 21088 31476 21140 31482
rect 21088 31418 21140 31424
rect 21008 29804 21128 29832
rect 20996 29708 21048 29714
rect 20996 29650 21048 29656
rect 20904 29300 20956 29306
rect 20904 29242 20956 29248
rect 20904 29164 20956 29170
rect 20904 29106 20956 29112
rect 20810 29064 20866 29073
rect 20810 28999 20866 29008
rect 20720 28756 20772 28762
rect 20720 28698 20772 28704
rect 20824 28694 20852 28999
rect 20812 28688 20864 28694
rect 20812 28630 20864 28636
rect 20628 28212 20680 28218
rect 20628 28154 20680 28160
rect 20628 28008 20680 28014
rect 20628 27950 20680 27956
rect 20640 27402 20668 27950
rect 20720 27872 20772 27878
rect 20720 27814 20772 27820
rect 20732 27470 20760 27814
rect 20720 27464 20772 27470
rect 20720 27406 20772 27412
rect 20628 27396 20680 27402
rect 20628 27338 20680 27344
rect 20640 26858 20668 27338
rect 20628 26852 20680 26858
rect 20628 26794 20680 26800
rect 20732 26466 20760 27406
rect 20916 26586 20944 29106
rect 21008 27606 21036 29650
rect 21100 29510 21128 29804
rect 21088 29504 21140 29510
rect 21088 29446 21140 29452
rect 21088 28484 21140 28490
rect 21088 28426 21140 28432
rect 21100 28082 21128 28426
rect 21088 28076 21140 28082
rect 21088 28018 21140 28024
rect 21100 27878 21128 28018
rect 21088 27872 21140 27878
rect 21088 27814 21140 27820
rect 21100 27606 21128 27814
rect 20996 27600 21048 27606
rect 20996 27542 21048 27548
rect 21088 27600 21140 27606
rect 21088 27542 21140 27548
rect 21088 27464 21140 27470
rect 21088 27406 21140 27412
rect 20812 26580 20864 26586
rect 20812 26522 20864 26528
rect 20904 26580 20956 26586
rect 20904 26522 20956 26528
rect 20640 26438 20760 26466
rect 20640 25838 20668 26438
rect 20720 26376 20772 26382
rect 20720 26318 20772 26324
rect 20628 25832 20680 25838
rect 20628 25774 20680 25780
rect 20732 25294 20760 26318
rect 20824 25906 20852 26522
rect 20916 26246 20944 26522
rect 20996 26444 21048 26450
rect 20996 26386 21048 26392
rect 20904 26240 20956 26246
rect 20904 26182 20956 26188
rect 21008 26042 21036 26386
rect 21100 26382 21128 27406
rect 21088 26376 21140 26382
rect 21088 26318 21140 26324
rect 20996 26036 21048 26042
rect 20996 25978 21048 25984
rect 20812 25900 20864 25906
rect 20812 25842 20864 25848
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20824 25158 20852 25842
rect 21008 25362 21036 25978
rect 20996 25356 21048 25362
rect 20996 25298 21048 25304
rect 20904 25288 20956 25294
rect 20904 25230 20956 25236
rect 20812 25152 20864 25158
rect 20812 25094 20864 25100
rect 20916 24818 20944 25230
rect 20904 24812 20956 24818
rect 20904 24754 20956 24760
rect 21100 24410 21128 26318
rect 21088 24404 21140 24410
rect 21088 24346 21140 24352
rect 20628 24064 20680 24070
rect 20628 24006 20680 24012
rect 20456 22066 20576 22094
rect 20352 22024 20404 22030
rect 20352 21966 20404 21972
rect 20260 19984 20312 19990
rect 20260 19926 20312 19932
rect 20456 19836 20484 22066
rect 20536 21344 20588 21350
rect 20536 21286 20588 21292
rect 20548 20806 20576 21286
rect 20536 20800 20588 20806
rect 20536 20742 20588 20748
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20548 20058 20576 20198
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20640 19938 20668 24006
rect 21192 23866 21220 32846
rect 21456 32836 21508 32842
rect 21456 32778 21508 32784
rect 21468 32026 21496 32778
rect 21456 32020 21508 32026
rect 21456 31962 21508 31968
rect 21928 31770 21956 33798
rect 22020 33658 22048 34546
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 22468 33992 22520 33998
rect 22468 33934 22520 33940
rect 22652 33992 22704 33998
rect 22652 33934 22704 33940
rect 22008 33652 22060 33658
rect 22008 33594 22060 33600
rect 22480 33590 22508 33934
rect 22468 33584 22520 33590
rect 22468 33526 22520 33532
rect 22376 33312 22428 33318
rect 22376 33254 22428 33260
rect 22388 32502 22416 33254
rect 22480 32978 22508 33526
rect 22468 32972 22520 32978
rect 22468 32914 22520 32920
rect 22664 32570 22692 33934
rect 23296 33856 23348 33862
rect 23296 33798 23348 33804
rect 23308 33590 23336 33798
rect 23296 33584 23348 33590
rect 23296 33526 23348 33532
rect 24400 33516 24452 33522
rect 24400 33458 24452 33464
rect 24216 33312 24268 33318
rect 24216 33254 24268 33260
rect 22652 32564 22704 32570
rect 22652 32506 22704 32512
rect 24228 32502 24256 33254
rect 24412 33114 24440 33458
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 24400 33108 24452 33114
rect 24400 33050 24452 33056
rect 24768 32972 24820 32978
rect 24768 32914 24820 32920
rect 24584 32904 24636 32910
rect 24584 32846 24636 32852
rect 22376 32496 22428 32502
rect 22376 32438 22428 32444
rect 24216 32496 24268 32502
rect 24216 32438 24268 32444
rect 22008 32428 22060 32434
rect 22008 32370 22060 32376
rect 22284 32428 22336 32434
rect 22284 32370 22336 32376
rect 22020 31890 22048 32370
rect 22296 32026 22324 32370
rect 22284 32020 22336 32026
rect 22284 31962 22336 31968
rect 22008 31884 22060 31890
rect 22008 31826 22060 31832
rect 21548 31748 21600 31754
rect 21548 31690 21600 31696
rect 21836 31742 21956 31770
rect 22020 31754 22048 31826
rect 22388 31754 22416 32438
rect 22560 32428 22612 32434
rect 22560 32370 22612 32376
rect 23480 32428 23532 32434
rect 23480 32370 23532 32376
rect 22468 31884 22520 31890
rect 22468 31826 22520 31832
rect 22008 31748 22060 31754
rect 21560 30802 21588 31690
rect 21836 31686 21864 31742
rect 22008 31690 22060 31696
rect 22296 31726 22416 31754
rect 22296 31686 22324 31726
rect 21824 31680 21876 31686
rect 21824 31622 21876 31628
rect 22284 31680 22336 31686
rect 22284 31622 22336 31628
rect 22376 31680 22428 31686
rect 22376 31622 22428 31628
rect 21836 31346 21864 31622
rect 21824 31340 21876 31346
rect 21824 31282 21876 31288
rect 21548 30796 21600 30802
rect 21548 30738 21600 30744
rect 21640 29504 21692 29510
rect 21640 29446 21692 29452
rect 21456 28620 21508 28626
rect 21456 28562 21508 28568
rect 21468 28422 21496 28562
rect 21456 28416 21508 28422
rect 21456 28358 21508 28364
rect 21272 28076 21324 28082
rect 21272 28018 21324 28024
rect 21284 27470 21312 28018
rect 21272 27464 21324 27470
rect 21272 27406 21324 27412
rect 21548 26376 21600 26382
rect 21548 26318 21600 26324
rect 21456 25832 21508 25838
rect 21456 25774 21508 25780
rect 21272 25764 21324 25770
rect 21272 25706 21324 25712
rect 21284 24886 21312 25706
rect 21364 25288 21416 25294
rect 21364 25230 21416 25236
rect 21272 24880 21324 24886
rect 21272 24822 21324 24828
rect 21284 24410 21312 24822
rect 21272 24404 21324 24410
rect 21272 24346 21324 24352
rect 21376 23866 21404 25230
rect 21468 24818 21496 25774
rect 21456 24812 21508 24818
rect 21456 24754 21508 24760
rect 21560 24614 21588 26318
rect 21548 24608 21600 24614
rect 21548 24550 21600 24556
rect 21560 24154 21588 24550
rect 21468 24126 21588 24154
rect 21468 24070 21496 24126
rect 21456 24064 21508 24070
rect 21456 24006 21508 24012
rect 21180 23860 21232 23866
rect 21180 23802 21232 23808
rect 21364 23860 21416 23866
rect 21364 23802 21416 23808
rect 21192 23118 21220 23802
rect 21548 23724 21600 23730
rect 21548 23666 21600 23672
rect 21180 23112 21232 23118
rect 21180 23054 21232 23060
rect 20720 23044 20772 23050
rect 20720 22986 20772 22992
rect 21088 23044 21140 23050
rect 21088 22986 21140 22992
rect 20732 22166 20760 22986
rect 20904 22500 20956 22506
rect 20904 22442 20956 22448
rect 20720 22160 20772 22166
rect 20720 22102 20772 22108
rect 20812 22024 20864 22030
rect 20812 21966 20864 21972
rect 20824 21690 20852 21966
rect 20812 21684 20864 21690
rect 20812 21626 20864 21632
rect 20812 20936 20864 20942
rect 20812 20878 20864 20884
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20364 19808 20484 19836
rect 20548 19910 20668 19938
rect 20260 19712 20312 19718
rect 20260 19654 20312 19660
rect 20168 19168 20220 19174
rect 20168 19110 20220 19116
rect 20168 17808 20220 17814
rect 20168 17750 20220 17756
rect 20074 17640 20130 17649
rect 20074 17575 20130 17584
rect 20076 17196 20128 17202
rect 20180 17184 20208 17750
rect 20272 17746 20300 19654
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 20364 17678 20392 19808
rect 20444 19712 20496 19718
rect 20444 19654 20496 19660
rect 20456 18358 20484 19654
rect 20548 18902 20576 19910
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20536 18896 20588 18902
rect 20536 18838 20588 18844
rect 20444 18352 20496 18358
rect 20444 18294 20496 18300
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20456 17678 20484 18022
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20444 17672 20496 17678
rect 20444 17614 20496 17620
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20364 17202 20392 17478
rect 20128 17156 20208 17184
rect 20352 17196 20404 17202
rect 20076 17138 20128 17144
rect 20352 17138 20404 17144
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 20352 16992 20404 16998
rect 20456 16969 20484 17070
rect 20352 16934 20404 16940
rect 20442 16960 20498 16969
rect 19800 16516 19852 16522
rect 19800 16458 19852 16464
rect 20364 16454 20392 16934
rect 20442 16895 20498 16904
rect 20352 16448 20404 16454
rect 20352 16390 20404 16396
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 19892 16108 19944 16114
rect 20168 16108 20220 16114
rect 19944 16068 20168 16096
rect 19892 16050 19944 16056
rect 20168 16050 20220 16056
rect 20168 15904 20220 15910
rect 20168 15846 20220 15852
rect 19522 15736 19578 15745
rect 19522 15671 19578 15680
rect 19536 15570 19564 15671
rect 19524 15564 19576 15570
rect 19524 15506 19576 15512
rect 19522 15464 19578 15473
rect 19522 15399 19524 15408
rect 19576 15399 19578 15408
rect 19982 15464 20038 15473
rect 20180 15434 20208 15846
rect 19982 15399 20038 15408
rect 20168 15428 20220 15434
rect 19524 15370 19576 15376
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 19536 13530 19564 13670
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19996 13326 20024 15399
rect 20168 15370 20220 15376
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 20088 13938 20116 14214
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 20180 13394 20208 14894
rect 20168 13388 20220 13394
rect 20168 13330 20220 13336
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 20076 13252 20128 13258
rect 20076 13194 20128 13200
rect 20168 13252 20220 13258
rect 20168 13194 20220 13200
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19524 11824 19576 11830
rect 19524 11766 19576 11772
rect 19536 11286 19564 11766
rect 19524 11280 19576 11286
rect 19524 11222 19576 11228
rect 19996 11150 20024 12174
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 19614 10704 19670 10713
rect 19614 10639 19670 10648
rect 19892 10668 19944 10674
rect 19628 10538 19656 10639
rect 19892 10610 19944 10616
rect 19904 10577 19932 10610
rect 19890 10568 19946 10577
rect 19616 10532 19668 10538
rect 19890 10503 19946 10512
rect 19616 10474 19668 10480
rect 19260 9982 19380 10010
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19260 9500 19288 9982
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19352 9654 19380 9862
rect 19444 9761 19472 9998
rect 19996 9994 20024 11086
rect 19984 9988 20036 9994
rect 19984 9930 20036 9936
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19430 9752 19486 9761
rect 19574 9744 19882 9764
rect 19430 9687 19486 9696
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19798 9616 19854 9625
rect 19260 9472 19380 9500
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 19260 7886 19288 9318
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 19352 6882 19380 9472
rect 19444 8566 19472 9590
rect 19798 9551 19800 9560
rect 19852 9551 19854 9560
rect 19800 9522 19852 9528
rect 20088 9489 20116 13194
rect 20180 10441 20208 13194
rect 20272 12102 20300 16186
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20350 14648 20406 14657
rect 20350 14583 20406 14592
rect 20364 14482 20392 14583
rect 20352 14476 20404 14482
rect 20352 14418 20404 14424
rect 20364 12306 20392 14418
rect 20456 12850 20484 15642
rect 20548 15162 20576 18838
rect 20640 17882 20668 19790
rect 20628 17876 20680 17882
rect 20628 17818 20680 17824
rect 20732 17762 20760 20742
rect 20824 20602 20852 20878
rect 20812 20596 20864 20602
rect 20812 20538 20864 20544
rect 20824 20262 20852 20538
rect 20812 20256 20864 20262
rect 20812 20198 20864 20204
rect 20824 19666 20852 20198
rect 20916 19854 20944 22442
rect 21100 22438 21128 22986
rect 21088 22432 21140 22438
rect 21088 22374 21140 22380
rect 21100 19938 21128 22374
rect 21192 20466 21220 23054
rect 21364 22976 21416 22982
rect 21364 22918 21416 22924
rect 21376 21962 21404 22918
rect 21456 22568 21508 22574
rect 21456 22510 21508 22516
rect 21468 22234 21496 22510
rect 21456 22228 21508 22234
rect 21456 22170 21508 22176
rect 21560 22098 21588 23666
rect 21548 22092 21600 22098
rect 21652 22094 21680 29446
rect 21732 28008 21784 28014
rect 21732 27950 21784 27956
rect 21744 27674 21772 27950
rect 21732 27668 21784 27674
rect 21732 27610 21784 27616
rect 21836 22094 21864 31282
rect 22100 30728 22152 30734
rect 22100 30670 22152 30676
rect 22112 30122 22140 30670
rect 22192 30252 22244 30258
rect 22192 30194 22244 30200
rect 22100 30116 22152 30122
rect 22100 30058 22152 30064
rect 22112 29594 22140 30058
rect 22020 29566 22140 29594
rect 21916 29504 21968 29510
rect 21916 29446 21968 29452
rect 21928 28694 21956 29446
rect 22020 28694 22048 29566
rect 22100 29504 22152 29510
rect 22100 29446 22152 29452
rect 21916 28688 21968 28694
rect 21916 28630 21968 28636
rect 22008 28688 22060 28694
rect 22008 28630 22060 28636
rect 21928 28422 21956 28630
rect 22112 28558 22140 29446
rect 22204 29306 22232 30194
rect 22296 29594 22324 31622
rect 22388 31414 22416 31622
rect 22376 31408 22428 31414
rect 22376 31350 22428 31356
rect 22376 31272 22428 31278
rect 22376 31214 22428 31220
rect 22388 29850 22416 31214
rect 22376 29844 22428 29850
rect 22376 29786 22428 29792
rect 22296 29566 22416 29594
rect 22192 29300 22244 29306
rect 22192 29242 22244 29248
rect 22284 29232 22336 29238
rect 22284 29174 22336 29180
rect 22192 29164 22244 29170
rect 22192 29106 22244 29112
rect 22204 29073 22232 29106
rect 22190 29064 22246 29073
rect 22190 28999 22246 29008
rect 22100 28552 22152 28558
rect 22100 28494 22152 28500
rect 21916 28416 21968 28422
rect 21916 28358 21968 28364
rect 21928 28014 21956 28358
rect 21916 28008 21968 28014
rect 21916 27950 21968 27956
rect 22204 27674 22232 28999
rect 22296 28082 22324 29174
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22192 27668 22244 27674
rect 22192 27610 22244 27616
rect 22008 27532 22060 27538
rect 22008 27474 22060 27480
rect 22020 26926 22048 27474
rect 22204 27470 22232 27610
rect 22192 27464 22244 27470
rect 22192 27406 22244 27412
rect 22204 27130 22232 27406
rect 22192 27124 22244 27130
rect 22192 27066 22244 27072
rect 22008 26920 22060 26926
rect 22008 26862 22060 26868
rect 22020 26450 22048 26862
rect 22100 26784 22152 26790
rect 22100 26726 22152 26732
rect 22112 26518 22140 26726
rect 22100 26512 22152 26518
rect 22100 26454 22152 26460
rect 22008 26444 22060 26450
rect 22008 26386 22060 26392
rect 22100 26376 22152 26382
rect 22100 26318 22152 26324
rect 22112 26234 22140 26318
rect 21928 26206 22140 26234
rect 21928 25838 21956 26206
rect 22296 26042 22324 28018
rect 22284 26036 22336 26042
rect 22284 25978 22336 25984
rect 22100 25900 22152 25906
rect 22100 25842 22152 25848
rect 22284 25900 22336 25906
rect 22284 25842 22336 25848
rect 21916 25832 21968 25838
rect 21916 25774 21968 25780
rect 21916 25696 21968 25702
rect 21916 25638 21968 25644
rect 21928 23050 21956 25638
rect 22112 25362 22140 25842
rect 22296 25498 22324 25842
rect 22284 25492 22336 25498
rect 22284 25434 22336 25440
rect 22100 25356 22152 25362
rect 22100 25298 22152 25304
rect 22192 25220 22244 25226
rect 22192 25162 22244 25168
rect 22204 24750 22232 25162
rect 22192 24744 22244 24750
rect 22192 24686 22244 24692
rect 22284 24744 22336 24750
rect 22284 24686 22336 24692
rect 22296 24410 22324 24686
rect 22284 24404 22336 24410
rect 22284 24346 22336 24352
rect 22284 24200 22336 24206
rect 22284 24142 22336 24148
rect 22296 24070 22324 24142
rect 22284 24064 22336 24070
rect 22284 24006 22336 24012
rect 22192 23724 22244 23730
rect 22192 23666 22244 23672
rect 22204 23322 22232 23666
rect 22284 23656 22336 23662
rect 22284 23598 22336 23604
rect 22192 23316 22244 23322
rect 22192 23258 22244 23264
rect 21916 23044 21968 23050
rect 21916 22986 21968 22992
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22112 22710 22140 22918
rect 22296 22778 22324 23598
rect 22284 22772 22336 22778
rect 22284 22714 22336 22720
rect 22100 22704 22152 22710
rect 22100 22646 22152 22652
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 21652 22066 21772 22094
rect 21836 22066 21956 22094
rect 21548 22034 21600 22040
rect 21364 21956 21416 21962
rect 21364 21898 21416 21904
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 21100 19910 21312 19938
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 20824 19638 20944 19666
rect 20916 18034 20944 19638
rect 20996 19372 21048 19378
rect 20996 19314 21048 19320
rect 21008 18154 21036 19314
rect 20996 18148 21048 18154
rect 20996 18090 21048 18096
rect 21192 18086 21220 19790
rect 21284 18306 21312 19910
rect 21376 18970 21404 21898
rect 21560 21622 21588 22034
rect 21548 21616 21600 21622
rect 21548 21558 21600 21564
rect 21640 21616 21692 21622
rect 21640 21558 21692 21564
rect 21548 20460 21600 20466
rect 21548 20402 21600 20408
rect 21560 19922 21588 20402
rect 21548 19916 21600 19922
rect 21548 19858 21600 19864
rect 21364 18964 21416 18970
rect 21364 18906 21416 18912
rect 21284 18278 21404 18306
rect 21272 18148 21324 18154
rect 21272 18090 21324 18096
rect 20640 17734 20760 17762
rect 20824 18006 20944 18034
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 20536 15156 20588 15162
rect 20536 15098 20588 15104
rect 20536 14000 20588 14006
rect 20536 13942 20588 13948
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 20352 12300 20404 12306
rect 20352 12242 20404 12248
rect 20444 12300 20496 12306
rect 20444 12242 20496 12248
rect 20456 12170 20484 12242
rect 20444 12164 20496 12170
rect 20444 12106 20496 12112
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 20258 11928 20314 11937
rect 20258 11863 20314 11872
rect 20166 10432 20222 10441
rect 20166 10367 20222 10376
rect 20180 9654 20208 10367
rect 20168 9648 20220 9654
rect 20168 9590 20220 9596
rect 20074 9480 20130 9489
rect 20074 9415 20130 9424
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19432 8560 19484 8566
rect 19432 8502 19484 8508
rect 20088 8498 20116 9318
rect 20272 8650 20300 11863
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20364 10130 20392 11698
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20444 9988 20496 9994
rect 20444 9930 20496 9936
rect 20350 9616 20406 9625
rect 20350 9551 20352 9560
rect 20404 9551 20406 9560
rect 20352 9522 20404 9528
rect 20272 8622 20392 8650
rect 20260 8560 20312 8566
rect 20258 8528 20260 8537
rect 20312 8528 20314 8537
rect 20076 8492 20128 8498
rect 20258 8463 20314 8472
rect 20076 8434 20128 8440
rect 19432 7812 19484 7818
rect 19432 7754 19484 7760
rect 19260 6854 19380 6882
rect 19260 6390 19288 6854
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19248 6384 19300 6390
rect 19248 6326 19300 6332
rect 19248 6248 19300 6254
rect 19246 6216 19248 6225
rect 19300 6216 19302 6225
rect 19156 6180 19208 6186
rect 19246 6151 19302 6160
rect 19156 6122 19208 6128
rect 19168 5914 19196 6122
rect 19352 6118 19380 6734
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19156 5908 19208 5914
rect 19156 5850 19208 5856
rect 19352 5234 19380 6054
rect 19444 5914 19472 7754
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 19616 6112 19668 6118
rect 19996 6089 20024 6258
rect 19616 6054 19668 6060
rect 19982 6080 20038 6089
rect 19628 5914 19656 6054
rect 19982 6015 20038 6024
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19616 5908 19668 5914
rect 19616 5850 19668 5856
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 19996 5574 20024 5714
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 19246 4992 19302 5001
rect 19246 4927 19302 4936
rect 18984 2746 19104 2774
rect 18984 1766 19012 2746
rect 18972 1760 19024 1766
rect 18972 1702 19024 1708
rect 19260 800 19288 4927
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 19352 2514 19380 4626
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19996 4282 20024 4558
rect 19984 4276 20036 4282
rect 19536 4236 19840 4264
rect 19432 4208 19484 4214
rect 19536 4196 19564 4236
rect 19484 4168 19564 4196
rect 19432 4150 19484 4156
rect 19616 4140 19668 4146
rect 19616 4082 19668 4088
rect 19430 4040 19486 4049
rect 19430 3975 19486 3984
rect 19524 4004 19576 4010
rect 19444 3534 19472 3975
rect 19524 3946 19576 3952
rect 19536 3913 19564 3946
rect 19522 3904 19578 3913
rect 19522 3839 19578 3848
rect 19628 3738 19656 4082
rect 19616 3732 19668 3738
rect 19616 3674 19668 3680
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19812 3466 19840 4236
rect 19984 4218 20036 4224
rect 19982 4040 20038 4049
rect 19982 3975 20038 3984
rect 19800 3460 19852 3466
rect 19800 3402 19852 3408
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19340 2508 19392 2514
rect 19340 2450 19392 2456
rect 19444 1034 19472 3334
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19444 1006 19656 1034
rect 19628 800 19656 1006
rect 19996 800 20024 3975
rect 20088 3058 20116 8434
rect 20168 8016 20220 8022
rect 20168 7958 20220 7964
rect 20180 6730 20208 7958
rect 20364 7936 20392 8622
rect 20272 7908 20392 7936
rect 20272 7392 20300 7908
rect 20456 7886 20484 9930
rect 20548 9654 20576 13942
rect 20640 13870 20668 17734
rect 20718 17640 20774 17649
rect 20718 17575 20774 17584
rect 20732 17202 20760 17575
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20824 16810 20852 18006
rect 20902 17912 20958 17921
rect 20902 17847 20958 17856
rect 20916 17338 20944 17847
rect 20904 17332 20956 17338
rect 20904 17274 20956 17280
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 21008 17066 21036 17274
rect 21088 17264 21140 17270
rect 21088 17206 21140 17212
rect 20996 17060 21048 17066
rect 20996 17002 21048 17008
rect 21100 16998 21128 17206
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 20824 16782 20944 16810
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20732 13546 20760 14962
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20824 14414 20852 14758
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20916 13870 20944 16782
rect 21088 15564 21140 15570
rect 21088 15506 21140 15512
rect 21100 15450 21128 15506
rect 21008 15422 21128 15450
rect 20904 13864 20956 13870
rect 20904 13806 20956 13812
rect 20640 13530 20760 13546
rect 20628 13524 20760 13530
rect 20680 13518 20760 13524
rect 20628 13466 20680 13472
rect 21008 13410 21036 15422
rect 21088 13728 21140 13734
rect 21088 13670 21140 13676
rect 20916 13382 21036 13410
rect 20916 12866 20944 13382
rect 20996 13252 21048 13258
rect 20996 13194 21048 13200
rect 21008 12986 21036 13194
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 20720 12844 20772 12850
rect 20916 12838 21036 12866
rect 20720 12786 20772 12792
rect 20628 12640 20680 12646
rect 20628 12582 20680 12588
rect 20640 9738 20668 12582
rect 20732 11558 20760 12786
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 20916 12442 20944 12718
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 20812 12096 20864 12102
rect 20812 12038 20864 12044
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20732 10742 20760 11494
rect 20720 10736 20772 10742
rect 20720 10678 20772 10684
rect 20640 9710 20760 9738
rect 20732 9654 20760 9710
rect 20536 9648 20588 9654
rect 20536 9590 20588 9596
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20720 9444 20772 9450
rect 20720 9386 20772 9392
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20640 8430 20668 8910
rect 20628 8424 20680 8430
rect 20628 8366 20680 8372
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20352 7812 20404 7818
rect 20352 7754 20404 7760
rect 20364 7546 20392 7754
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20272 7364 20392 7392
rect 20260 7268 20312 7274
rect 20260 7210 20312 7216
rect 20168 6724 20220 6730
rect 20168 6666 20220 6672
rect 20168 6384 20220 6390
rect 20168 6326 20220 6332
rect 20180 3942 20208 6326
rect 20272 5302 20300 7210
rect 20364 5370 20392 7364
rect 20444 7336 20496 7342
rect 20444 7278 20496 7284
rect 20456 6322 20484 7278
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20442 6216 20498 6225
rect 20442 6151 20498 6160
rect 20456 5710 20484 6151
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 20352 5364 20404 5370
rect 20404 5324 20484 5352
rect 20352 5306 20404 5312
rect 20260 5296 20312 5302
rect 20260 5238 20312 5244
rect 20350 5128 20406 5137
rect 20350 5063 20406 5072
rect 20364 4214 20392 5063
rect 20352 4208 20404 4214
rect 20352 4150 20404 4156
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 20180 3534 20208 3878
rect 20272 3602 20300 4014
rect 20260 3596 20312 3602
rect 20260 3538 20312 3544
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 20272 3058 20300 3538
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 20260 3052 20312 3058
rect 20260 2994 20312 3000
rect 20364 800 20392 4014
rect 20456 3913 20484 5324
rect 20548 4758 20576 7686
rect 20640 6798 20668 8366
rect 20732 8022 20760 9386
rect 20720 8016 20772 8022
rect 20720 7958 20772 7964
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 20732 6662 20760 7686
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20720 5704 20772 5710
rect 20720 5646 20772 5652
rect 20536 4752 20588 4758
rect 20536 4694 20588 4700
rect 20548 4622 20576 4694
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20442 3904 20498 3913
rect 20442 3839 20498 3848
rect 20548 3194 20576 4082
rect 20640 3670 20668 4422
rect 20628 3664 20680 3670
rect 20628 3606 20680 3612
rect 20628 3460 20680 3466
rect 20628 3402 20680 3408
rect 20536 3188 20588 3194
rect 20536 3130 20588 3136
rect 20640 3126 20668 3402
rect 20732 3194 20760 5646
rect 20824 4214 20852 12038
rect 20916 11150 20944 12378
rect 21008 11354 21036 12838
rect 21100 12442 21128 13670
rect 21192 13462 21220 18022
rect 21180 13456 21232 13462
rect 21180 13398 21232 13404
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 21192 12782 21220 13262
rect 21180 12776 21232 12782
rect 21180 12718 21232 12724
rect 21088 12436 21140 12442
rect 21088 12378 21140 12384
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 20996 11076 21048 11082
rect 20996 11018 21048 11024
rect 20904 11008 20956 11014
rect 20904 10950 20956 10956
rect 20916 9926 20944 10950
rect 21008 10538 21036 11018
rect 20996 10532 21048 10538
rect 20996 10474 21048 10480
rect 21100 10266 21128 12378
rect 21178 11792 21234 11801
rect 21178 11727 21234 11736
rect 21088 10260 21140 10266
rect 21088 10202 21140 10208
rect 21192 9926 21220 11727
rect 21284 10690 21312 18090
rect 21376 15094 21404 18278
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21468 17202 21496 17614
rect 21456 17196 21508 17202
rect 21456 17138 21508 17144
rect 21548 16448 21600 16454
rect 21548 16390 21600 16396
rect 21560 15570 21588 16390
rect 21652 16046 21680 21558
rect 21744 19378 21772 22066
rect 21824 22024 21876 22030
rect 21824 21966 21876 21972
rect 21836 21554 21864 21966
rect 21824 21548 21876 21554
rect 21824 21490 21876 21496
rect 21836 20942 21864 21490
rect 21824 20936 21876 20942
rect 21824 20878 21876 20884
rect 21928 20516 21956 22066
rect 22100 22024 22152 22030
rect 22098 21992 22100 22001
rect 22152 21992 22154 22001
rect 22098 21927 22154 21936
rect 22100 21888 22152 21894
rect 22006 21856 22062 21865
rect 22100 21830 22152 21836
rect 22006 21791 22062 21800
rect 22020 21350 22048 21791
rect 22112 21729 22140 21830
rect 22098 21720 22154 21729
rect 22098 21655 22154 21664
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 22008 21344 22060 21350
rect 22008 21286 22060 21292
rect 22112 21026 22140 21490
rect 22204 21146 22232 22578
rect 22284 21956 22336 21962
rect 22284 21898 22336 21904
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 22296 21026 22324 21898
rect 22112 20998 22324 21026
rect 22008 20936 22060 20942
rect 22060 20884 22140 20890
rect 22008 20878 22140 20884
rect 22020 20862 22140 20878
rect 22296 20874 22324 20998
rect 22112 20618 22140 20862
rect 22284 20868 22336 20874
rect 22284 20810 22336 20816
rect 22112 20602 22232 20618
rect 22112 20596 22244 20602
rect 22112 20590 22192 20596
rect 22192 20538 22244 20544
rect 21928 20488 22048 20516
rect 21732 19372 21784 19378
rect 21732 19314 21784 19320
rect 21916 19372 21968 19378
rect 21916 19314 21968 19320
rect 21928 19242 21956 19314
rect 21916 19236 21968 19242
rect 21916 19178 21968 19184
rect 21732 19168 21784 19174
rect 21732 19110 21784 19116
rect 21744 17377 21772 19110
rect 21824 18692 21876 18698
rect 21824 18634 21876 18640
rect 21836 17882 21864 18634
rect 21928 18222 21956 19178
rect 22020 18426 22048 20488
rect 22388 19378 22416 29566
rect 22480 28762 22508 31826
rect 22572 31822 22600 32370
rect 23492 31958 23520 32370
rect 23572 32224 23624 32230
rect 23572 32166 23624 32172
rect 23480 31952 23532 31958
rect 23480 31894 23532 31900
rect 23388 31884 23440 31890
rect 23388 31826 23440 31832
rect 22560 31816 22612 31822
rect 22560 31758 22612 31764
rect 23204 31816 23256 31822
rect 23204 31758 23256 31764
rect 23020 31204 23072 31210
rect 23020 31146 23072 31152
rect 22560 30320 22612 30326
rect 22560 30262 22612 30268
rect 22468 28756 22520 28762
rect 22468 28698 22520 28704
rect 22572 26790 22600 30262
rect 22836 29776 22888 29782
rect 22836 29718 22888 29724
rect 22744 29504 22796 29510
rect 22744 29446 22796 29452
rect 22652 28620 22704 28626
rect 22652 28562 22704 28568
rect 22664 28422 22692 28562
rect 22756 28558 22784 29446
rect 22848 28966 22876 29718
rect 23032 29306 23060 31146
rect 23216 30122 23244 31758
rect 23296 31272 23348 31278
rect 23296 31214 23348 31220
rect 23308 30938 23336 31214
rect 23296 30932 23348 30938
rect 23296 30874 23348 30880
rect 23308 30394 23336 30874
rect 23400 30802 23428 31826
rect 23584 31754 23612 32166
rect 24596 32026 24624 32846
rect 24584 32020 24636 32026
rect 24584 31962 24636 31968
rect 24400 31884 24452 31890
rect 24400 31826 24452 31832
rect 23492 31748 23624 31754
rect 23492 31726 23572 31748
rect 23388 30796 23440 30802
rect 23388 30738 23440 30744
rect 23492 30682 23520 31726
rect 23572 31690 23624 31696
rect 24216 31680 24268 31686
rect 24216 31622 24268 31628
rect 24228 31346 24256 31622
rect 24216 31340 24268 31346
rect 24216 31282 24268 31288
rect 24032 31272 24084 31278
rect 24032 31214 24084 31220
rect 23400 30654 23520 30682
rect 23296 30388 23348 30394
rect 23296 30330 23348 30336
rect 23400 30274 23428 30654
rect 23480 30592 23532 30598
rect 23480 30534 23532 30540
rect 23308 30258 23428 30274
rect 23296 30252 23428 30258
rect 23348 30246 23428 30252
rect 23296 30194 23348 30200
rect 23204 30116 23256 30122
rect 23204 30058 23256 30064
rect 23308 30002 23336 30194
rect 23388 30184 23440 30190
rect 23388 30126 23440 30132
rect 23216 29974 23336 30002
rect 23112 29572 23164 29578
rect 23112 29514 23164 29520
rect 23020 29300 23072 29306
rect 23020 29242 23072 29248
rect 23124 29238 23152 29514
rect 23112 29232 23164 29238
rect 23112 29174 23164 29180
rect 22836 28960 22888 28966
rect 22836 28902 22888 28908
rect 22744 28552 22796 28558
rect 22744 28494 22796 28500
rect 22652 28416 22704 28422
rect 22652 28358 22704 28364
rect 22664 27402 22692 28358
rect 22756 27849 22784 28494
rect 22742 27840 22798 27849
rect 22742 27775 22798 27784
rect 22756 27470 22784 27775
rect 22744 27464 22796 27470
rect 22744 27406 22796 27412
rect 22652 27396 22704 27402
rect 22652 27338 22704 27344
rect 22560 26784 22612 26790
rect 22560 26726 22612 26732
rect 22572 25906 22600 26726
rect 22664 26382 22692 27338
rect 22756 27130 22784 27406
rect 22744 27124 22796 27130
rect 22744 27066 22796 27072
rect 22744 26988 22796 26994
rect 22744 26930 22796 26936
rect 22652 26376 22704 26382
rect 22652 26318 22704 26324
rect 22560 25900 22612 25906
rect 22560 25842 22612 25848
rect 22756 25294 22784 26930
rect 22848 26586 22876 28902
rect 23020 28416 23072 28422
rect 23020 28358 23072 28364
rect 22928 27464 22980 27470
rect 22928 27406 22980 27412
rect 22940 26994 22968 27406
rect 22928 26988 22980 26994
rect 22928 26930 22980 26936
rect 22928 26784 22980 26790
rect 22928 26726 22980 26732
rect 22836 26580 22888 26586
rect 22836 26522 22888 26528
rect 22940 25430 22968 26726
rect 23032 26518 23060 28358
rect 23124 26994 23152 29174
rect 23112 26988 23164 26994
rect 23112 26930 23164 26936
rect 23112 26852 23164 26858
rect 23112 26794 23164 26800
rect 23020 26512 23072 26518
rect 23020 26454 23072 26460
rect 22928 25424 22980 25430
rect 22928 25366 22980 25372
rect 23124 25294 23152 26794
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 23112 25288 23164 25294
rect 23112 25230 23164 25236
rect 22756 24970 22784 25230
rect 22560 24948 22612 24954
rect 22560 24890 22612 24896
rect 22664 24942 22784 24970
rect 22466 24848 22522 24857
rect 22466 24783 22468 24792
rect 22520 24783 22522 24792
rect 22468 24754 22520 24760
rect 22572 24410 22600 24890
rect 22664 24682 22692 24942
rect 23124 24834 23152 25230
rect 22756 24818 23152 24834
rect 22744 24812 23152 24818
rect 22796 24806 23152 24812
rect 22744 24754 22796 24760
rect 22652 24676 22704 24682
rect 22652 24618 22704 24624
rect 22560 24404 22612 24410
rect 22560 24346 22612 24352
rect 22664 24206 22692 24618
rect 22468 24200 22520 24206
rect 22468 24142 22520 24148
rect 22652 24200 22704 24206
rect 22652 24142 22704 24148
rect 23112 24200 23164 24206
rect 23112 24142 23164 24148
rect 22480 23730 22508 24142
rect 22468 23724 22520 23730
rect 22468 23666 22520 23672
rect 22664 23662 22692 24142
rect 22744 24132 22796 24138
rect 22744 24074 22796 24080
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22560 22976 22612 22982
rect 22560 22918 22612 22924
rect 22468 22160 22520 22166
rect 22468 22102 22520 22108
rect 22480 22030 22508 22102
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 22480 21554 22508 21966
rect 22468 21548 22520 21554
rect 22468 21490 22520 21496
rect 22572 21486 22600 22918
rect 22756 22001 22784 24074
rect 23124 24070 23152 24142
rect 23112 24064 23164 24070
rect 23112 24006 23164 24012
rect 23124 23186 23152 24006
rect 23112 23180 23164 23186
rect 23112 23122 23164 23128
rect 22928 22976 22980 22982
rect 22928 22918 22980 22924
rect 22940 22778 22968 22918
rect 22928 22772 22980 22778
rect 22928 22714 22980 22720
rect 22928 22636 22980 22642
rect 22928 22578 22980 22584
rect 22940 22030 22968 22578
rect 23216 22094 23244 29974
rect 23400 29850 23428 30126
rect 23388 29844 23440 29850
rect 23388 29786 23440 29792
rect 23296 29640 23348 29646
rect 23296 29582 23348 29588
rect 23308 28558 23336 29582
rect 23492 29034 23520 30534
rect 24044 30394 24072 31214
rect 24412 30802 24440 31826
rect 24584 31748 24636 31754
rect 24584 31690 24636 31696
rect 24596 31346 24624 31690
rect 24780 31346 24808 32914
rect 25412 32428 25464 32434
rect 25412 32370 25464 32376
rect 25228 32224 25280 32230
rect 25228 32166 25280 32172
rect 25240 31822 25268 32166
rect 25228 31816 25280 31822
rect 25228 31758 25280 31764
rect 25044 31680 25096 31686
rect 25044 31622 25096 31628
rect 25056 31414 25084 31622
rect 25424 31482 25452 32370
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 25412 31476 25464 31482
rect 25412 31418 25464 31424
rect 25044 31408 25096 31414
rect 25044 31350 25096 31356
rect 24584 31340 24636 31346
rect 24584 31282 24636 31288
rect 24768 31340 24820 31346
rect 24768 31282 24820 31288
rect 24400 30796 24452 30802
rect 24400 30738 24452 30744
rect 24584 30728 24636 30734
rect 24584 30670 24636 30676
rect 24032 30388 24084 30394
rect 24032 30330 24084 30336
rect 24032 30252 24084 30258
rect 24032 30194 24084 30200
rect 23664 30048 23716 30054
rect 23664 29990 23716 29996
rect 23676 29306 23704 29990
rect 23664 29300 23716 29306
rect 23664 29242 23716 29248
rect 24044 29170 24072 30194
rect 24596 29238 24624 30670
rect 24860 30252 24912 30258
rect 24860 30194 24912 30200
rect 24584 29232 24636 29238
rect 24584 29174 24636 29180
rect 24032 29164 24084 29170
rect 24032 29106 24084 29112
rect 23480 29028 23532 29034
rect 23480 28970 23532 28976
rect 23296 28552 23348 28558
rect 23296 28494 23348 28500
rect 23664 28552 23716 28558
rect 23664 28494 23716 28500
rect 23848 28552 23900 28558
rect 23848 28494 23900 28500
rect 23308 27674 23336 28494
rect 23676 28150 23704 28494
rect 23664 28144 23716 28150
rect 23664 28086 23716 28092
rect 23756 28076 23808 28082
rect 23756 28018 23808 28024
rect 23296 27668 23348 27674
rect 23296 27610 23348 27616
rect 23768 27402 23796 28018
rect 23860 27606 23888 28494
rect 23940 28484 23992 28490
rect 23940 28426 23992 28432
rect 23952 28014 23980 28426
rect 23940 28008 23992 28014
rect 23940 27950 23992 27956
rect 23848 27600 23900 27606
rect 23848 27542 23900 27548
rect 23756 27396 23808 27402
rect 23756 27338 23808 27344
rect 23664 26444 23716 26450
rect 23664 26386 23716 26392
rect 23296 26376 23348 26382
rect 23296 26318 23348 26324
rect 23308 23322 23336 26318
rect 23480 26240 23532 26246
rect 23480 26182 23532 26188
rect 23388 25968 23440 25974
rect 23388 25910 23440 25916
rect 23400 25786 23428 25910
rect 23492 25906 23520 26182
rect 23676 26042 23704 26386
rect 23664 26036 23716 26042
rect 23664 25978 23716 25984
rect 24044 25906 24072 29106
rect 24400 29028 24452 29034
rect 24400 28970 24452 28976
rect 24412 27470 24440 28970
rect 24596 28082 24624 29174
rect 24872 29102 24900 30194
rect 25056 29730 25084 31350
rect 26240 31340 26292 31346
rect 26240 31282 26292 31288
rect 26056 31136 26108 31142
rect 26056 31078 26108 31084
rect 26068 30666 26096 31078
rect 26056 30660 26108 30666
rect 26056 30602 26108 30608
rect 26252 30394 26280 31282
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 26424 30728 26476 30734
rect 26424 30670 26476 30676
rect 26240 30388 26292 30394
rect 26240 30330 26292 30336
rect 25136 30252 25188 30258
rect 25136 30194 25188 30200
rect 25320 30252 25372 30258
rect 25320 30194 25372 30200
rect 25148 29850 25176 30194
rect 25136 29844 25188 29850
rect 25136 29786 25188 29792
rect 25056 29702 25176 29730
rect 24952 29504 25004 29510
rect 24952 29446 25004 29452
rect 24964 29238 24992 29446
rect 24952 29232 25004 29238
rect 24952 29174 25004 29180
rect 24860 29096 24912 29102
rect 24860 29038 24912 29044
rect 24768 28620 24820 28626
rect 24768 28562 24820 28568
rect 24584 28076 24636 28082
rect 24584 28018 24636 28024
rect 24584 27872 24636 27878
rect 24584 27814 24636 27820
rect 24596 27470 24624 27814
rect 24780 27470 24808 28562
rect 24400 27464 24452 27470
rect 24400 27406 24452 27412
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 24768 27464 24820 27470
rect 24768 27406 24820 27412
rect 24952 27328 25004 27334
rect 24952 27270 25004 27276
rect 24676 26852 24728 26858
rect 24676 26794 24728 26800
rect 24400 26376 24452 26382
rect 24400 26318 24452 26324
rect 23480 25900 23532 25906
rect 23480 25842 23532 25848
rect 23664 25900 23716 25906
rect 23664 25842 23716 25848
rect 24032 25900 24084 25906
rect 24032 25842 24084 25848
rect 23676 25786 23704 25842
rect 23400 25758 23704 25786
rect 24044 25702 24072 25842
rect 24412 25702 24440 26318
rect 24688 25838 24716 26794
rect 24964 26382 24992 27270
rect 24952 26376 25004 26382
rect 24952 26318 25004 26324
rect 24676 25832 24728 25838
rect 24676 25774 24728 25780
rect 24032 25696 24084 25702
rect 24032 25638 24084 25644
rect 24400 25696 24452 25702
rect 24400 25638 24452 25644
rect 24412 25294 24440 25638
rect 24400 25288 24452 25294
rect 24400 25230 24452 25236
rect 24584 25288 24636 25294
rect 24584 25230 24636 25236
rect 23664 25152 23716 25158
rect 23664 25094 23716 25100
rect 23676 24886 23704 25094
rect 23664 24880 23716 24886
rect 23664 24822 23716 24828
rect 23480 24064 23532 24070
rect 23480 24006 23532 24012
rect 23296 23316 23348 23322
rect 23296 23258 23348 23264
rect 23308 22574 23336 23258
rect 23296 22568 23348 22574
rect 23296 22510 23348 22516
rect 23032 22066 23244 22094
rect 22928 22024 22980 22030
rect 22742 21992 22798 22001
rect 23032 22012 23060 22066
rect 23032 21984 23336 22012
rect 22928 21966 22980 21972
rect 22742 21927 22798 21936
rect 22836 21956 22888 21962
rect 22652 21888 22704 21894
rect 22652 21830 22704 21836
rect 22560 21480 22612 21486
rect 22560 21422 22612 21428
rect 22468 21344 22520 21350
rect 22468 21286 22520 21292
rect 22480 20534 22508 21286
rect 22468 20528 22520 20534
rect 22468 20470 22520 20476
rect 22664 19854 22692 21830
rect 22756 20058 22784 21927
rect 22836 21898 22888 21904
rect 22848 21865 22876 21898
rect 23020 21888 23072 21894
rect 22834 21856 22890 21865
rect 23020 21830 23072 21836
rect 22834 21791 22890 21800
rect 22928 21616 22980 21622
rect 22928 21558 22980 21564
rect 22836 21480 22888 21486
rect 22836 21422 22888 21428
rect 22848 20330 22876 21422
rect 22940 20942 22968 21558
rect 22928 20936 22980 20942
rect 22928 20878 22980 20884
rect 22836 20324 22888 20330
rect 22836 20266 22888 20272
rect 22744 20052 22796 20058
rect 22744 19994 22796 20000
rect 22652 19848 22704 19854
rect 22652 19790 22704 19796
rect 23032 19666 23060 21830
rect 23204 20936 23256 20942
rect 23204 20878 23256 20884
rect 23216 20602 23244 20878
rect 23308 20754 23336 21984
rect 23388 20936 23440 20942
rect 23492 20924 23520 24006
rect 24308 23792 24360 23798
rect 24308 23734 24360 23740
rect 23572 23724 23624 23730
rect 23572 23666 23624 23672
rect 23756 23724 23808 23730
rect 23756 23666 23808 23672
rect 23584 23050 23612 23666
rect 23768 23186 23796 23666
rect 23940 23656 23992 23662
rect 23940 23598 23992 23604
rect 23756 23180 23808 23186
rect 23756 23122 23808 23128
rect 23572 23044 23624 23050
rect 23572 22986 23624 22992
rect 23584 22710 23612 22986
rect 23572 22704 23624 22710
rect 23572 22646 23624 22652
rect 23768 22642 23796 23122
rect 23756 22636 23808 22642
rect 23756 22578 23808 22584
rect 23768 22030 23796 22578
rect 23756 22024 23808 22030
rect 23756 21966 23808 21972
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 23676 21554 23704 21830
rect 23756 21616 23808 21622
rect 23756 21558 23808 21564
rect 23664 21548 23716 21554
rect 23664 21490 23716 21496
rect 23664 21412 23716 21418
rect 23664 21354 23716 21360
rect 23676 21078 23704 21354
rect 23664 21072 23716 21078
rect 23664 21014 23716 21020
rect 23440 20896 23520 20924
rect 23388 20878 23440 20884
rect 23308 20726 23428 20754
rect 23204 20596 23256 20602
rect 23204 20538 23256 20544
rect 22664 19638 23060 19666
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 22376 19372 22428 19378
rect 22376 19314 22428 19320
rect 22008 18420 22060 18426
rect 22008 18362 22060 18368
rect 22112 18358 22140 19314
rect 22296 19242 22508 19258
rect 22192 19236 22244 19242
rect 22192 19178 22244 19184
rect 22296 19236 22520 19242
rect 22296 19230 22468 19236
rect 22100 18352 22152 18358
rect 22100 18294 22152 18300
rect 21916 18216 21968 18222
rect 21916 18158 21968 18164
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 21824 17876 21876 17882
rect 21824 17818 21876 17824
rect 22112 17678 22140 18022
rect 22100 17672 22152 17678
rect 22100 17614 22152 17620
rect 21730 17368 21786 17377
rect 22204 17354 22232 19178
rect 22296 18902 22324 19230
rect 22468 19178 22520 19184
rect 22376 19168 22428 19174
rect 22376 19110 22428 19116
rect 22284 18896 22336 18902
rect 22284 18838 22336 18844
rect 22284 17672 22336 17678
rect 22284 17614 22336 17620
rect 22112 17338 22232 17354
rect 21730 17303 21786 17312
rect 22100 17332 22232 17338
rect 22152 17326 22232 17332
rect 22100 17274 22152 17280
rect 22296 17270 22324 17614
rect 22192 17264 22244 17270
rect 22190 17232 22192 17241
rect 22284 17264 22336 17270
rect 22244 17232 22246 17241
rect 22284 17206 22336 17212
rect 22190 17167 22246 17176
rect 21824 17128 21876 17134
rect 21822 17096 21824 17105
rect 21876 17096 21878 17105
rect 21822 17031 21878 17040
rect 21824 16788 21876 16794
rect 21824 16730 21876 16736
rect 21640 16040 21692 16046
rect 21640 15982 21692 15988
rect 21652 15638 21680 15982
rect 21640 15632 21692 15638
rect 21640 15574 21692 15580
rect 21548 15564 21600 15570
rect 21548 15506 21600 15512
rect 21548 15428 21600 15434
rect 21548 15370 21600 15376
rect 21364 15088 21416 15094
rect 21364 15030 21416 15036
rect 21376 14550 21404 15030
rect 21364 14544 21416 14550
rect 21364 14486 21416 14492
rect 21456 13184 21508 13190
rect 21456 13126 21508 13132
rect 21364 12912 21416 12918
rect 21364 12854 21416 12860
rect 21376 11286 21404 12854
rect 21468 12102 21496 13126
rect 21560 12442 21588 15370
rect 21652 13394 21680 15574
rect 21836 14958 21864 16730
rect 22192 16516 22244 16522
rect 22192 16458 22244 16464
rect 22100 16448 22152 16454
rect 22100 16390 22152 16396
rect 22008 16040 22060 16046
rect 22008 15982 22060 15988
rect 21916 15496 21968 15502
rect 22020 15450 22048 15982
rect 22112 15638 22140 16390
rect 22100 15632 22152 15638
rect 22100 15574 22152 15580
rect 21968 15444 22048 15450
rect 21916 15438 22048 15444
rect 21928 15422 22048 15438
rect 21824 14952 21876 14958
rect 21824 14894 21876 14900
rect 22020 14618 22048 15422
rect 22204 15162 22232 16458
rect 22284 15972 22336 15978
rect 22284 15914 22336 15920
rect 22296 15638 22324 15914
rect 22284 15632 22336 15638
rect 22284 15574 22336 15580
rect 22192 15156 22244 15162
rect 22192 15098 22244 15104
rect 22388 15026 22416 19110
rect 22468 18828 22520 18834
rect 22468 18770 22520 18776
rect 22480 16590 22508 18770
rect 22560 18760 22612 18766
rect 22560 18702 22612 18708
rect 22572 17678 22600 18702
rect 22560 17672 22612 17678
rect 22560 17614 22612 17620
rect 22468 16584 22520 16590
rect 22468 16526 22520 16532
rect 22468 15564 22520 15570
rect 22468 15506 22520 15512
rect 22376 15020 22428 15026
rect 22376 14962 22428 14968
rect 22100 14884 22152 14890
rect 22100 14826 22152 14832
rect 22008 14612 22060 14618
rect 22008 14554 22060 14560
rect 21824 14408 21876 14414
rect 21824 14350 21876 14356
rect 21732 14340 21784 14346
rect 21732 14282 21784 14288
rect 21640 13388 21692 13394
rect 21640 13330 21692 13336
rect 21744 13326 21772 14282
rect 21836 13734 21864 14350
rect 21916 13932 21968 13938
rect 22020 13920 22048 14554
rect 21968 13892 22048 13920
rect 21916 13874 21968 13880
rect 21824 13728 21876 13734
rect 21824 13670 21876 13676
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21928 12850 21956 13874
rect 22008 13184 22060 13190
rect 22008 13126 22060 13132
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 21548 12436 21600 12442
rect 21548 12378 21600 12384
rect 21640 12368 21692 12374
rect 21640 12310 21692 12316
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21364 11280 21416 11286
rect 21364 11222 21416 11228
rect 21284 10662 21404 10690
rect 20904 9920 20956 9926
rect 21180 9920 21232 9926
rect 20956 9868 21036 9874
rect 20904 9862 21036 9868
rect 21180 9862 21232 9868
rect 20916 9846 21036 9862
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20916 5914 20944 7346
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20812 4208 20864 4214
rect 20812 4150 20864 4156
rect 20812 3936 20864 3942
rect 20812 3878 20864 3884
rect 20720 3188 20772 3194
rect 20720 3130 20772 3136
rect 20628 3120 20680 3126
rect 20628 3062 20680 3068
rect 20824 2446 20852 3878
rect 20916 3398 20944 4966
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 21008 3058 21036 9846
rect 21376 9738 21404 10662
rect 21100 9710 21404 9738
rect 21100 3534 21128 9710
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 21192 9178 21220 9522
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 21284 8090 21312 9522
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 21376 9178 21404 9318
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21468 8294 21496 11698
rect 21548 11552 21600 11558
rect 21548 11494 21600 11500
rect 21560 9994 21588 11494
rect 21652 11354 21680 12310
rect 21928 11762 21956 12786
rect 22020 12782 22048 13126
rect 22008 12776 22060 12782
rect 22008 12718 22060 12724
rect 21916 11756 21968 11762
rect 21916 11698 21968 11704
rect 21732 11620 21784 11626
rect 21732 11562 21784 11568
rect 21640 11348 21692 11354
rect 21640 11290 21692 11296
rect 21640 11144 21692 11150
rect 21640 11086 21692 11092
rect 21548 9988 21600 9994
rect 21548 9930 21600 9936
rect 21456 8288 21508 8294
rect 21456 8230 21508 8236
rect 21652 8106 21680 11086
rect 21272 8084 21324 8090
rect 21272 8026 21324 8032
rect 21468 8078 21680 8106
rect 21468 6866 21496 8078
rect 21548 8016 21600 8022
rect 21548 7958 21600 7964
rect 21456 6860 21508 6866
rect 21456 6802 21508 6808
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 21364 6656 21416 6662
rect 21364 6598 21416 6604
rect 21180 6384 21232 6390
rect 21180 6326 21232 6332
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 20996 3052 21048 3058
rect 20996 2994 21048 3000
rect 21192 2938 21220 6326
rect 21284 5846 21312 6598
rect 21272 5840 21324 5846
rect 21272 5782 21324 5788
rect 21376 5710 21404 6598
rect 21456 6248 21508 6254
rect 21456 6190 21508 6196
rect 21468 5846 21496 6190
rect 21456 5840 21508 5846
rect 21456 5782 21508 5788
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 21454 4312 21510 4321
rect 21454 4247 21510 4256
rect 21272 4004 21324 4010
rect 21272 3946 21324 3952
rect 21284 3738 21312 3946
rect 21272 3732 21324 3738
rect 21272 3674 21324 3680
rect 21272 3392 21324 3398
rect 21272 3334 21324 3340
rect 21008 2910 21220 2938
rect 21284 2922 21312 3334
rect 21272 2916 21324 2922
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 20732 870 20852 898
rect 20732 800 20760 870
rect 17052 734 17356 762
rect 17406 0 17462 800
rect 17774 0 17830 800
rect 18142 0 18198 800
rect 18510 0 18566 800
rect 18878 0 18934 800
rect 19246 0 19302 800
rect 19614 0 19670 800
rect 19982 0 20038 800
rect 20350 0 20406 800
rect 20718 0 20774 800
rect 20824 762 20852 870
rect 21008 762 21036 2910
rect 21272 2858 21324 2864
rect 21088 2848 21140 2854
rect 21088 2790 21140 2796
rect 21180 2848 21232 2854
rect 21180 2790 21232 2796
rect 21100 2446 21128 2790
rect 21088 2440 21140 2446
rect 21088 2382 21140 2388
rect 21192 1034 21220 2790
rect 21100 1006 21220 1034
rect 21100 800 21128 1006
rect 21468 800 21496 4247
rect 21560 2650 21588 7958
rect 21744 7154 21772 11562
rect 21914 9480 21970 9489
rect 21914 9415 21970 9424
rect 21822 9208 21878 9217
rect 21822 9143 21878 9152
rect 21836 8906 21864 9143
rect 21928 9110 21956 9415
rect 21916 9104 21968 9110
rect 21916 9046 21968 9052
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 21652 7126 21772 7154
rect 21652 6322 21680 7126
rect 21732 6996 21784 7002
rect 21732 6938 21784 6944
rect 21640 6316 21692 6322
rect 21640 6258 21692 6264
rect 21744 4826 21772 6938
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 21836 6322 21864 6734
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 21914 5808 21970 5817
rect 21914 5743 21970 5752
rect 21928 5710 21956 5743
rect 21916 5704 21968 5710
rect 21916 5646 21968 5652
rect 21824 5568 21876 5574
rect 21824 5510 21876 5516
rect 21836 5234 21864 5510
rect 21824 5228 21876 5234
rect 21824 5170 21876 5176
rect 21732 4820 21784 4826
rect 21732 4762 21784 4768
rect 21824 4752 21876 4758
rect 21824 4694 21876 4700
rect 21732 3528 21784 3534
rect 21732 3470 21784 3476
rect 21744 3194 21772 3470
rect 21732 3188 21784 3194
rect 21732 3130 21784 3136
rect 21744 3058 21772 3130
rect 21732 3052 21784 3058
rect 21732 2994 21784 3000
rect 21548 2644 21600 2650
rect 21548 2586 21600 2592
rect 21836 800 21864 4694
rect 21914 3904 21970 3913
rect 21914 3839 21970 3848
rect 21928 3602 21956 3839
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 21928 2990 21956 3538
rect 22020 3534 22048 12718
rect 22112 12306 22140 14826
rect 22480 14482 22508 15506
rect 22572 15434 22600 17614
rect 22664 16454 22692 19638
rect 23020 19508 23072 19514
rect 23020 19450 23072 19456
rect 22928 18352 22980 18358
rect 22928 18294 22980 18300
rect 22836 18284 22888 18290
rect 22836 18226 22888 18232
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 22652 16448 22704 16454
rect 22652 16390 22704 16396
rect 22652 16176 22704 16182
rect 22652 16118 22704 16124
rect 22664 15706 22692 16118
rect 22652 15700 22704 15706
rect 22652 15642 22704 15648
rect 22756 15502 22784 17478
rect 22744 15496 22796 15502
rect 22744 15438 22796 15444
rect 22560 15428 22612 15434
rect 22560 15370 22612 15376
rect 22468 14476 22520 14482
rect 22468 14418 22520 14424
rect 22652 14408 22704 14414
rect 22652 14350 22704 14356
rect 22468 14272 22520 14278
rect 22468 14214 22520 14220
rect 22192 13728 22244 13734
rect 22192 13670 22244 13676
rect 22204 13326 22232 13670
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 22376 12640 22428 12646
rect 22376 12582 22428 12588
rect 22100 12300 22152 12306
rect 22100 12242 22152 12248
rect 22388 12238 22416 12582
rect 22376 12232 22428 12238
rect 22376 12174 22428 12180
rect 22192 11552 22244 11558
rect 22190 11520 22192 11529
rect 22284 11552 22336 11558
rect 22244 11520 22246 11529
rect 22284 11494 22336 11500
rect 22190 11455 22246 11464
rect 22296 10674 22324 11494
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22376 10056 22428 10062
rect 22376 9998 22428 10004
rect 22100 9512 22152 9518
rect 22098 9480 22100 9489
rect 22152 9480 22154 9489
rect 22098 9415 22154 9424
rect 22192 9444 22244 9450
rect 22192 9386 22244 9392
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 22112 8090 22140 8434
rect 22204 8294 22232 9386
rect 22284 9172 22336 9178
rect 22284 9114 22336 9120
rect 22192 8288 22244 8294
rect 22192 8230 22244 8236
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 22204 7954 22232 8230
rect 22296 8090 22324 9114
rect 22284 8084 22336 8090
rect 22284 8026 22336 8032
rect 22192 7948 22244 7954
rect 22192 7890 22244 7896
rect 22388 7546 22416 9998
rect 22480 9586 22508 14214
rect 22664 13938 22692 14350
rect 22652 13932 22704 13938
rect 22652 13874 22704 13880
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22572 13326 22600 13466
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 22664 12850 22692 13874
rect 22652 12844 22704 12850
rect 22652 12786 22704 12792
rect 22652 12096 22704 12102
rect 22652 12038 22704 12044
rect 22664 11082 22692 12038
rect 22652 11076 22704 11082
rect 22652 11018 22704 11024
rect 22664 10826 22692 11018
rect 22572 10798 22692 10826
rect 22468 9580 22520 9586
rect 22468 9522 22520 9528
rect 22468 7812 22520 7818
rect 22468 7754 22520 7760
rect 22376 7540 22428 7546
rect 22376 7482 22428 7488
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22112 5642 22140 7346
rect 22284 6316 22336 6322
rect 22284 6258 22336 6264
rect 22100 5636 22152 5642
rect 22100 5578 22152 5584
rect 22296 5166 22324 6258
rect 22374 5944 22430 5953
rect 22374 5879 22430 5888
rect 22388 5574 22416 5879
rect 22376 5568 22428 5574
rect 22376 5510 22428 5516
rect 22284 5160 22336 5166
rect 22284 5102 22336 5108
rect 22192 5024 22244 5030
rect 22192 4966 22244 4972
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 22112 4146 22140 4762
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 22100 3936 22152 3942
rect 22098 3904 22100 3913
rect 22152 3904 22154 3913
rect 22098 3839 22154 3848
rect 22204 3754 22232 4966
rect 22296 4214 22324 5102
rect 22480 4826 22508 7754
rect 22468 4820 22520 4826
rect 22468 4762 22520 4768
rect 22376 4616 22428 4622
rect 22376 4558 22428 4564
rect 22284 4208 22336 4214
rect 22284 4150 22336 4156
rect 22112 3726 22232 3754
rect 22008 3528 22060 3534
rect 22008 3470 22060 3476
rect 21916 2984 21968 2990
rect 21916 2926 21968 2932
rect 22112 2854 22140 3726
rect 22192 3664 22244 3670
rect 22192 3606 22244 3612
rect 22204 3058 22232 3606
rect 22296 3602 22324 4150
rect 22284 3596 22336 3602
rect 22284 3538 22336 3544
rect 22192 3052 22244 3058
rect 22192 2994 22244 3000
rect 22284 2984 22336 2990
rect 22284 2926 22336 2932
rect 22100 2848 22152 2854
rect 22100 2790 22152 2796
rect 22296 2774 22324 2926
rect 22388 2922 22416 4558
rect 22468 4276 22520 4282
rect 22468 4218 22520 4224
rect 22376 2916 22428 2922
rect 22376 2858 22428 2864
rect 22296 2746 22416 2774
rect 22388 2514 22416 2746
rect 22376 2508 22428 2514
rect 22376 2450 22428 2456
rect 22204 870 22324 898
rect 22204 800 22232 870
rect 20824 734 21036 762
rect 21086 0 21142 800
rect 21454 0 21510 800
rect 21822 0 21878 800
rect 22190 0 22246 800
rect 22296 762 22324 870
rect 22480 762 22508 4218
rect 22572 2446 22600 10798
rect 22652 10192 22704 10198
rect 22652 10134 22704 10140
rect 22664 9058 22692 10134
rect 22848 9738 22876 18226
rect 22940 17678 22968 18294
rect 22928 17672 22980 17678
rect 22928 17614 22980 17620
rect 23032 17490 23060 19450
rect 23216 19378 23244 20538
rect 23204 19372 23256 19378
rect 23204 19314 23256 19320
rect 23400 19174 23428 20726
rect 23492 20602 23520 20896
rect 23572 20868 23624 20874
rect 23572 20810 23624 20816
rect 23480 20596 23532 20602
rect 23480 20538 23532 20544
rect 23584 19334 23612 20810
rect 23676 20466 23704 21014
rect 23768 20942 23796 21558
rect 23952 21554 23980 23598
rect 24032 23520 24084 23526
rect 24032 23462 24084 23468
rect 24044 23118 24072 23462
rect 24032 23112 24084 23118
rect 24032 23054 24084 23060
rect 24124 22432 24176 22438
rect 24124 22374 24176 22380
rect 24136 21554 24164 22374
rect 23940 21548 23992 21554
rect 23940 21490 23992 21496
rect 24124 21548 24176 21554
rect 24124 21490 24176 21496
rect 23756 20936 23808 20942
rect 23756 20878 23808 20884
rect 23940 20800 23992 20806
rect 23940 20742 23992 20748
rect 23952 20466 23980 20742
rect 23664 20460 23716 20466
rect 23664 20402 23716 20408
rect 23940 20460 23992 20466
rect 23940 20402 23992 20408
rect 23584 19306 23888 19334
rect 23388 19168 23440 19174
rect 23388 19110 23440 19116
rect 23860 18630 23888 19306
rect 23940 18760 23992 18766
rect 23940 18702 23992 18708
rect 23664 18624 23716 18630
rect 23664 18566 23716 18572
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23112 18284 23164 18290
rect 23112 18226 23164 18232
rect 23124 17678 23152 18226
rect 23480 18216 23532 18222
rect 23676 18193 23704 18566
rect 23480 18158 23532 18164
rect 23662 18184 23718 18193
rect 23492 17882 23520 18158
rect 23662 18119 23718 18128
rect 23296 17876 23348 17882
rect 23480 17876 23532 17882
rect 23296 17818 23348 17824
rect 23400 17836 23480 17864
rect 23204 17808 23256 17814
rect 23204 17750 23256 17756
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 23032 17462 23152 17490
rect 22928 16992 22980 16998
rect 22928 16934 22980 16940
rect 22940 11898 22968 16934
rect 23020 16448 23072 16454
rect 23020 16390 23072 16396
rect 23032 15026 23060 16390
rect 23020 15020 23072 15026
rect 23020 14962 23072 14968
rect 23032 12782 23060 14962
rect 23020 12776 23072 12782
rect 23020 12718 23072 12724
rect 23124 12434 23152 17462
rect 23216 17270 23244 17750
rect 23204 17264 23256 17270
rect 23204 17206 23256 17212
rect 23216 13308 23244 17206
rect 23308 16096 23336 17818
rect 23400 17338 23428 17836
rect 23480 17818 23532 17824
rect 23860 17814 23888 18566
rect 23848 17808 23900 17814
rect 23848 17750 23900 17756
rect 23388 17332 23440 17338
rect 23388 17274 23440 17280
rect 23480 17332 23532 17338
rect 23480 17274 23532 17280
rect 23492 17241 23520 17274
rect 23478 17232 23534 17241
rect 23952 17202 23980 18702
rect 24216 18216 24268 18222
rect 24216 18158 24268 18164
rect 23478 17167 23534 17176
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 23572 17060 23624 17066
rect 23572 17002 23624 17008
rect 23388 16108 23440 16114
rect 23308 16068 23388 16096
rect 23308 15706 23336 16068
rect 23388 16050 23440 16056
rect 23388 15972 23440 15978
rect 23388 15914 23440 15920
rect 23296 15700 23348 15706
rect 23296 15642 23348 15648
rect 23308 14958 23336 15642
rect 23400 15570 23428 15914
rect 23478 15736 23534 15745
rect 23584 15706 23612 17002
rect 23756 16448 23808 16454
rect 23756 16390 23808 16396
rect 23478 15671 23534 15680
rect 23572 15700 23624 15706
rect 23388 15564 23440 15570
rect 23388 15506 23440 15512
rect 23492 15502 23520 15671
rect 23572 15642 23624 15648
rect 23480 15496 23532 15502
rect 23480 15438 23532 15444
rect 23572 15020 23624 15026
rect 23572 14962 23624 14968
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 23296 14816 23348 14822
rect 23296 14758 23348 14764
rect 23308 14006 23336 14758
rect 23480 14408 23532 14414
rect 23480 14350 23532 14356
rect 23296 14000 23348 14006
rect 23296 13942 23348 13948
rect 23296 13320 23348 13326
rect 23216 13280 23296 13308
rect 23296 13262 23348 13268
rect 23124 12406 23428 12434
rect 23296 12232 23348 12238
rect 23296 12174 23348 12180
rect 23112 12164 23164 12170
rect 23112 12106 23164 12112
rect 22928 11892 22980 11898
rect 22928 11834 22980 11840
rect 23124 11694 23152 12106
rect 23308 11898 23336 12174
rect 23296 11892 23348 11898
rect 23296 11834 23348 11840
rect 23112 11688 23164 11694
rect 23112 11630 23164 11636
rect 23124 11218 23152 11630
rect 23296 11280 23348 11286
rect 23296 11222 23348 11228
rect 23112 11212 23164 11218
rect 23112 11154 23164 11160
rect 23308 11098 23336 11222
rect 22940 11082 23336 11098
rect 22928 11076 23336 11082
rect 22980 11070 23336 11076
rect 22928 11018 22980 11024
rect 23296 10736 23348 10742
rect 23296 10678 23348 10684
rect 23308 10266 23336 10678
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 22848 9710 23336 9738
rect 22836 9580 22888 9586
rect 22836 9522 22888 9528
rect 22744 9376 22796 9382
rect 22744 9318 22796 9324
rect 22756 9178 22784 9318
rect 22848 9178 22876 9522
rect 22928 9444 22980 9450
rect 22928 9386 22980 9392
rect 22744 9172 22796 9178
rect 22744 9114 22796 9120
rect 22836 9172 22888 9178
rect 22836 9114 22888 9120
rect 22664 9030 22876 9058
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22650 6352 22706 6361
rect 22650 6287 22706 6296
rect 22664 5710 22692 6287
rect 22652 5704 22704 5710
rect 22652 5646 22704 5652
rect 22652 4820 22704 4826
rect 22652 4762 22704 4768
rect 22664 4282 22692 4762
rect 22652 4276 22704 4282
rect 22652 4218 22704 4224
rect 22756 3466 22784 7482
rect 22848 6322 22876 9030
rect 22940 7886 22968 9386
rect 22928 7880 22980 7886
rect 22928 7822 22980 7828
rect 22836 6316 22888 6322
rect 22836 6258 22888 6264
rect 22744 3460 22796 3466
rect 22744 3402 22796 3408
rect 22652 3120 22704 3126
rect 22652 3062 22704 3068
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 22664 2258 22692 3062
rect 22940 3058 22968 7822
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 22928 3052 22980 3058
rect 22928 2994 22980 3000
rect 22928 2916 22980 2922
rect 22928 2858 22980 2864
rect 22572 2230 22692 2258
rect 22572 800 22600 2230
rect 22940 800 22968 2858
rect 23032 2650 23060 7346
rect 23204 7200 23256 7206
rect 23204 7142 23256 7148
rect 23216 4622 23244 7142
rect 23308 6730 23336 9710
rect 23296 6724 23348 6730
rect 23296 6666 23348 6672
rect 23400 6662 23428 12406
rect 23492 10266 23520 14350
rect 23584 12986 23612 14962
rect 23664 13184 23716 13190
rect 23664 13126 23716 13132
rect 23572 12980 23624 12986
rect 23572 12922 23624 12928
rect 23676 12918 23704 13126
rect 23664 12912 23716 12918
rect 23664 12854 23716 12860
rect 23676 12442 23704 12854
rect 23664 12436 23716 12442
rect 23664 12378 23716 12384
rect 23664 12300 23716 12306
rect 23664 12242 23716 12248
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 23584 10810 23612 11086
rect 23572 10804 23624 10810
rect 23572 10746 23624 10752
rect 23480 10260 23532 10266
rect 23480 10202 23532 10208
rect 23492 9654 23520 10202
rect 23572 9920 23624 9926
rect 23572 9862 23624 9868
rect 23480 9648 23532 9654
rect 23480 9590 23532 9596
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 23492 6186 23520 7890
rect 23480 6180 23532 6186
rect 23308 6140 23480 6168
rect 23308 5642 23336 6140
rect 23480 6122 23532 6128
rect 23386 6080 23442 6089
rect 23386 6015 23442 6024
rect 23400 5642 23428 6015
rect 23296 5636 23348 5642
rect 23296 5578 23348 5584
rect 23388 5636 23440 5642
rect 23388 5578 23440 5584
rect 23584 5302 23612 9862
rect 23676 7954 23704 12242
rect 23768 11762 23796 16390
rect 24030 15600 24086 15609
rect 24030 15535 24086 15544
rect 23940 14816 23992 14822
rect 23940 14758 23992 14764
rect 23848 14340 23900 14346
rect 23848 14282 23900 14288
rect 23860 11898 23888 14282
rect 23952 13938 23980 14758
rect 23940 13932 23992 13938
rect 23940 13874 23992 13880
rect 24044 13818 24072 15535
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 23952 13790 24072 13818
rect 23952 12434 23980 13790
rect 24032 13184 24084 13190
rect 24032 13126 24084 13132
rect 24044 12850 24072 13126
rect 24136 12986 24164 14962
rect 24124 12980 24176 12986
rect 24124 12922 24176 12928
rect 24032 12844 24084 12850
rect 24032 12786 24084 12792
rect 24124 12708 24176 12714
rect 24124 12650 24176 12656
rect 23952 12406 24072 12434
rect 23848 11892 23900 11898
rect 23848 11834 23900 11840
rect 23860 11778 23888 11834
rect 23756 11756 23808 11762
rect 23860 11750 23980 11778
rect 23756 11698 23808 11704
rect 23952 11694 23980 11750
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 23754 11520 23810 11529
rect 23754 11455 23810 11464
rect 23768 11082 23796 11455
rect 23756 11076 23808 11082
rect 23756 11018 23808 11024
rect 23756 10124 23808 10130
rect 23756 10066 23808 10072
rect 23768 9178 23796 10066
rect 23848 9988 23900 9994
rect 23848 9930 23900 9936
rect 23756 9172 23808 9178
rect 23756 9114 23808 9120
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 23756 7744 23808 7750
rect 23756 7686 23808 7692
rect 23664 7404 23716 7410
rect 23664 7346 23716 7352
rect 23572 5296 23624 5302
rect 23572 5238 23624 5244
rect 23572 4752 23624 4758
rect 23572 4694 23624 4700
rect 23204 4616 23256 4622
rect 23204 4558 23256 4564
rect 23480 4480 23532 4486
rect 23480 4422 23532 4428
rect 23204 3936 23256 3942
rect 23204 3878 23256 3884
rect 23296 3936 23348 3942
rect 23296 3878 23348 3884
rect 23216 3738 23244 3878
rect 23204 3732 23256 3738
rect 23204 3674 23256 3680
rect 23112 3460 23164 3466
rect 23112 3402 23164 3408
rect 23124 2854 23152 3402
rect 23308 2922 23336 3878
rect 23492 3126 23520 4422
rect 23480 3120 23532 3126
rect 23480 3062 23532 3068
rect 23296 2916 23348 2922
rect 23296 2858 23348 2864
rect 23112 2848 23164 2854
rect 23112 2790 23164 2796
rect 23584 2774 23612 4694
rect 23676 4690 23704 7346
rect 23768 6798 23796 7686
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 23860 5914 23888 9930
rect 23940 9376 23992 9382
rect 23940 9318 23992 9324
rect 23952 8498 23980 9318
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 23952 7342 23980 7822
rect 24044 7478 24072 12406
rect 24136 12186 24164 12650
rect 24228 12306 24256 18158
rect 24320 15978 24348 23734
rect 24412 23662 24440 25230
rect 24492 24404 24544 24410
rect 24492 24346 24544 24352
rect 24400 23656 24452 23662
rect 24400 23598 24452 23604
rect 24504 23118 24532 24346
rect 24596 23866 24624 25230
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 25044 24608 25096 24614
rect 25044 24550 25096 24556
rect 24688 24274 24716 24550
rect 24676 24268 24728 24274
rect 24676 24210 24728 24216
rect 24952 24132 25004 24138
rect 24952 24074 25004 24080
rect 24964 23882 24992 24074
rect 24584 23860 24636 23866
rect 24584 23802 24636 23808
rect 24872 23854 24992 23882
rect 24872 23338 24900 23854
rect 25056 23798 25084 24550
rect 25044 23792 25096 23798
rect 25044 23734 25096 23740
rect 24952 23724 25004 23730
rect 24952 23666 25004 23672
rect 24780 23310 24900 23338
rect 24964 23322 24992 23666
rect 24952 23316 25004 23322
rect 24780 23254 24808 23310
rect 24952 23258 25004 23264
rect 24768 23248 24820 23254
rect 24768 23190 24820 23196
rect 24492 23112 24544 23118
rect 24492 23054 24544 23060
rect 24676 23044 24728 23050
rect 24676 22986 24728 22992
rect 24492 22568 24544 22574
rect 24492 22510 24544 22516
rect 24400 21956 24452 21962
rect 24400 21898 24452 21904
rect 24412 21350 24440 21898
rect 24400 21344 24452 21350
rect 24400 21286 24452 21292
rect 24412 20942 24440 21286
rect 24400 20936 24452 20942
rect 24400 20878 24452 20884
rect 24504 19922 24532 22510
rect 24688 22094 24716 22986
rect 25148 22094 25176 29702
rect 25228 29708 25280 29714
rect 25228 29650 25280 29656
rect 25240 28762 25268 29650
rect 25228 28756 25280 28762
rect 25228 28698 25280 28704
rect 25332 28558 25360 30194
rect 26436 29714 26464 30670
rect 26608 30592 26660 30598
rect 26608 30534 26660 30540
rect 26620 30326 26648 30534
rect 26608 30320 26660 30326
rect 26608 30262 26660 30268
rect 26424 29708 26476 29714
rect 26424 29650 26476 29656
rect 25872 29504 25924 29510
rect 25872 29446 25924 29452
rect 25884 29050 25912 29446
rect 26332 29232 26384 29238
rect 25976 29180 26332 29186
rect 25976 29174 26384 29180
rect 25976 29170 26372 29174
rect 25964 29164 26372 29170
rect 26016 29158 26372 29164
rect 25964 29106 26016 29112
rect 26056 29096 26108 29102
rect 25884 29044 26056 29050
rect 25884 29038 26108 29044
rect 25688 29028 25740 29034
rect 25688 28970 25740 28976
rect 25884 29022 26096 29038
rect 25320 28552 25372 28558
rect 25320 28494 25372 28500
rect 25332 28218 25360 28494
rect 25320 28212 25372 28218
rect 25320 28154 25372 28160
rect 25700 28082 25728 28970
rect 25884 28490 25912 29022
rect 26148 28960 26200 28966
rect 26148 28902 26200 28908
rect 25872 28484 25924 28490
rect 25872 28426 25924 28432
rect 25688 28076 25740 28082
rect 25688 28018 25740 28024
rect 25700 27470 25728 28018
rect 25780 28008 25832 28014
rect 25884 27996 25912 28426
rect 26056 28416 26108 28422
rect 26056 28358 26108 28364
rect 26068 28150 26096 28358
rect 26160 28218 26188 28902
rect 26332 28756 26384 28762
rect 26332 28698 26384 28704
rect 26344 28422 26372 28698
rect 26436 28558 26464 29650
rect 26620 29510 26648 30262
rect 27528 30252 27580 30258
rect 27528 30194 27580 30200
rect 26976 30184 27028 30190
rect 26976 30126 27028 30132
rect 26608 29504 26660 29510
rect 26608 29446 26660 29452
rect 26424 28552 26476 28558
rect 26424 28494 26476 28500
rect 26332 28416 26384 28422
rect 26332 28358 26384 28364
rect 26148 28212 26200 28218
rect 26148 28154 26200 28160
rect 26056 28144 26108 28150
rect 26056 28086 26108 28092
rect 25832 27968 25912 27996
rect 25780 27950 25832 27956
rect 25688 27464 25740 27470
rect 25688 27406 25740 27412
rect 25780 27464 25832 27470
rect 25780 27406 25832 27412
rect 25228 27396 25280 27402
rect 25228 27338 25280 27344
rect 25504 27396 25556 27402
rect 25504 27338 25556 27344
rect 25240 26790 25268 27338
rect 25516 27130 25544 27338
rect 25504 27124 25556 27130
rect 25504 27066 25556 27072
rect 25700 26926 25728 27406
rect 25792 27130 25820 27406
rect 25884 27146 25912 27968
rect 26160 27470 26188 28154
rect 26344 28014 26372 28358
rect 26332 28008 26384 28014
rect 26332 27950 26384 27956
rect 26148 27464 26200 27470
rect 26148 27406 26200 27412
rect 25884 27130 26096 27146
rect 25780 27124 25832 27130
rect 25780 27066 25832 27072
rect 25884 27124 26108 27130
rect 25884 27118 26056 27124
rect 25780 26988 25832 26994
rect 25780 26930 25832 26936
rect 25688 26920 25740 26926
rect 25688 26862 25740 26868
rect 25228 26784 25280 26790
rect 25228 26726 25280 26732
rect 24596 22066 24716 22094
rect 25056 22066 25176 22094
rect 24492 19916 24544 19922
rect 24492 19858 24544 19864
rect 24504 18766 24532 19858
rect 24492 18760 24544 18766
rect 24492 18702 24544 18708
rect 24504 18154 24532 18702
rect 24492 18148 24544 18154
rect 24492 18090 24544 18096
rect 24596 16522 24624 22066
rect 24676 22024 24728 22030
rect 24676 21966 24728 21972
rect 24688 21622 24716 21966
rect 24676 21616 24728 21622
rect 24676 21558 24728 21564
rect 24952 19168 25004 19174
rect 24952 19110 25004 19116
rect 24768 18284 24820 18290
rect 24820 18244 24900 18272
rect 24768 18226 24820 18232
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24584 16516 24636 16522
rect 24584 16458 24636 16464
rect 24688 16250 24716 17682
rect 24872 17678 24900 18244
rect 24964 17678 24992 19110
rect 25056 18290 25084 22066
rect 25136 20936 25188 20942
rect 25136 20878 25188 20884
rect 25148 20602 25176 20878
rect 25136 20596 25188 20602
rect 25136 20538 25188 20544
rect 25044 18284 25096 18290
rect 25044 18226 25096 18232
rect 24860 17672 24912 17678
rect 24860 17614 24912 17620
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 24858 17096 24914 17105
rect 24858 17031 24914 17040
rect 24872 16658 24900 17031
rect 25136 16992 25188 16998
rect 25136 16934 25188 16940
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 24676 16244 24728 16250
rect 24676 16186 24728 16192
rect 24584 16040 24636 16046
rect 24584 15982 24636 15988
rect 24308 15972 24360 15978
rect 24308 15914 24360 15920
rect 24596 15502 24624 15982
rect 24674 15600 24730 15609
rect 24872 15570 24900 16594
rect 24952 16108 25004 16114
rect 24952 16050 25004 16056
rect 24674 15535 24730 15544
rect 24860 15564 24912 15570
rect 24688 15502 24716 15535
rect 24860 15506 24912 15512
rect 24964 15552 24992 16050
rect 25044 15564 25096 15570
rect 24964 15524 25044 15552
rect 24584 15496 24636 15502
rect 24584 15438 24636 15444
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24860 15020 24912 15026
rect 24860 14962 24912 14968
rect 24584 14952 24636 14958
rect 24584 14894 24636 14900
rect 24596 14006 24624 14894
rect 24872 14618 24900 14962
rect 24964 14618 24992 15524
rect 25044 15506 25096 15512
rect 25044 15360 25096 15366
rect 25044 15302 25096 15308
rect 24860 14612 24912 14618
rect 24860 14554 24912 14560
rect 24952 14612 25004 14618
rect 24952 14554 25004 14560
rect 25056 14414 25084 15302
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 24584 14000 24636 14006
rect 24584 13942 24636 13948
rect 24596 13530 24624 13942
rect 24952 13728 25004 13734
rect 24952 13670 25004 13676
rect 24584 13524 24636 13530
rect 24584 13466 24636 13472
rect 24964 13258 24992 13670
rect 24952 13252 25004 13258
rect 24952 13194 25004 13200
rect 24584 12844 24636 12850
rect 24584 12786 24636 12792
rect 24308 12368 24360 12374
rect 24308 12310 24360 12316
rect 24216 12300 24268 12306
rect 24216 12242 24268 12248
rect 24136 12170 24256 12186
rect 24136 12164 24268 12170
rect 24136 12158 24216 12164
rect 24216 12106 24268 12112
rect 24228 11694 24256 12106
rect 24216 11688 24268 11694
rect 24216 11630 24268 11636
rect 24228 11286 24256 11630
rect 24216 11280 24268 11286
rect 24216 11222 24268 11228
rect 24320 11218 24348 12310
rect 24308 11212 24360 11218
rect 24308 11154 24360 11160
rect 24216 11144 24268 11150
rect 24216 11086 24268 11092
rect 24400 11144 24452 11150
rect 24400 11086 24452 11092
rect 24124 11076 24176 11082
rect 24124 11018 24176 11024
rect 24032 7472 24084 7478
rect 24032 7414 24084 7420
rect 23940 7336 23992 7342
rect 24136 7290 24164 11018
rect 24228 10742 24256 11086
rect 24308 11076 24360 11082
rect 24308 11018 24360 11024
rect 24216 10736 24268 10742
rect 24216 10678 24268 10684
rect 24320 10470 24348 11018
rect 24308 10464 24360 10470
rect 24308 10406 24360 10412
rect 24308 9716 24360 9722
rect 24308 9658 24360 9664
rect 24320 8838 24348 9658
rect 24412 9654 24440 11086
rect 24492 10600 24544 10606
rect 24492 10542 24544 10548
rect 24504 10305 24532 10542
rect 24490 10296 24546 10305
rect 24490 10231 24546 10240
rect 24400 9648 24452 9654
rect 24400 9590 24452 9596
rect 24412 9042 24440 9590
rect 24492 9580 24544 9586
rect 24492 9522 24544 9528
rect 24400 9036 24452 9042
rect 24400 8978 24452 8984
rect 24308 8832 24360 8838
rect 24308 8774 24360 8780
rect 24320 8498 24348 8774
rect 24504 8634 24532 9522
rect 24492 8628 24544 8634
rect 24492 8570 24544 8576
rect 24308 8492 24360 8498
rect 24308 8434 24360 8440
rect 24492 7812 24544 7818
rect 24492 7754 24544 7760
rect 24504 7478 24532 7754
rect 24216 7472 24268 7478
rect 24216 7414 24268 7420
rect 24492 7472 24544 7478
rect 24492 7414 24544 7420
rect 23940 7278 23992 7284
rect 24044 7262 24164 7290
rect 24044 7188 24072 7262
rect 23952 7160 24072 7188
rect 24124 7200 24176 7206
rect 23848 5908 23900 5914
rect 23848 5850 23900 5856
rect 23952 5030 23980 7160
rect 24124 7142 24176 7148
rect 24032 6928 24084 6934
rect 24032 6870 24084 6876
rect 23940 5024 23992 5030
rect 23940 4966 23992 4972
rect 23664 4684 23716 4690
rect 23664 4626 23716 4632
rect 23664 3392 23716 3398
rect 23664 3334 23716 3340
rect 23848 3392 23900 3398
rect 23848 3334 23900 3340
rect 23676 3126 23704 3334
rect 23860 3194 23888 3334
rect 23848 3188 23900 3194
rect 23848 3130 23900 3136
rect 23664 3120 23716 3126
rect 23664 3062 23716 3068
rect 23848 2916 23900 2922
rect 23848 2858 23900 2864
rect 23400 2746 23612 2774
rect 23020 2644 23072 2650
rect 23020 2586 23072 2592
rect 23400 800 23428 2746
rect 23860 1986 23888 2858
rect 24044 2446 24072 6870
rect 24136 5710 24164 7142
rect 24124 5704 24176 5710
rect 24124 5646 24176 5652
rect 24228 5370 24256 7414
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 24320 6866 24348 7346
rect 24400 7268 24452 7274
rect 24400 7210 24452 7216
rect 24412 6934 24440 7210
rect 24400 6928 24452 6934
rect 24400 6870 24452 6876
rect 24308 6860 24360 6866
rect 24308 6802 24360 6808
rect 24492 6792 24544 6798
rect 24492 6734 24544 6740
rect 24400 6656 24452 6662
rect 24400 6598 24452 6604
rect 24308 6316 24360 6322
rect 24308 6258 24360 6264
rect 24320 5642 24348 6258
rect 24412 5710 24440 6598
rect 24400 5704 24452 5710
rect 24400 5646 24452 5652
rect 24308 5636 24360 5642
rect 24308 5578 24360 5584
rect 24216 5364 24268 5370
rect 24216 5306 24268 5312
rect 24400 5092 24452 5098
rect 24400 5034 24452 5040
rect 24216 5024 24268 5030
rect 24216 4966 24268 4972
rect 24228 2514 24256 4966
rect 24412 4078 24440 5034
rect 24400 4072 24452 4078
rect 24400 4014 24452 4020
rect 24412 3602 24440 4014
rect 24400 3596 24452 3602
rect 24400 3538 24452 3544
rect 24412 2990 24440 3538
rect 24504 3194 24532 6734
rect 24596 3534 24624 12786
rect 25148 12434 25176 16934
rect 25240 15502 25268 26726
rect 25792 25770 25820 26930
rect 25884 26382 25912 27118
rect 26056 27066 26108 27072
rect 26160 26926 26188 27406
rect 26148 26920 26200 26926
rect 26148 26862 26200 26868
rect 25872 26376 25924 26382
rect 25872 26318 25924 26324
rect 26148 26308 26200 26314
rect 26148 26250 26200 26256
rect 26160 25906 26188 26250
rect 26240 26036 26292 26042
rect 26240 25978 26292 25984
rect 26148 25900 26200 25906
rect 26148 25842 26200 25848
rect 25504 25764 25556 25770
rect 25504 25706 25556 25712
rect 25780 25764 25832 25770
rect 25780 25706 25832 25712
rect 25516 24954 25544 25706
rect 25688 25220 25740 25226
rect 25688 25162 25740 25168
rect 26148 25220 26200 25226
rect 26148 25162 26200 25168
rect 25504 24948 25556 24954
rect 25504 24890 25556 24896
rect 25700 23866 25728 25162
rect 26160 24857 26188 25162
rect 26146 24848 26202 24857
rect 26146 24783 26202 24792
rect 26160 24750 26188 24783
rect 25964 24744 26016 24750
rect 25964 24686 26016 24692
rect 26148 24744 26200 24750
rect 26148 24686 26200 24692
rect 25976 23866 26004 24686
rect 26252 24682 26280 25978
rect 26240 24676 26292 24682
rect 26240 24618 26292 24624
rect 26056 24064 26108 24070
rect 26056 24006 26108 24012
rect 25688 23860 25740 23866
rect 25688 23802 25740 23808
rect 25964 23860 26016 23866
rect 25964 23802 26016 23808
rect 25596 23112 25648 23118
rect 25596 23054 25648 23060
rect 25412 22976 25464 22982
rect 25412 22918 25464 22924
rect 25424 22710 25452 22918
rect 25412 22704 25464 22710
rect 25412 22646 25464 22652
rect 25608 21690 25636 23054
rect 25596 21684 25648 21690
rect 25596 21626 25648 21632
rect 25872 21140 25924 21146
rect 25792 21100 25872 21128
rect 25688 20460 25740 20466
rect 25688 20402 25740 20408
rect 25700 20058 25728 20402
rect 25688 20052 25740 20058
rect 25688 19994 25740 20000
rect 25792 19378 25820 21100
rect 25872 21082 25924 21088
rect 25872 20324 25924 20330
rect 25872 20266 25924 20272
rect 25964 20324 26016 20330
rect 25964 20266 26016 20272
rect 25780 19372 25832 19378
rect 25780 19314 25832 19320
rect 25780 18692 25832 18698
rect 25780 18634 25832 18640
rect 25320 18352 25372 18358
rect 25320 18294 25372 18300
rect 25332 17678 25360 18294
rect 25596 18216 25648 18222
rect 25596 18158 25648 18164
rect 25608 17814 25636 18158
rect 25596 17808 25648 17814
rect 25596 17750 25648 17756
rect 25504 17740 25556 17746
rect 25504 17682 25556 17688
rect 25320 17672 25372 17678
rect 25320 17614 25372 17620
rect 25320 17536 25372 17542
rect 25320 17478 25372 17484
rect 25332 16998 25360 17478
rect 25320 16992 25372 16998
rect 25320 16934 25372 16940
rect 25412 16992 25464 16998
rect 25412 16934 25464 16940
rect 25424 15978 25452 16934
rect 25412 15972 25464 15978
rect 25412 15914 25464 15920
rect 25228 15496 25280 15502
rect 25228 15438 25280 15444
rect 25320 14068 25372 14074
rect 25320 14010 25372 14016
rect 25332 12850 25360 14010
rect 25320 12844 25372 12850
rect 25320 12786 25372 12792
rect 24964 12406 25176 12434
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24872 11830 24900 12038
rect 24860 11824 24912 11830
rect 24860 11766 24912 11772
rect 24964 11506 24992 12406
rect 25412 12300 25464 12306
rect 25412 12242 25464 12248
rect 25044 11688 25096 11694
rect 25044 11630 25096 11636
rect 24872 11478 24992 11506
rect 24872 10674 24900 11478
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 25056 10606 25084 11630
rect 25320 10668 25372 10674
rect 25320 10610 25372 10616
rect 25044 10600 25096 10606
rect 25044 10542 25096 10548
rect 25332 10305 25360 10610
rect 25424 10470 25452 12242
rect 25412 10464 25464 10470
rect 25412 10406 25464 10412
rect 25318 10296 25374 10305
rect 25318 10231 25374 10240
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 25412 10056 25464 10062
rect 25412 9998 25464 10004
rect 24860 9648 24912 9654
rect 24766 9616 24822 9625
rect 24860 9590 24912 9596
rect 24766 9551 24768 9560
rect 24820 9551 24822 9560
rect 24768 9522 24820 9528
rect 24676 9512 24728 9518
rect 24674 9480 24676 9489
rect 24728 9480 24730 9489
rect 24674 9415 24730 9424
rect 24766 9072 24822 9081
rect 24766 9007 24822 9016
rect 24780 7410 24808 9007
rect 24872 8838 24900 9590
rect 24964 9450 24992 9998
rect 25044 9988 25096 9994
rect 25044 9930 25096 9936
rect 24952 9444 25004 9450
rect 24952 9386 25004 9392
rect 24860 8832 24912 8838
rect 24860 8774 24912 8780
rect 24872 8430 24900 8774
rect 25056 8498 25084 9930
rect 25424 9722 25452 9998
rect 25320 9716 25372 9722
rect 25320 9658 25372 9664
rect 25412 9716 25464 9722
rect 25412 9658 25464 9664
rect 25332 9586 25360 9658
rect 25320 9580 25372 9586
rect 25320 9522 25372 9528
rect 25136 9444 25188 9450
rect 25136 9386 25188 9392
rect 25044 8492 25096 8498
rect 25044 8434 25096 8440
rect 24860 8424 24912 8430
rect 24860 8366 24912 8372
rect 25148 7886 25176 9386
rect 25516 9382 25544 17682
rect 25792 17338 25820 18634
rect 25884 18408 25912 20266
rect 25976 19417 26004 20266
rect 26068 20058 26096 24006
rect 26240 23112 26292 23118
rect 26240 23054 26292 23060
rect 26252 21962 26280 23054
rect 26240 21956 26292 21962
rect 26240 21898 26292 21904
rect 26252 21729 26280 21898
rect 26238 21720 26294 21729
rect 26238 21655 26294 21664
rect 26252 21622 26280 21655
rect 26240 21616 26292 21622
rect 26240 21558 26292 21564
rect 26240 20868 26292 20874
rect 26240 20810 26292 20816
rect 26148 20256 26200 20262
rect 26148 20198 26200 20204
rect 26056 20052 26108 20058
rect 26056 19994 26108 20000
rect 26160 19854 26188 20198
rect 26148 19848 26200 19854
rect 26148 19790 26200 19796
rect 26252 19514 26280 20810
rect 26240 19508 26292 19514
rect 26240 19450 26292 19456
rect 25962 19408 26018 19417
rect 26238 19408 26294 19417
rect 25962 19343 26018 19352
rect 26056 19372 26108 19378
rect 26238 19343 26240 19352
rect 26056 19314 26108 19320
rect 26292 19343 26294 19352
rect 26240 19314 26292 19320
rect 25884 18380 26004 18408
rect 25872 17672 25924 17678
rect 25872 17614 25924 17620
rect 25780 17332 25832 17338
rect 25780 17274 25832 17280
rect 25780 16652 25832 16658
rect 25884 16640 25912 17614
rect 25976 17542 26004 18380
rect 25964 17536 26016 17542
rect 25964 17478 26016 17484
rect 25962 17368 26018 17377
rect 25962 17303 26018 17312
rect 25976 17202 26004 17303
rect 25964 17196 26016 17202
rect 25964 17138 26016 17144
rect 25832 16612 25912 16640
rect 25780 16594 25832 16600
rect 25792 16114 25820 16594
rect 25780 16108 25832 16114
rect 25780 16050 25832 16056
rect 25596 15632 25648 15638
rect 25596 15574 25648 15580
rect 25608 13938 25636 15574
rect 26068 15162 26096 19314
rect 26240 19168 26292 19174
rect 26240 19110 26292 19116
rect 26252 18766 26280 19110
rect 26240 18760 26292 18766
rect 26240 18702 26292 18708
rect 26240 18624 26292 18630
rect 26240 18566 26292 18572
rect 26148 18216 26200 18222
rect 26146 18184 26148 18193
rect 26200 18184 26202 18193
rect 26252 18170 26280 18566
rect 26344 18290 26372 27950
rect 26516 24880 26568 24886
rect 26516 24822 26568 24828
rect 26528 24410 26556 24822
rect 26516 24404 26568 24410
rect 26516 24346 26568 24352
rect 26620 24290 26648 29446
rect 26700 29232 26752 29238
rect 26700 29174 26752 29180
rect 26528 24262 26648 24290
rect 26424 23588 26476 23594
rect 26424 23530 26476 23536
rect 26436 23186 26464 23530
rect 26424 23180 26476 23186
rect 26424 23122 26476 23128
rect 26424 22976 26476 22982
rect 26424 22918 26476 22924
rect 26436 22710 26464 22918
rect 26424 22704 26476 22710
rect 26424 22646 26476 22652
rect 26424 18828 26476 18834
rect 26424 18770 26476 18776
rect 26332 18284 26384 18290
rect 26332 18226 26384 18232
rect 26252 18142 26372 18170
rect 26146 18119 26202 18128
rect 26160 17814 26188 18119
rect 26148 17808 26200 17814
rect 26148 17750 26200 17756
rect 26148 17672 26200 17678
rect 26200 17632 26280 17660
rect 26148 17614 26200 17620
rect 26148 16584 26200 16590
rect 26148 16526 26200 16532
rect 26160 16402 26188 16526
rect 26252 16522 26280 17632
rect 26344 17134 26372 18142
rect 26436 17882 26464 18770
rect 26424 17876 26476 17882
rect 26424 17818 26476 17824
rect 26528 17678 26556 24262
rect 26712 24154 26740 29174
rect 26884 28552 26936 28558
rect 26884 28494 26936 28500
rect 26896 27062 26924 28494
rect 26988 28082 27016 30126
rect 27252 29504 27304 29510
rect 27252 29446 27304 29452
rect 27264 29170 27292 29446
rect 27540 29306 27568 30194
rect 28448 30048 28500 30054
rect 28448 29990 28500 29996
rect 28460 29646 28488 29990
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 28448 29640 28500 29646
rect 28448 29582 28500 29588
rect 27528 29300 27580 29306
rect 27528 29242 27580 29248
rect 27252 29164 27304 29170
rect 27252 29106 27304 29112
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 27804 28484 27856 28490
rect 27804 28426 27856 28432
rect 27816 28218 27844 28426
rect 27804 28212 27856 28218
rect 27804 28154 27856 28160
rect 26976 28076 27028 28082
rect 26976 28018 27028 28024
rect 26988 27538 27016 28018
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 28172 27600 28224 27606
rect 28172 27542 28224 27548
rect 26976 27532 27028 27538
rect 26976 27474 27028 27480
rect 26884 27056 26936 27062
rect 26884 26998 26936 27004
rect 26896 26450 26924 26998
rect 26988 26790 27016 27474
rect 27068 27328 27120 27334
rect 27068 27270 27120 27276
rect 27528 27328 27580 27334
rect 27528 27270 27580 27276
rect 26976 26784 27028 26790
rect 26976 26726 27028 26732
rect 26884 26444 26936 26450
rect 26884 26386 26936 26392
rect 26896 26042 26924 26386
rect 26976 26308 27028 26314
rect 26976 26250 27028 26256
rect 26884 26036 26936 26042
rect 26884 25978 26936 25984
rect 26792 25968 26844 25974
rect 26792 25910 26844 25916
rect 26620 24126 26740 24154
rect 26516 17672 26568 17678
rect 26516 17614 26568 17620
rect 26424 17332 26476 17338
rect 26424 17274 26476 17280
rect 26332 17128 26384 17134
rect 26332 17070 26384 17076
rect 26240 16516 26292 16522
rect 26240 16458 26292 16464
rect 26160 16374 26280 16402
rect 26252 16114 26280 16374
rect 26240 16108 26292 16114
rect 26240 16050 26292 16056
rect 26252 15434 26280 16050
rect 26344 15978 26372 17070
rect 26332 15972 26384 15978
rect 26332 15914 26384 15920
rect 26240 15428 26292 15434
rect 26240 15370 26292 15376
rect 26436 15178 26464 17274
rect 26620 16250 26648 24126
rect 26700 23792 26752 23798
rect 26700 23734 26752 23740
rect 26712 22438 26740 23734
rect 26700 22432 26752 22438
rect 26700 22374 26752 22380
rect 26712 22030 26740 22374
rect 26700 22024 26752 22030
rect 26700 21966 26752 21972
rect 26804 20874 26832 25910
rect 26988 25498 27016 26250
rect 26976 25492 27028 25498
rect 26976 25434 27028 25440
rect 27080 25294 27108 27270
rect 27160 26988 27212 26994
rect 27160 26930 27212 26936
rect 27172 26586 27200 26930
rect 27160 26580 27212 26586
rect 27160 26522 27212 26528
rect 27540 25974 27568 27270
rect 28184 26518 28212 27542
rect 28356 27464 28408 27470
rect 28356 27406 28408 27412
rect 28368 27130 28396 27406
rect 28356 27124 28408 27130
rect 28356 27066 28408 27072
rect 28448 27056 28500 27062
rect 28448 26998 28500 27004
rect 28172 26512 28224 26518
rect 28172 26454 28224 26460
rect 27528 25968 27580 25974
rect 27528 25910 27580 25916
rect 26884 25288 26936 25294
rect 26884 25230 26936 25236
rect 27068 25288 27120 25294
rect 27068 25230 27120 25236
rect 26896 21690 26924 25230
rect 27436 24676 27488 24682
rect 27436 24618 27488 24624
rect 26976 24608 27028 24614
rect 26976 24550 27028 24556
rect 26988 24274 27016 24550
rect 26976 24268 27028 24274
rect 26976 24210 27028 24216
rect 27160 24268 27212 24274
rect 27160 24210 27212 24216
rect 26988 23186 27016 24210
rect 27068 23724 27120 23730
rect 27068 23666 27120 23672
rect 26976 23180 27028 23186
rect 26976 23122 27028 23128
rect 26884 21684 26936 21690
rect 26884 21626 26936 21632
rect 26884 21344 26936 21350
rect 26884 21286 26936 21292
rect 26792 20868 26844 20874
rect 26792 20810 26844 20816
rect 26804 20058 26832 20810
rect 26896 20602 26924 21286
rect 27080 21146 27108 23666
rect 27172 23662 27200 24210
rect 27344 24132 27396 24138
rect 27344 24074 27396 24080
rect 27252 23724 27304 23730
rect 27252 23666 27304 23672
rect 27160 23656 27212 23662
rect 27160 23598 27212 23604
rect 27160 21548 27212 21554
rect 27160 21490 27212 21496
rect 27068 21140 27120 21146
rect 27068 21082 27120 21088
rect 26884 20596 26936 20602
rect 26884 20538 26936 20544
rect 26884 20460 26936 20466
rect 26884 20402 26936 20408
rect 26792 20052 26844 20058
rect 26792 19994 26844 20000
rect 26700 19780 26752 19786
rect 26700 19722 26752 19728
rect 26712 18970 26740 19722
rect 26700 18964 26752 18970
rect 26700 18906 26752 18912
rect 26608 16244 26660 16250
rect 26608 16186 26660 16192
rect 26516 16040 26568 16046
rect 26516 15982 26568 15988
rect 26056 15156 26108 15162
rect 26056 15098 26108 15104
rect 26344 15150 26464 15178
rect 26068 14482 26096 15098
rect 25688 14476 25740 14482
rect 25688 14418 25740 14424
rect 26056 14476 26108 14482
rect 26056 14418 26108 14424
rect 25700 13938 25728 14418
rect 25596 13932 25648 13938
rect 25596 13874 25648 13880
rect 25688 13932 25740 13938
rect 25688 13874 25740 13880
rect 25872 13932 25924 13938
rect 26056 13932 26108 13938
rect 25872 13874 25924 13880
rect 25976 13892 26056 13920
rect 25780 13796 25832 13802
rect 25780 13738 25832 13744
rect 25688 13184 25740 13190
rect 25688 13126 25740 13132
rect 25700 12918 25728 13126
rect 25688 12912 25740 12918
rect 25688 12854 25740 12860
rect 25792 12442 25820 13738
rect 25884 12782 25912 13874
rect 25976 13258 26004 13892
rect 26056 13874 26108 13880
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 26252 13326 26280 13670
rect 26240 13320 26292 13326
rect 26240 13262 26292 13268
rect 25964 13252 26016 13258
rect 25964 13194 26016 13200
rect 25976 12850 26004 13194
rect 25964 12844 26016 12850
rect 25964 12786 26016 12792
rect 25872 12776 25924 12782
rect 25872 12718 25924 12724
rect 25872 12640 25924 12646
rect 25872 12582 25924 12588
rect 25780 12436 25832 12442
rect 25780 12378 25832 12384
rect 25884 12170 25912 12582
rect 25976 12306 26004 12786
rect 26148 12436 26200 12442
rect 26148 12378 26200 12384
rect 25964 12300 26016 12306
rect 25964 12242 26016 12248
rect 25688 12164 25740 12170
rect 25688 12106 25740 12112
rect 25872 12164 25924 12170
rect 25872 12106 25924 12112
rect 25596 9444 25648 9450
rect 25596 9386 25648 9392
rect 25504 9376 25556 9382
rect 25504 9318 25556 9324
rect 25516 9110 25544 9318
rect 25504 9104 25556 9110
rect 25504 9046 25556 9052
rect 25608 8498 25636 9386
rect 25596 8492 25648 8498
rect 25596 8434 25648 8440
rect 25136 7880 25188 7886
rect 25136 7822 25188 7828
rect 25412 7880 25464 7886
rect 25412 7822 25464 7828
rect 25044 7812 25096 7818
rect 25044 7754 25096 7760
rect 24768 7404 24820 7410
rect 24768 7346 24820 7352
rect 24952 7200 25004 7206
rect 24952 7142 25004 7148
rect 24964 6934 24992 7142
rect 25056 6934 25084 7754
rect 25320 7404 25372 7410
rect 25320 7346 25372 7352
rect 24676 6928 24728 6934
rect 24676 6870 24728 6876
rect 24952 6928 25004 6934
rect 24952 6870 25004 6876
rect 25044 6928 25096 6934
rect 25044 6870 25096 6876
rect 24688 6458 24716 6870
rect 24768 6792 24820 6798
rect 24766 6760 24768 6769
rect 24820 6760 24822 6769
rect 24766 6695 24822 6704
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 24688 5234 24716 6394
rect 24860 6248 24912 6254
rect 24860 6190 24912 6196
rect 24768 6180 24820 6186
rect 24768 6122 24820 6128
rect 24780 5953 24808 6122
rect 24766 5944 24822 5953
rect 24766 5879 24822 5888
rect 24768 5636 24820 5642
rect 24768 5578 24820 5584
rect 24780 5545 24808 5578
rect 24766 5536 24822 5545
rect 24766 5471 24822 5480
rect 24872 5370 24900 6190
rect 24964 5846 24992 6870
rect 24952 5840 25004 5846
rect 24952 5782 25004 5788
rect 24860 5364 24912 5370
rect 24860 5306 24912 5312
rect 24676 5228 24728 5234
rect 24676 5170 24728 5176
rect 24964 5166 24992 5782
rect 24952 5160 25004 5166
rect 24952 5102 25004 5108
rect 24768 4548 24820 4554
rect 24768 4490 24820 4496
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24492 3188 24544 3194
rect 24492 3130 24544 3136
rect 24490 3088 24546 3097
rect 24490 3023 24546 3032
rect 24400 2984 24452 2990
rect 24400 2926 24452 2932
rect 24308 2848 24360 2854
rect 24308 2790 24360 2796
rect 24216 2508 24268 2514
rect 24216 2450 24268 2456
rect 24032 2440 24084 2446
rect 24032 2382 24084 2388
rect 24320 2378 24348 2790
rect 24308 2372 24360 2378
rect 24308 2314 24360 2320
rect 24124 2304 24176 2310
rect 24124 2246 24176 2252
rect 23768 1958 23888 1986
rect 23768 800 23796 1958
rect 24136 800 24164 2246
rect 24504 800 24532 3023
rect 24780 2854 24808 4490
rect 24952 4072 25004 4078
rect 24952 4014 25004 4020
rect 24768 2848 24820 2854
rect 24768 2790 24820 2796
rect 24964 2650 24992 4014
rect 25056 3602 25084 6870
rect 25136 6724 25188 6730
rect 25136 6666 25188 6672
rect 25148 4622 25176 6666
rect 25228 6656 25280 6662
rect 25228 6598 25280 6604
rect 25136 4616 25188 4622
rect 25136 4558 25188 4564
rect 25136 3732 25188 3738
rect 25136 3674 25188 3680
rect 25044 3596 25096 3602
rect 25044 3538 25096 3544
rect 25148 2990 25176 3674
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 24952 2644 25004 2650
rect 24952 2586 25004 2592
rect 24860 2576 24912 2582
rect 24860 2518 24912 2524
rect 24872 800 24900 2518
rect 25240 2446 25268 6598
rect 25332 4146 25360 7346
rect 25424 5545 25452 7822
rect 25504 7744 25556 7750
rect 25504 7686 25556 7692
rect 25516 6322 25544 7686
rect 25596 6792 25648 6798
rect 25596 6734 25648 6740
rect 25504 6316 25556 6322
rect 25504 6258 25556 6264
rect 25502 6216 25558 6225
rect 25502 6151 25558 6160
rect 25410 5536 25466 5545
rect 25410 5471 25466 5480
rect 25320 4140 25372 4146
rect 25320 4082 25372 4088
rect 25318 4040 25374 4049
rect 25318 3975 25374 3984
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 25332 2258 25360 3975
rect 25516 3738 25544 6151
rect 25504 3732 25556 3738
rect 25504 3674 25556 3680
rect 25608 3194 25636 6734
rect 25700 4214 25728 12106
rect 26160 11082 26188 12378
rect 26240 12232 26292 12238
rect 26240 12174 26292 12180
rect 26252 11354 26280 12174
rect 26240 11348 26292 11354
rect 26240 11290 26292 11296
rect 26148 11076 26200 11082
rect 26148 11018 26200 11024
rect 25780 11008 25832 11014
rect 25780 10950 25832 10956
rect 25792 10538 25820 10950
rect 25780 10532 25832 10538
rect 25780 10474 25832 10480
rect 25872 10464 25924 10470
rect 25872 10406 25924 10412
rect 25780 8492 25832 8498
rect 25780 8434 25832 8440
rect 25792 6746 25820 8434
rect 25884 6882 25912 10406
rect 26056 9580 26108 9586
rect 26056 9522 26108 9528
rect 26068 9489 26096 9522
rect 26054 9480 26110 9489
rect 26054 9415 26110 9424
rect 25964 9376 26016 9382
rect 25964 9318 26016 9324
rect 26056 9376 26108 9382
rect 26056 9318 26108 9324
rect 25976 8974 26004 9318
rect 25964 8968 26016 8974
rect 25964 8910 26016 8916
rect 26068 8634 26096 9318
rect 26056 8628 26108 8634
rect 26056 8570 26108 8576
rect 25964 8560 26016 8566
rect 26160 8514 26188 11018
rect 26240 10464 26292 10470
rect 26238 10432 26240 10441
rect 26292 10432 26294 10441
rect 26238 10367 26294 10376
rect 26240 9104 26292 9110
rect 26238 9072 26240 9081
rect 26292 9072 26294 9081
rect 26238 9007 26294 9016
rect 26344 8974 26372 15150
rect 26424 14068 26476 14074
rect 26424 14010 26476 14016
rect 26436 11762 26464 14010
rect 26528 12434 26556 15982
rect 26712 13326 26740 18906
rect 26896 18766 26924 20402
rect 26976 19848 27028 19854
rect 26976 19790 27028 19796
rect 26988 19378 27016 19790
rect 27172 19514 27200 21490
rect 27264 20330 27292 23666
rect 27356 23594 27384 24074
rect 27344 23588 27396 23594
rect 27344 23530 27396 23536
rect 27356 21418 27384 23530
rect 27448 23186 27476 24618
rect 27528 23792 27580 23798
rect 27528 23734 27580 23740
rect 27436 23180 27488 23186
rect 27436 23122 27488 23128
rect 27448 22778 27476 23122
rect 27540 22982 27568 23734
rect 28080 23112 28132 23118
rect 28080 23054 28132 23060
rect 27620 23044 27672 23050
rect 27620 22986 27672 22992
rect 27528 22976 27580 22982
rect 27528 22918 27580 22924
rect 27436 22772 27488 22778
rect 27436 22714 27488 22720
rect 27540 22642 27568 22918
rect 27528 22636 27580 22642
rect 27528 22578 27580 22584
rect 27344 21412 27396 21418
rect 27344 21354 27396 21360
rect 27528 20868 27580 20874
rect 27528 20810 27580 20816
rect 27436 20800 27488 20806
rect 27436 20742 27488 20748
rect 27344 20596 27396 20602
rect 27344 20538 27396 20544
rect 27252 20324 27304 20330
rect 27252 20266 27304 20272
rect 27264 20058 27292 20266
rect 27252 20052 27304 20058
rect 27252 19994 27304 20000
rect 27252 19712 27304 19718
rect 27252 19654 27304 19660
rect 27160 19508 27212 19514
rect 27160 19450 27212 19456
rect 26976 19372 27028 19378
rect 26976 19314 27028 19320
rect 26884 18760 26936 18766
rect 26884 18702 26936 18708
rect 26792 18420 26844 18426
rect 26792 18362 26844 18368
rect 26804 17134 26832 18362
rect 26988 18222 27016 19314
rect 27172 18766 27200 19450
rect 27160 18760 27212 18766
rect 27160 18702 27212 18708
rect 27160 18624 27212 18630
rect 27264 18612 27292 19654
rect 27356 19310 27384 20538
rect 27448 20466 27476 20742
rect 27540 20534 27568 20810
rect 27528 20528 27580 20534
rect 27528 20470 27580 20476
rect 27436 20460 27488 20466
rect 27436 20402 27488 20408
rect 27448 19417 27476 20402
rect 27632 20346 27660 22986
rect 27804 22704 27856 22710
rect 27804 22646 27856 22652
rect 27712 21548 27764 21554
rect 27712 21490 27764 21496
rect 27724 20942 27752 21490
rect 27712 20936 27764 20942
rect 27712 20878 27764 20884
rect 27528 20324 27580 20330
rect 27632 20318 27752 20346
rect 27528 20266 27580 20272
rect 27540 19854 27568 20266
rect 27620 20256 27672 20262
rect 27620 20198 27672 20204
rect 27528 19848 27580 19854
rect 27528 19790 27580 19796
rect 27632 19786 27660 20198
rect 27620 19780 27672 19786
rect 27620 19722 27672 19728
rect 27724 19718 27752 20318
rect 27712 19712 27764 19718
rect 27712 19654 27764 19660
rect 27434 19408 27490 19417
rect 27434 19343 27490 19352
rect 27712 19372 27764 19378
rect 27344 19304 27396 19310
rect 27344 19246 27396 19252
rect 27212 18584 27292 18612
rect 27160 18566 27212 18572
rect 27356 18578 27384 19246
rect 27448 18766 27476 19343
rect 27712 19314 27764 19320
rect 27724 18970 27752 19314
rect 27712 18964 27764 18970
rect 27712 18906 27764 18912
rect 27816 18902 27844 22646
rect 28092 22506 28120 23054
rect 28080 22500 28132 22506
rect 28080 22442 28132 22448
rect 28092 22098 28120 22442
rect 28080 22092 28132 22098
rect 28080 22034 28132 22040
rect 27896 21888 27948 21894
rect 27896 21830 27948 21836
rect 27988 21888 28040 21894
rect 27988 21830 28040 21836
rect 27908 20942 27936 21830
rect 28000 21010 28028 21830
rect 27988 21004 28040 21010
rect 27988 20946 28040 20952
rect 28092 20942 28120 22034
rect 27896 20936 27948 20942
rect 27896 20878 27948 20884
rect 28080 20936 28132 20942
rect 28080 20878 28132 20884
rect 27988 20868 28040 20874
rect 27988 20810 28040 20816
rect 27804 18896 27856 18902
rect 27804 18838 27856 18844
rect 27436 18760 27488 18766
rect 27436 18702 27488 18708
rect 27896 18692 27948 18698
rect 27896 18634 27948 18640
rect 27436 18624 27488 18630
rect 27356 18572 27436 18578
rect 27356 18566 27488 18572
rect 27356 18550 27476 18566
rect 26976 18216 27028 18222
rect 26976 18158 27028 18164
rect 26988 17746 27016 18158
rect 27252 18080 27304 18086
rect 27252 18022 27304 18028
rect 27068 17808 27120 17814
rect 27068 17750 27120 17756
rect 26976 17740 27028 17746
rect 26976 17682 27028 17688
rect 26884 17196 26936 17202
rect 26884 17138 26936 17144
rect 26792 17128 26844 17134
rect 26792 17070 26844 17076
rect 26804 16794 26832 17070
rect 26792 16788 26844 16794
rect 26792 16730 26844 16736
rect 26792 16652 26844 16658
rect 26792 16594 26844 16600
rect 26700 13320 26752 13326
rect 26700 13262 26752 13268
rect 26528 12406 26648 12434
rect 26516 11824 26568 11830
rect 26516 11766 26568 11772
rect 26424 11756 26476 11762
rect 26424 11698 26476 11704
rect 26528 11150 26556 11766
rect 26516 11144 26568 11150
rect 26516 11086 26568 11092
rect 26528 10742 26556 11086
rect 26516 10736 26568 10742
rect 26516 10678 26568 10684
rect 26620 9330 26648 12406
rect 26712 10266 26740 13262
rect 26804 12646 26832 16594
rect 26896 16114 26924 17138
rect 27080 17116 27108 17750
rect 27264 17338 27292 18022
rect 27528 17672 27580 17678
rect 27528 17614 27580 17620
rect 27160 17332 27212 17338
rect 27160 17274 27212 17280
rect 27252 17332 27304 17338
rect 27252 17274 27304 17280
rect 27172 17218 27200 17274
rect 27172 17202 27292 17218
rect 27540 17202 27568 17614
rect 27620 17536 27672 17542
rect 27620 17478 27672 17484
rect 27712 17536 27764 17542
rect 27712 17478 27764 17484
rect 27172 17196 27304 17202
rect 27172 17190 27252 17196
rect 27252 17138 27304 17144
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 27632 17134 27660 17478
rect 27344 17128 27396 17134
rect 27080 17088 27200 17116
rect 27068 16720 27120 16726
rect 27068 16662 27120 16668
rect 26976 16652 27028 16658
rect 26976 16594 27028 16600
rect 26884 16108 26936 16114
rect 26884 16050 26936 16056
rect 26988 15026 27016 16594
rect 27080 16114 27108 16662
rect 27068 16108 27120 16114
rect 27068 16050 27120 16056
rect 26976 15020 27028 15026
rect 26976 14962 27028 14968
rect 26988 14618 27016 14962
rect 26976 14612 27028 14618
rect 26976 14554 27028 14560
rect 26988 13530 27016 14554
rect 26976 13524 27028 13530
rect 26976 13466 27028 13472
rect 26988 12850 27016 13466
rect 27068 13388 27120 13394
rect 27068 13330 27120 13336
rect 26976 12844 27028 12850
rect 26896 12804 26976 12832
rect 26792 12640 26844 12646
rect 26792 12582 26844 12588
rect 26792 11756 26844 11762
rect 26792 11698 26844 11704
rect 26700 10260 26752 10266
rect 26700 10202 26752 10208
rect 26700 9512 26752 9518
rect 26700 9454 26752 9460
rect 26528 9302 26648 9330
rect 26332 8968 26384 8974
rect 26332 8910 26384 8916
rect 26344 8634 26372 8910
rect 26332 8628 26384 8634
rect 26332 8570 26384 8576
rect 25964 8502 26016 8508
rect 25976 8430 26004 8502
rect 26068 8486 26188 8514
rect 25964 8424 26016 8430
rect 25964 8366 26016 8372
rect 25964 7404 26016 7410
rect 25964 7346 26016 7352
rect 25976 7002 26004 7346
rect 25964 6996 26016 7002
rect 25964 6938 26016 6944
rect 25884 6854 26004 6882
rect 25792 6718 25912 6746
rect 25884 6225 25912 6718
rect 25870 6216 25926 6225
rect 25870 6151 25926 6160
rect 25780 5228 25832 5234
rect 25780 5170 25832 5176
rect 25688 4208 25740 4214
rect 25688 4150 25740 4156
rect 25792 4146 25820 5170
rect 25872 5160 25924 5166
rect 25872 5102 25924 5108
rect 25884 4758 25912 5102
rect 25872 4752 25924 4758
rect 25872 4694 25924 4700
rect 25780 4140 25832 4146
rect 25780 4082 25832 4088
rect 25872 3936 25924 3942
rect 25872 3878 25924 3884
rect 25596 3188 25648 3194
rect 25596 3130 25648 3136
rect 25504 2916 25556 2922
rect 25504 2858 25556 2864
rect 25516 2446 25544 2858
rect 25884 2774 25912 3878
rect 25976 3058 26004 6854
rect 26068 6066 26096 8486
rect 26528 7698 26556 9302
rect 26712 9058 26740 9454
rect 26620 9030 26740 9058
rect 26620 8974 26648 9030
rect 26608 8968 26660 8974
rect 26608 8910 26660 8916
rect 26700 8968 26752 8974
rect 26700 8910 26752 8916
rect 26608 8832 26660 8838
rect 26608 8774 26660 8780
rect 26620 7954 26648 8774
rect 26608 7948 26660 7954
rect 26608 7890 26660 7896
rect 26712 7886 26740 8910
rect 26700 7880 26752 7886
rect 26700 7822 26752 7828
rect 26700 7744 26752 7750
rect 26528 7670 26648 7698
rect 26700 7686 26752 7692
rect 26148 6792 26200 6798
rect 26148 6734 26200 6740
rect 26332 6792 26384 6798
rect 26332 6734 26384 6740
rect 26160 6186 26188 6734
rect 26240 6384 26292 6390
rect 26240 6326 26292 6332
rect 26148 6180 26200 6186
rect 26148 6122 26200 6128
rect 26068 6038 26188 6066
rect 26056 5092 26108 5098
rect 26056 5034 26108 5040
rect 26068 4622 26096 5034
rect 26056 4616 26108 4622
rect 26056 4558 26108 4564
rect 26068 4146 26096 4558
rect 26160 4146 26188 6038
rect 26252 5710 26280 6326
rect 26240 5704 26292 5710
rect 26240 5646 26292 5652
rect 26344 4146 26372 6734
rect 26516 6724 26568 6730
rect 26516 6666 26568 6672
rect 26424 6656 26476 6662
rect 26424 6598 26476 6604
rect 26056 4140 26108 4146
rect 26056 4082 26108 4088
rect 26148 4140 26200 4146
rect 26148 4082 26200 4088
rect 26332 4140 26384 4146
rect 26332 4082 26384 4088
rect 26068 3670 26096 4082
rect 26056 3664 26108 3670
rect 26056 3606 26108 3612
rect 25964 3052 26016 3058
rect 25964 2994 26016 3000
rect 26068 2922 26096 3606
rect 26436 3534 26464 6598
rect 26240 3528 26292 3534
rect 26240 3470 26292 3476
rect 26424 3528 26476 3534
rect 26424 3470 26476 3476
rect 26056 2916 26108 2922
rect 26056 2858 26108 2864
rect 25884 2746 26004 2774
rect 25596 2576 25648 2582
rect 25596 2518 25648 2524
rect 25504 2440 25556 2446
rect 25504 2382 25556 2388
rect 25240 2230 25360 2258
rect 25240 800 25268 2230
rect 25608 800 25636 2518
rect 25976 800 26004 2746
rect 26252 2446 26280 3470
rect 26332 3392 26384 3398
rect 26332 3334 26384 3340
rect 26240 2440 26292 2446
rect 26240 2382 26292 2388
rect 26344 800 26372 3334
rect 26528 2446 26556 6666
rect 26620 5914 26648 7670
rect 26608 5908 26660 5914
rect 26608 5850 26660 5856
rect 26620 5302 26648 5850
rect 26712 5642 26740 7686
rect 26700 5636 26752 5642
rect 26700 5578 26752 5584
rect 26608 5296 26660 5302
rect 26608 5238 26660 5244
rect 26804 4622 26832 11698
rect 26896 11626 26924 12804
rect 26976 12786 27028 12792
rect 26976 12640 27028 12646
rect 26976 12582 27028 12588
rect 26884 11620 26936 11626
rect 26884 11562 26936 11568
rect 26896 10130 26924 11562
rect 26988 10266 27016 12582
rect 27080 11354 27108 13330
rect 27172 12102 27200 17088
rect 27342 17096 27344 17105
rect 27620 17128 27672 17134
rect 27396 17096 27398 17105
rect 27620 17070 27672 17076
rect 27342 17031 27398 17040
rect 27344 16516 27396 16522
rect 27344 16458 27396 16464
rect 27356 16114 27384 16458
rect 27344 16108 27396 16114
rect 27344 16050 27396 16056
rect 27344 15972 27396 15978
rect 27344 15914 27396 15920
rect 27252 13184 27304 13190
rect 27252 13126 27304 13132
rect 27160 12096 27212 12102
rect 27160 12038 27212 12044
rect 27264 11830 27292 13126
rect 27252 11824 27304 11830
rect 27252 11766 27304 11772
rect 27068 11348 27120 11354
rect 27068 11290 27120 11296
rect 27068 11076 27120 11082
rect 27068 11018 27120 11024
rect 26976 10260 27028 10266
rect 26976 10202 27028 10208
rect 26884 10124 26936 10130
rect 26884 10066 26936 10072
rect 26884 9988 26936 9994
rect 26884 9930 26936 9936
rect 26896 9722 26924 9930
rect 26976 9920 27028 9926
rect 26976 9862 27028 9868
rect 26884 9716 26936 9722
rect 26884 9658 26936 9664
rect 26988 9586 27016 9862
rect 26976 9580 27028 9586
rect 26976 9522 27028 9528
rect 26884 8832 26936 8838
rect 26884 8774 26936 8780
rect 26896 7041 26924 8774
rect 26974 8256 27030 8265
rect 26974 8191 27030 8200
rect 26882 7032 26938 7041
rect 26882 6967 26938 6976
rect 26882 5944 26938 5953
rect 26882 5879 26884 5888
rect 26936 5879 26938 5888
rect 26884 5850 26936 5856
rect 26988 5624 27016 8191
rect 27080 7410 27108 11018
rect 27158 10296 27214 10305
rect 27158 10231 27214 10240
rect 27252 10260 27304 10266
rect 27172 9722 27200 10231
rect 27252 10202 27304 10208
rect 27160 9716 27212 9722
rect 27160 9658 27212 9664
rect 27264 9625 27292 10202
rect 27250 9616 27306 9625
rect 27250 9551 27306 9560
rect 27356 8974 27384 15914
rect 27620 15904 27672 15910
rect 27620 15846 27672 15852
rect 27632 15502 27660 15846
rect 27620 15496 27672 15502
rect 27620 15438 27672 15444
rect 27436 15360 27488 15366
rect 27436 15302 27488 15308
rect 27448 15094 27476 15302
rect 27436 15088 27488 15094
rect 27436 15030 27488 15036
rect 27528 14000 27580 14006
rect 27528 13942 27580 13948
rect 27436 13456 27488 13462
rect 27436 13398 27488 13404
rect 27448 12986 27476 13398
rect 27540 12986 27568 13942
rect 27620 13320 27672 13326
rect 27620 13262 27672 13268
rect 27436 12980 27488 12986
rect 27436 12922 27488 12928
rect 27528 12980 27580 12986
rect 27528 12922 27580 12928
rect 27436 12232 27488 12238
rect 27436 12174 27488 12180
rect 27448 10713 27476 12174
rect 27528 12096 27580 12102
rect 27528 12038 27580 12044
rect 27434 10704 27490 10713
rect 27434 10639 27436 10648
rect 27488 10639 27490 10648
rect 27436 10610 27488 10616
rect 27436 9988 27488 9994
rect 27436 9930 27488 9936
rect 27344 8968 27396 8974
rect 27344 8910 27396 8916
rect 27448 8838 27476 9930
rect 27436 8832 27488 8838
rect 27436 8774 27488 8780
rect 27540 8616 27568 12038
rect 27632 11150 27660 13262
rect 27724 13172 27752 17478
rect 27804 16448 27856 16454
rect 27804 16390 27856 16396
rect 27816 13308 27844 16390
rect 27908 15570 27936 18634
rect 28000 16454 28028 20810
rect 28080 18624 28132 18630
rect 28080 18566 28132 18572
rect 28092 17678 28120 18566
rect 28080 17672 28132 17678
rect 28080 17614 28132 17620
rect 28184 17610 28212 26454
rect 28460 26382 28488 26998
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 28448 26376 28500 26382
rect 28448 26318 28500 26324
rect 28460 25702 28488 26318
rect 28448 25696 28500 25702
rect 28448 25638 28500 25644
rect 28356 24812 28408 24818
rect 28356 24754 28408 24760
rect 28368 24410 28396 24754
rect 28356 24404 28408 24410
rect 28356 24346 28408 24352
rect 28356 23724 28408 23730
rect 28356 23666 28408 23672
rect 28264 23656 28316 23662
rect 28264 23598 28316 23604
rect 28276 23118 28304 23598
rect 28368 23322 28396 23666
rect 28356 23316 28408 23322
rect 28356 23258 28408 23264
rect 28460 23202 28488 25638
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 28540 24200 28592 24206
rect 28540 24142 28592 24148
rect 28552 23866 28580 24142
rect 28540 23860 28592 23866
rect 28540 23802 28592 23808
rect 29184 23724 29236 23730
rect 29184 23666 29236 23672
rect 29920 23724 29972 23730
rect 29920 23666 29972 23672
rect 29000 23520 29052 23526
rect 29000 23462 29052 23468
rect 28368 23174 28488 23202
rect 28264 23112 28316 23118
rect 28264 23054 28316 23060
rect 28276 22234 28304 23054
rect 28264 22228 28316 22234
rect 28264 22170 28316 22176
rect 28368 21978 28396 23174
rect 29012 23118 29040 23462
rect 29196 23322 29224 23666
rect 29644 23520 29696 23526
rect 29644 23462 29696 23468
rect 29184 23316 29236 23322
rect 29184 23258 29236 23264
rect 28448 23112 28500 23118
rect 28448 23054 28500 23060
rect 29000 23112 29052 23118
rect 29000 23054 29052 23060
rect 28460 22778 28488 23054
rect 28448 22772 28500 22778
rect 28448 22714 28500 22720
rect 29656 22710 29684 23462
rect 29644 22704 29696 22710
rect 29644 22646 29696 22652
rect 28632 22228 28684 22234
rect 28632 22170 28684 22176
rect 28644 22098 28672 22170
rect 29932 22098 29960 23666
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 28632 22092 28684 22098
rect 28632 22034 28684 22040
rect 29920 22092 29972 22098
rect 29920 22034 29972 22040
rect 28724 22024 28776 22030
rect 28368 21950 28488 21978
rect 28724 21966 28776 21972
rect 28356 21888 28408 21894
rect 28356 21830 28408 21836
rect 28368 21554 28396 21830
rect 28356 21548 28408 21554
rect 28356 21490 28408 21496
rect 28356 21004 28408 21010
rect 28356 20946 28408 20952
rect 28368 20516 28396 20946
rect 28460 20618 28488 21950
rect 28736 21146 28764 21966
rect 28816 21480 28868 21486
rect 28816 21422 28868 21428
rect 28724 21140 28776 21146
rect 28724 21082 28776 21088
rect 28460 20590 28764 20618
rect 28368 20488 28488 20516
rect 28356 20392 28408 20398
rect 28356 20334 28408 20340
rect 28368 18222 28396 20334
rect 28356 18216 28408 18222
rect 28356 18158 28408 18164
rect 28264 18080 28316 18086
rect 28264 18022 28316 18028
rect 28172 17604 28224 17610
rect 28172 17546 28224 17552
rect 28080 16992 28132 16998
rect 28080 16934 28132 16940
rect 27988 16448 28040 16454
rect 27988 16390 28040 16396
rect 27896 15564 27948 15570
rect 27896 15506 27948 15512
rect 27908 15162 27936 15506
rect 28092 15502 28120 16934
rect 28172 16516 28224 16522
rect 28172 16458 28224 16464
rect 28184 16250 28212 16458
rect 28172 16244 28224 16250
rect 28172 16186 28224 16192
rect 28080 15496 28132 15502
rect 28080 15438 28132 15444
rect 27896 15156 27948 15162
rect 27896 15098 27948 15104
rect 27908 13376 27936 15098
rect 28080 14612 28132 14618
rect 28080 14554 28132 14560
rect 27908 13348 28028 13376
rect 27816 13280 27936 13308
rect 27724 13144 27844 13172
rect 27712 12844 27764 12850
rect 27712 12786 27764 12792
rect 27724 11898 27752 12786
rect 27712 11892 27764 11898
rect 27712 11834 27764 11840
rect 27620 11144 27672 11150
rect 27620 11086 27672 11092
rect 27712 10668 27764 10674
rect 27712 10610 27764 10616
rect 27620 10464 27672 10470
rect 27620 10406 27672 10412
rect 27632 9217 27660 10406
rect 27618 9208 27674 9217
rect 27618 9143 27674 9152
rect 27264 8588 27568 8616
rect 27158 8392 27214 8401
rect 27158 8327 27214 8336
rect 27068 7404 27120 7410
rect 27068 7346 27120 7352
rect 27080 6322 27108 7346
rect 27068 6316 27120 6322
rect 27068 6258 27120 6264
rect 26988 5596 27108 5624
rect 26792 4616 26844 4622
rect 26792 4558 26844 4564
rect 26976 4072 27028 4078
rect 26976 4014 27028 4020
rect 26988 3602 27016 4014
rect 26884 3596 26936 3602
rect 26884 3538 26936 3544
rect 26976 3596 27028 3602
rect 26976 3538 27028 3544
rect 26896 3058 26924 3538
rect 26884 3052 26936 3058
rect 26884 2994 26936 3000
rect 26516 2440 26568 2446
rect 26516 2382 26568 2388
rect 27080 1578 27108 5596
rect 27172 2774 27200 8327
rect 27264 6769 27292 8588
rect 27724 8537 27752 10610
rect 27816 8974 27844 13144
rect 27908 9586 27936 13280
rect 28000 12238 28028 13348
rect 28092 12374 28120 14554
rect 28276 13462 28304 18022
rect 28356 16788 28408 16794
rect 28356 16730 28408 16736
rect 28368 16114 28396 16730
rect 28356 16108 28408 16114
rect 28356 16050 28408 16056
rect 28460 15570 28488 20488
rect 28540 18760 28592 18766
rect 28540 18702 28592 18708
rect 28552 17542 28580 18702
rect 28632 18692 28684 18698
rect 28632 18634 28684 18640
rect 28644 18086 28672 18634
rect 28632 18080 28684 18086
rect 28632 18022 28684 18028
rect 28540 17536 28592 17542
rect 28540 17478 28592 17484
rect 28644 17354 28672 18022
rect 28552 17326 28672 17354
rect 28552 15910 28580 17326
rect 28736 16590 28764 20590
rect 28828 20330 28856 21422
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 28816 20324 28868 20330
rect 28816 20266 28868 20272
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 28724 16584 28776 16590
rect 28724 16526 28776 16532
rect 28632 16448 28684 16454
rect 28632 16390 28684 16396
rect 28644 16114 28672 16390
rect 28632 16108 28684 16114
rect 28632 16050 28684 16056
rect 28540 15904 28592 15910
rect 28540 15846 28592 15852
rect 28552 15638 28580 15846
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 28540 15632 28592 15638
rect 28540 15574 28592 15580
rect 28448 15564 28500 15570
rect 28448 15506 28500 15512
rect 28356 15360 28408 15366
rect 28356 15302 28408 15308
rect 28368 14414 28396 15302
rect 28460 14618 28488 15506
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 28448 14612 28500 14618
rect 28448 14554 28500 14560
rect 28356 14408 28408 14414
rect 28356 14350 28408 14356
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 28264 13456 28316 13462
rect 28264 13398 28316 13404
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 28080 12368 28132 12374
rect 28080 12310 28132 12316
rect 27988 12232 28040 12238
rect 27988 12174 28040 12180
rect 28080 12164 28132 12170
rect 28080 12106 28132 12112
rect 28264 12164 28316 12170
rect 28264 12106 28316 12112
rect 28092 11762 28120 12106
rect 28276 11898 28304 12106
rect 28448 12096 28500 12102
rect 28448 12038 28500 12044
rect 28264 11892 28316 11898
rect 28264 11834 28316 11840
rect 28080 11756 28132 11762
rect 28080 11698 28132 11704
rect 27988 10260 28040 10266
rect 27988 10202 28040 10208
rect 28000 9654 28028 10202
rect 27988 9648 28040 9654
rect 27988 9590 28040 9596
rect 27896 9580 27948 9586
rect 27896 9522 27948 9528
rect 27804 8968 27856 8974
rect 27804 8910 27856 8916
rect 27710 8528 27766 8537
rect 27436 8492 27488 8498
rect 27710 8463 27766 8472
rect 27436 8434 27488 8440
rect 27448 8090 27476 8434
rect 27436 8084 27488 8090
rect 27436 8026 27488 8032
rect 27620 8016 27672 8022
rect 27540 7964 27620 7970
rect 27540 7958 27672 7964
rect 27344 7948 27396 7954
rect 27344 7890 27396 7896
rect 27540 7942 27660 7958
rect 27356 7546 27384 7890
rect 27540 7886 27568 7942
rect 27528 7880 27580 7886
rect 27528 7822 27580 7828
rect 27620 7880 27672 7886
rect 27620 7822 27672 7828
rect 27344 7540 27396 7546
rect 27344 7482 27396 7488
rect 27250 6760 27306 6769
rect 27250 6695 27306 6704
rect 27264 6118 27292 6695
rect 27528 6316 27580 6322
rect 27632 6304 27660 7822
rect 27580 6276 27660 6304
rect 27528 6258 27580 6264
rect 27252 6112 27304 6118
rect 27252 6054 27304 6060
rect 27804 6112 27856 6118
rect 27804 6054 27856 6060
rect 27712 5704 27764 5710
rect 27712 5646 27764 5652
rect 27344 5228 27396 5234
rect 27344 5170 27396 5176
rect 27356 3738 27384 5170
rect 27724 5166 27752 5646
rect 27712 5160 27764 5166
rect 27712 5102 27764 5108
rect 27620 5024 27672 5030
rect 27620 4966 27672 4972
rect 27632 4690 27660 4966
rect 27620 4684 27672 4690
rect 27620 4626 27672 4632
rect 27724 4622 27752 5102
rect 27712 4616 27764 4622
rect 27712 4558 27764 4564
rect 27620 4480 27672 4486
rect 27620 4422 27672 4428
rect 27632 4146 27660 4422
rect 27620 4140 27672 4146
rect 27620 4082 27672 4088
rect 27344 3732 27396 3738
rect 27344 3674 27396 3680
rect 27528 3732 27580 3738
rect 27528 3674 27580 3680
rect 27540 3398 27568 3674
rect 27528 3392 27580 3398
rect 27528 3334 27580 3340
rect 27816 3194 27844 6054
rect 27896 5364 27948 5370
rect 27896 5306 27948 5312
rect 27804 3188 27856 3194
rect 27804 3130 27856 3136
rect 27172 2746 27476 2774
rect 26988 1550 27108 1578
rect 26712 870 26832 898
rect 26712 800 26740 870
rect 22296 734 22508 762
rect 22558 0 22614 800
rect 22926 0 22982 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 25226 0 25282 800
rect 25594 0 25650 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26698 0 26754 800
rect 26804 762 26832 870
rect 26988 762 27016 1550
rect 27068 1420 27120 1426
rect 27068 1362 27120 1368
rect 27080 800 27108 1362
rect 27448 800 27476 2746
rect 27908 2650 27936 5306
rect 28000 3126 28028 9590
rect 28092 9586 28120 11698
rect 28460 11150 28488 12038
rect 28998 11792 29054 11801
rect 28998 11727 29000 11736
rect 29052 11727 29054 11736
rect 29000 11698 29052 11704
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 29552 11280 29604 11286
rect 29552 11222 29604 11228
rect 28448 11144 28500 11150
rect 28448 11086 28500 11092
rect 29000 10736 29052 10742
rect 28920 10684 29000 10690
rect 28920 10678 29052 10684
rect 28448 10668 28500 10674
rect 28448 10610 28500 10616
rect 28920 10662 29040 10678
rect 28460 10441 28488 10610
rect 28632 10600 28684 10606
rect 28632 10542 28684 10548
rect 28722 10568 28778 10577
rect 28446 10432 28502 10441
rect 28446 10367 28502 10376
rect 28080 9580 28132 9586
rect 28080 9522 28132 9528
rect 28092 8974 28120 9522
rect 28080 8968 28132 8974
rect 28080 8910 28132 8916
rect 28356 8968 28408 8974
rect 28356 8910 28408 8916
rect 28092 7818 28120 8910
rect 28172 8900 28224 8906
rect 28172 8842 28224 8848
rect 28184 8634 28212 8842
rect 28368 8634 28396 8910
rect 28172 8628 28224 8634
rect 28172 8570 28224 8576
rect 28356 8628 28408 8634
rect 28356 8570 28408 8576
rect 28184 8514 28212 8570
rect 28184 8486 28396 8514
rect 28368 8430 28396 8486
rect 28356 8424 28408 8430
rect 28356 8366 28408 8372
rect 28264 8288 28316 8294
rect 28262 8256 28264 8265
rect 28316 8256 28318 8265
rect 28262 8191 28318 8200
rect 28460 7970 28488 10367
rect 28644 9586 28672 10542
rect 28722 10503 28724 10512
rect 28776 10503 28778 10512
rect 28816 10532 28868 10538
rect 28724 10474 28776 10480
rect 28816 10474 28868 10480
rect 28724 10124 28776 10130
rect 28724 10066 28776 10072
rect 28632 9580 28684 9586
rect 28632 9522 28684 9528
rect 28644 8974 28672 9522
rect 28632 8968 28684 8974
rect 28632 8910 28684 8916
rect 28644 8022 28672 8910
rect 28368 7942 28488 7970
rect 28632 8016 28684 8022
rect 28632 7958 28684 7964
rect 28368 7834 28396 7942
rect 28276 7818 28396 7834
rect 28080 7812 28132 7818
rect 28080 7754 28132 7760
rect 28264 7812 28396 7818
rect 28316 7806 28396 7812
rect 28264 7754 28316 7760
rect 28080 7472 28132 7478
rect 28080 7414 28132 7420
rect 28092 7342 28120 7414
rect 28080 7336 28132 7342
rect 28080 7278 28132 7284
rect 28080 6792 28132 6798
rect 28080 6734 28132 6740
rect 28092 4078 28120 6734
rect 28276 5778 28304 7754
rect 28736 6984 28764 10066
rect 28460 6956 28764 6984
rect 28354 5808 28410 5817
rect 28264 5772 28316 5778
rect 28354 5743 28356 5752
rect 28264 5714 28316 5720
rect 28408 5743 28410 5752
rect 28356 5714 28408 5720
rect 28460 4826 28488 6956
rect 28540 6724 28592 6730
rect 28540 6666 28592 6672
rect 28552 6118 28580 6666
rect 28540 6112 28592 6118
rect 28540 6054 28592 6060
rect 28448 4820 28500 4826
rect 28448 4762 28500 4768
rect 28356 4480 28408 4486
rect 28356 4422 28408 4428
rect 28448 4480 28500 4486
rect 28448 4422 28500 4428
rect 28080 4072 28132 4078
rect 28080 4014 28132 4020
rect 28368 3942 28396 4422
rect 28356 3936 28408 3942
rect 28356 3878 28408 3884
rect 28080 3188 28132 3194
rect 28080 3130 28132 3136
rect 27988 3120 28040 3126
rect 27988 3062 28040 3068
rect 28092 2922 28120 3130
rect 28080 2916 28132 2922
rect 28080 2858 28132 2864
rect 27896 2644 27948 2650
rect 27896 2586 27948 2592
rect 27804 2576 27856 2582
rect 27804 2518 27856 2524
rect 27816 800 27844 2518
rect 28092 2446 28120 2858
rect 28080 2440 28132 2446
rect 28080 2382 28132 2388
rect 28368 2378 28396 3878
rect 28460 3466 28488 4422
rect 28448 3460 28500 3466
rect 28448 3402 28500 3408
rect 28552 3126 28580 6054
rect 28724 5160 28776 5166
rect 28828 5137 28856 10474
rect 28920 10266 28948 10662
rect 29368 10464 29420 10470
rect 29368 10406 29420 10412
rect 28908 10260 28960 10266
rect 28908 10202 28960 10208
rect 29184 10192 29236 10198
rect 29182 10160 29184 10169
rect 29236 10160 29238 10169
rect 29182 10095 29238 10104
rect 29380 10062 29408 10406
rect 29368 10056 29420 10062
rect 29368 9998 29420 10004
rect 29000 9920 29052 9926
rect 29000 9862 29052 9868
rect 29012 9654 29040 9862
rect 29000 9648 29052 9654
rect 29000 9590 29052 9596
rect 29276 9580 29328 9586
rect 29276 9522 29328 9528
rect 29368 9580 29420 9586
rect 29368 9522 29420 9528
rect 29184 9036 29236 9042
rect 29184 8978 29236 8984
rect 29196 8634 29224 8978
rect 29184 8628 29236 8634
rect 29184 8570 29236 8576
rect 29092 8084 29144 8090
rect 29092 8026 29144 8032
rect 29000 8016 29052 8022
rect 29000 7958 29052 7964
rect 28908 7744 28960 7750
rect 28908 7686 28960 7692
rect 28920 7342 28948 7686
rect 28908 7336 28960 7342
rect 28908 7278 28960 7284
rect 29012 6322 29040 7958
rect 29104 6866 29132 8026
rect 29288 7954 29316 9522
rect 29276 7948 29328 7954
rect 29276 7890 29328 7896
rect 29182 7848 29238 7857
rect 29182 7783 29238 7792
rect 29196 7410 29224 7783
rect 29276 7540 29328 7546
rect 29276 7482 29328 7488
rect 29184 7404 29236 7410
rect 29184 7346 29236 7352
rect 29184 7200 29236 7206
rect 29184 7142 29236 7148
rect 29196 7002 29224 7142
rect 29184 6996 29236 7002
rect 29184 6938 29236 6944
rect 29092 6860 29144 6866
rect 29092 6802 29144 6808
rect 29196 6746 29224 6938
rect 29288 6798 29316 7482
rect 29104 6718 29224 6746
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 29000 6316 29052 6322
rect 29000 6258 29052 6264
rect 29000 5840 29052 5846
rect 29000 5782 29052 5788
rect 28908 5568 28960 5574
rect 28908 5510 28960 5516
rect 28724 5102 28776 5108
rect 28814 5128 28870 5137
rect 28736 4622 28764 5102
rect 28814 5063 28870 5072
rect 28920 4706 28948 5510
rect 29012 5302 29040 5782
rect 29000 5296 29052 5302
rect 29000 5238 29052 5244
rect 29104 5030 29132 6718
rect 29288 5846 29316 6734
rect 29276 5840 29328 5846
rect 29276 5782 29328 5788
rect 29380 5624 29408 9522
rect 29460 7948 29512 7954
rect 29460 7890 29512 7896
rect 29472 6934 29500 7890
rect 29460 6928 29512 6934
rect 29460 6870 29512 6876
rect 29460 6112 29512 6118
rect 29460 6054 29512 6060
rect 29196 5596 29408 5624
rect 29092 5024 29144 5030
rect 29092 4966 29144 4972
rect 28920 4678 29132 4706
rect 28724 4616 28776 4622
rect 28724 4558 28776 4564
rect 28816 4480 28868 4486
rect 28816 4422 28868 4428
rect 28724 4072 28776 4078
rect 28724 4014 28776 4020
rect 28540 3120 28592 3126
rect 28540 3062 28592 3068
rect 28540 2916 28592 2922
rect 28540 2858 28592 2864
rect 28356 2372 28408 2378
rect 28356 2314 28408 2320
rect 28552 800 28580 2858
rect 28736 2854 28764 4014
rect 28828 3398 28856 4422
rect 28816 3392 28868 3398
rect 28816 3334 28868 3340
rect 28828 3126 28856 3334
rect 28920 3194 28948 4678
rect 29000 4616 29052 4622
rect 29000 4558 29052 4564
rect 29012 4078 29040 4558
rect 29104 4486 29132 4678
rect 29092 4480 29144 4486
rect 29092 4422 29144 4428
rect 29000 4072 29052 4078
rect 29000 4014 29052 4020
rect 28908 3188 28960 3194
rect 28908 3130 28960 3136
rect 28816 3120 28868 3126
rect 28816 3062 28868 3068
rect 29196 2990 29224 5596
rect 29472 5370 29500 6054
rect 29564 5778 29592 11222
rect 29736 11144 29788 11150
rect 29734 11112 29736 11121
rect 29788 11112 29790 11121
rect 29734 11047 29790 11056
rect 36280 11014 36308 46854
rect 36268 11008 36320 11014
rect 36268 10950 36320 10956
rect 30196 10668 30248 10674
rect 30196 10610 30248 10616
rect 30288 10668 30340 10674
rect 30288 10610 30340 10616
rect 29736 10056 29788 10062
rect 30208 10033 30236 10610
rect 29736 9998 29788 10004
rect 30194 10024 30250 10033
rect 29748 9761 29776 9998
rect 30194 9959 30250 9968
rect 30104 9920 30156 9926
rect 30104 9862 30156 9868
rect 29734 9752 29790 9761
rect 29734 9687 29790 9696
rect 29920 8900 29972 8906
rect 29920 8842 29972 8848
rect 29736 8832 29788 8838
rect 29736 8774 29788 8780
rect 29748 8634 29776 8774
rect 29736 8628 29788 8634
rect 29736 8570 29788 8576
rect 29828 8492 29880 8498
rect 29828 8434 29880 8440
rect 29840 7818 29868 8434
rect 29828 7812 29880 7818
rect 29828 7754 29880 7760
rect 29932 6882 29960 8842
rect 30012 8356 30064 8362
rect 30012 8298 30064 8304
rect 29656 6854 29960 6882
rect 29552 5772 29604 5778
rect 29552 5714 29604 5720
rect 29460 5364 29512 5370
rect 29460 5306 29512 5312
rect 29276 5228 29328 5234
rect 29276 5170 29328 5176
rect 29184 2984 29236 2990
rect 29184 2926 29236 2932
rect 28632 2848 28684 2854
rect 28632 2790 28684 2796
rect 28724 2848 28776 2854
rect 28724 2790 28776 2796
rect 28908 2848 28960 2854
rect 28908 2790 28960 2796
rect 28644 2650 28672 2790
rect 28920 2650 28948 2790
rect 28632 2644 28684 2650
rect 28632 2586 28684 2592
rect 28908 2644 28960 2650
rect 28908 2586 28960 2592
rect 29288 2514 29316 5170
rect 29472 4554 29500 5306
rect 29552 5024 29604 5030
rect 29552 4966 29604 4972
rect 29460 4548 29512 4554
rect 29460 4490 29512 4496
rect 29460 4140 29512 4146
rect 29460 4082 29512 4088
rect 29368 3392 29420 3398
rect 29368 3334 29420 3340
rect 29276 2508 29328 2514
rect 29276 2450 29328 2456
rect 28816 2304 28868 2310
rect 28816 2246 28868 2252
rect 28828 1426 28856 2246
rect 28816 1420 28868 1426
rect 28816 1362 28868 1368
rect 29380 800 29408 3334
rect 29472 2854 29500 4082
rect 29460 2848 29512 2854
rect 29460 2790 29512 2796
rect 29564 2446 29592 4966
rect 29656 3058 29684 6854
rect 29736 6792 29788 6798
rect 29736 6734 29788 6740
rect 29748 6390 29776 6734
rect 30024 6730 30052 8298
rect 29828 6724 29880 6730
rect 30012 6724 30064 6730
rect 29880 6684 29960 6712
rect 29828 6666 29880 6672
rect 29736 6384 29788 6390
rect 29736 6326 29788 6332
rect 29828 6384 29880 6390
rect 29828 6326 29880 6332
rect 29734 5808 29790 5817
rect 29734 5743 29790 5752
rect 29748 5710 29776 5743
rect 29736 5704 29788 5710
rect 29736 5646 29788 5652
rect 29736 5024 29788 5030
rect 29736 4966 29788 4972
rect 29748 4826 29776 4966
rect 29736 4820 29788 4826
rect 29736 4762 29788 4768
rect 29748 4146 29776 4762
rect 29736 4140 29788 4146
rect 29736 4082 29788 4088
rect 29736 3528 29788 3534
rect 29736 3470 29788 3476
rect 29748 3058 29776 3470
rect 29644 3052 29696 3058
rect 29644 2994 29696 3000
rect 29736 3052 29788 3058
rect 29736 2994 29788 3000
rect 29552 2440 29604 2446
rect 29552 2382 29604 2388
rect 29840 2378 29868 6326
rect 29932 2514 29960 6684
rect 30012 6666 30064 6672
rect 30116 5692 30144 9862
rect 30196 8968 30248 8974
rect 30196 8910 30248 8916
rect 30208 7342 30236 8910
rect 30196 7336 30248 7342
rect 30196 7278 30248 7284
rect 30116 5664 30236 5692
rect 30012 5568 30064 5574
rect 30012 5510 30064 5516
rect 30024 4214 30052 5510
rect 30208 5250 30236 5664
rect 30300 5574 30328 10610
rect 30656 10464 30708 10470
rect 30656 10406 30708 10412
rect 30668 9761 30696 10406
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 31024 9920 31076 9926
rect 31022 9888 31024 9897
rect 31076 9888 31078 9897
rect 31022 9823 31078 9832
rect 30654 9752 30710 9761
rect 30654 9687 30710 9696
rect 32496 9716 32548 9722
rect 32496 9658 32548 9664
rect 30932 9580 30984 9586
rect 30932 9522 30984 9528
rect 31208 9580 31260 9586
rect 31208 9522 31260 9528
rect 30748 9376 30800 9382
rect 30748 9318 30800 9324
rect 30656 8968 30708 8974
rect 30656 8910 30708 8916
rect 30564 8832 30616 8838
rect 30564 8774 30616 8780
rect 30472 7880 30524 7886
rect 30472 7822 30524 7828
rect 30380 7744 30432 7750
rect 30380 7686 30432 7692
rect 30392 6322 30420 7686
rect 30484 6662 30512 7822
rect 30472 6656 30524 6662
rect 30472 6598 30524 6604
rect 30380 6316 30432 6322
rect 30380 6258 30432 6264
rect 30380 5636 30432 5642
rect 30380 5578 30432 5584
rect 30288 5568 30340 5574
rect 30288 5510 30340 5516
rect 30392 5370 30420 5578
rect 30380 5364 30432 5370
rect 30380 5306 30432 5312
rect 30116 5222 30236 5250
rect 30288 5228 30340 5234
rect 30012 4208 30064 4214
rect 30012 4150 30064 4156
rect 30116 4026 30144 5222
rect 30288 5170 30340 5176
rect 30196 5160 30248 5166
rect 30196 5102 30248 5108
rect 30208 4078 30236 5102
rect 30300 4146 30328 5170
rect 30576 4826 30604 8774
rect 30564 4820 30616 4826
rect 30564 4762 30616 4768
rect 30380 4480 30432 4486
rect 30380 4422 30432 4428
rect 30288 4140 30340 4146
rect 30288 4082 30340 4088
rect 30024 3998 30144 4026
rect 30196 4072 30248 4078
rect 30196 4014 30248 4020
rect 30024 3738 30052 3998
rect 30104 3936 30156 3942
rect 30104 3878 30156 3884
rect 30012 3732 30064 3738
rect 30012 3674 30064 3680
rect 30116 3466 30144 3878
rect 30104 3460 30156 3466
rect 30104 3402 30156 3408
rect 29920 2508 29972 2514
rect 29920 2450 29972 2456
rect 30392 2446 30420 4422
rect 30472 4140 30524 4146
rect 30472 4082 30524 4088
rect 30484 3738 30512 4082
rect 30668 4010 30696 8910
rect 30760 5914 30788 9318
rect 30840 8492 30892 8498
rect 30840 8434 30892 8440
rect 30852 7546 30880 8434
rect 30840 7540 30892 7546
rect 30840 7482 30892 7488
rect 30748 5908 30800 5914
rect 30748 5850 30800 5856
rect 30944 5681 30972 9522
rect 31220 9081 31248 9522
rect 31206 9072 31262 9081
rect 31206 9007 31262 9016
rect 31208 8968 31260 8974
rect 31208 8910 31260 8916
rect 31852 8968 31904 8974
rect 31852 8910 31904 8916
rect 31220 8401 31248 8910
rect 31206 8392 31262 8401
rect 31206 8327 31262 8336
rect 31024 7880 31076 7886
rect 31024 7822 31076 7828
rect 31668 7880 31720 7886
rect 31668 7822 31720 7828
rect 30930 5672 30986 5681
rect 30930 5607 30986 5616
rect 31036 5098 31064 7822
rect 31208 7404 31260 7410
rect 31208 7346 31260 7352
rect 31220 6662 31248 7346
rect 31208 6656 31260 6662
rect 31208 6598 31260 6604
rect 31024 5092 31076 5098
rect 31024 5034 31076 5040
rect 31220 4554 31248 6598
rect 31680 6089 31708 7822
rect 31760 6792 31812 6798
rect 31760 6734 31812 6740
rect 31666 6080 31722 6089
rect 31666 6015 31722 6024
rect 31576 5568 31628 5574
rect 31628 5528 31708 5556
rect 31576 5510 31628 5516
rect 31588 5302 31616 5510
rect 31576 5296 31628 5302
rect 31576 5238 31628 5244
rect 31392 5024 31444 5030
rect 31392 4966 31444 4972
rect 31404 4826 31432 4966
rect 31392 4820 31444 4826
rect 31392 4762 31444 4768
rect 31680 4554 31708 5528
rect 31772 4826 31800 6734
rect 31864 6458 31892 8910
rect 32404 8356 32456 8362
rect 32404 8298 32456 8304
rect 31944 7268 31996 7274
rect 31944 7210 31996 7216
rect 31852 6452 31904 6458
rect 31852 6394 31904 6400
rect 31852 6112 31904 6118
rect 31852 6054 31904 6060
rect 31760 4820 31812 4826
rect 31760 4762 31812 4768
rect 31208 4548 31260 4554
rect 31208 4490 31260 4496
rect 31668 4548 31720 4554
rect 31668 4490 31720 4496
rect 31392 4140 31444 4146
rect 31392 4082 31444 4088
rect 30656 4004 30708 4010
rect 30656 3946 30708 3952
rect 31024 3936 31076 3942
rect 31024 3878 31076 3884
rect 30472 3732 30524 3738
rect 30472 3674 30524 3680
rect 30484 3466 30512 3674
rect 30748 3596 30800 3602
rect 30748 3538 30800 3544
rect 30472 3460 30524 3466
rect 30472 3402 30524 3408
rect 30760 3194 30788 3538
rect 30748 3188 30800 3194
rect 30748 3130 30800 3136
rect 31036 3126 31064 3878
rect 31300 3392 31352 3398
rect 31300 3334 31352 3340
rect 31024 3120 31076 3126
rect 31024 3062 31076 3068
rect 31312 3058 31340 3334
rect 31404 3194 31432 4082
rect 31392 3188 31444 3194
rect 31392 3130 31444 3136
rect 30840 3052 30892 3058
rect 30840 2994 30892 3000
rect 31300 3052 31352 3058
rect 31300 2994 31352 3000
rect 31760 3052 31812 3058
rect 31760 2994 31812 3000
rect 30748 2848 30800 2854
rect 30748 2790 30800 2796
rect 30760 2650 30788 2790
rect 30748 2644 30800 2650
rect 30748 2586 30800 2592
rect 30380 2440 30432 2446
rect 30380 2382 30432 2388
rect 29828 2372 29880 2378
rect 29828 2314 29880 2320
rect 30104 2372 30156 2378
rect 30104 2314 30156 2320
rect 30116 800 30144 2314
rect 30852 800 30880 2994
rect 31576 2848 31628 2854
rect 31576 2790 31628 2796
rect 31588 800 31616 2790
rect 31772 2310 31800 2994
rect 31864 2774 31892 6054
rect 31956 5778 31984 7210
rect 32128 7200 32180 7206
rect 32128 7142 32180 7148
rect 32140 6882 32168 7142
rect 32140 6854 32260 6882
rect 32128 6724 32180 6730
rect 32128 6666 32180 6672
rect 32140 6254 32168 6666
rect 32128 6248 32180 6254
rect 32128 6190 32180 6196
rect 31944 5772 31996 5778
rect 31944 5714 31996 5720
rect 32036 5772 32088 5778
rect 32036 5714 32088 5720
rect 32048 3738 32076 5714
rect 32140 5642 32168 6190
rect 32128 5636 32180 5642
rect 32128 5578 32180 5584
rect 32140 3942 32168 5578
rect 32232 5030 32260 6854
rect 32312 6792 32364 6798
rect 32312 6734 32364 6740
rect 32324 5778 32352 6734
rect 32416 6322 32444 8298
rect 32508 7410 32536 9658
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 32772 9172 32824 9178
rect 32772 9114 32824 9120
rect 32680 8628 32732 8634
rect 32680 8570 32732 8576
rect 32496 7404 32548 7410
rect 32496 7346 32548 7352
rect 32508 6866 32536 7346
rect 32496 6860 32548 6866
rect 32496 6802 32548 6808
rect 32404 6316 32456 6322
rect 32404 6258 32456 6264
rect 32312 5772 32364 5778
rect 32312 5714 32364 5720
rect 32404 5636 32456 5642
rect 32404 5578 32456 5584
rect 32220 5024 32272 5030
rect 32220 4966 32272 4972
rect 32232 4826 32260 4966
rect 32220 4820 32272 4826
rect 32272 4780 32352 4808
rect 32220 4762 32272 4768
rect 32220 4480 32272 4486
rect 32220 4422 32272 4428
rect 32128 3936 32180 3942
rect 32128 3878 32180 3884
rect 32036 3732 32088 3738
rect 32036 3674 32088 3680
rect 32140 3534 32168 3878
rect 32128 3528 32180 3534
rect 32128 3470 32180 3476
rect 32232 3398 32260 4422
rect 32324 3670 32352 4780
rect 32312 3664 32364 3670
rect 32312 3606 32364 3612
rect 32416 3466 32444 5578
rect 32508 5302 32536 6802
rect 32496 5296 32548 5302
rect 32496 5238 32548 5244
rect 32692 4146 32720 8570
rect 32784 7478 32812 9114
rect 33140 8492 33192 8498
rect 33140 8434 33192 8440
rect 34704 8492 34756 8498
rect 34704 8434 34756 8440
rect 32956 8424 33008 8430
rect 32956 8366 33008 8372
rect 32968 7886 32996 8366
rect 32956 7880 33008 7886
rect 32956 7822 33008 7828
rect 32864 7812 32916 7818
rect 32864 7754 32916 7760
rect 32876 7546 32904 7754
rect 32864 7540 32916 7546
rect 32864 7482 32916 7488
rect 32772 7472 32824 7478
rect 32772 7414 32824 7420
rect 32968 7342 32996 7822
rect 33048 7744 33100 7750
rect 33048 7686 33100 7692
rect 33060 7410 33088 7686
rect 33048 7404 33100 7410
rect 33048 7346 33100 7352
rect 32956 7336 33008 7342
rect 32956 7278 33008 7284
rect 32772 6792 32824 6798
rect 32772 6734 32824 6740
rect 32784 5817 32812 6734
rect 32864 6656 32916 6662
rect 32864 6598 32916 6604
rect 32770 5808 32826 5817
rect 32770 5743 32826 5752
rect 32784 5234 32812 5743
rect 32772 5228 32824 5234
rect 32772 5170 32824 5176
rect 32784 4593 32812 5170
rect 32770 4584 32826 4593
rect 32770 4519 32826 4528
rect 32680 4140 32732 4146
rect 32680 4082 32732 4088
rect 32404 3460 32456 3466
rect 32404 3402 32456 3408
rect 32220 3392 32272 3398
rect 32220 3334 32272 3340
rect 32876 3058 32904 6598
rect 32968 6390 32996 7278
rect 32956 6384 33008 6390
rect 32956 6326 33008 6332
rect 33048 6112 33100 6118
rect 33048 6054 33100 6060
rect 33060 5642 33088 6054
rect 33048 5636 33100 5642
rect 33048 5578 33100 5584
rect 32956 5568 33008 5574
rect 32956 5510 33008 5516
rect 32968 4486 32996 5510
rect 33152 4826 33180 8434
rect 33600 8356 33652 8362
rect 33600 8298 33652 8304
rect 33416 7200 33468 7206
rect 33416 7142 33468 7148
rect 33428 5914 33456 7142
rect 33508 6724 33560 6730
rect 33508 6666 33560 6672
rect 33416 5908 33468 5914
rect 33416 5850 33468 5856
rect 33428 5386 33456 5850
rect 33244 5358 33456 5386
rect 33048 4820 33100 4826
rect 33048 4762 33100 4768
rect 33140 4820 33192 4826
rect 33140 4762 33192 4768
rect 33060 4706 33088 4762
rect 33244 4706 33272 5358
rect 33416 5228 33468 5234
rect 33416 5170 33468 5176
rect 33324 5024 33376 5030
rect 33324 4966 33376 4972
rect 33060 4678 33272 4706
rect 32956 4480 33008 4486
rect 32956 4422 33008 4428
rect 33232 4480 33284 4486
rect 33232 4422 33284 4428
rect 32864 3052 32916 3058
rect 32864 2994 32916 3000
rect 32312 2984 32364 2990
rect 32312 2926 32364 2932
rect 32324 2854 32352 2926
rect 32312 2848 32364 2854
rect 32312 2790 32364 2796
rect 31864 2746 32076 2774
rect 32048 2446 32076 2746
rect 32312 2576 32364 2582
rect 32312 2518 32364 2524
rect 32036 2440 32088 2446
rect 32036 2382 32088 2388
rect 31760 2304 31812 2310
rect 31760 2246 31812 2252
rect 32324 800 32352 2518
rect 33244 2446 33272 4422
rect 33336 2990 33364 4966
rect 33428 3602 33456 5170
rect 33520 4706 33548 6666
rect 33612 5914 33640 8298
rect 34716 8090 34744 8434
rect 35440 8288 35492 8294
rect 35440 8230 35492 8236
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34704 8084 34756 8090
rect 34704 8026 34756 8032
rect 35164 7880 35216 7886
rect 35164 7822 35216 7828
rect 34704 7744 34756 7750
rect 34704 7686 34756 7692
rect 34716 7546 34744 7686
rect 34704 7540 34756 7546
rect 34704 7482 34756 7488
rect 34612 6996 34664 7002
rect 34612 6938 34664 6944
rect 34060 6792 34112 6798
rect 34060 6734 34112 6740
rect 33876 6656 33928 6662
rect 33876 6598 33928 6604
rect 33600 5908 33652 5914
rect 33600 5850 33652 5856
rect 33520 4678 33640 4706
rect 33508 4548 33560 4554
rect 33508 4490 33560 4496
rect 33520 4282 33548 4490
rect 33508 4276 33560 4282
rect 33508 4218 33560 4224
rect 33416 3596 33468 3602
rect 33416 3538 33468 3544
rect 33520 3534 33548 4218
rect 33508 3528 33560 3534
rect 33508 3470 33560 3476
rect 33324 2984 33376 2990
rect 33324 2926 33376 2932
rect 33612 2774 33640 4678
rect 33888 3194 33916 6598
rect 34072 5778 34100 6734
rect 34624 5914 34652 6938
rect 34716 6730 34744 7482
rect 35176 7410 35204 7822
rect 35452 7750 35480 8230
rect 35440 7744 35492 7750
rect 35440 7686 35492 7692
rect 35624 7744 35676 7750
rect 35624 7686 35676 7692
rect 36084 7744 36136 7750
rect 36084 7686 36136 7692
rect 35164 7404 35216 7410
rect 35164 7346 35216 7352
rect 35452 7290 35480 7686
rect 35636 7478 35664 7686
rect 36096 7546 36124 7686
rect 36084 7540 36136 7546
rect 36084 7482 36136 7488
rect 35624 7472 35676 7478
rect 35624 7414 35676 7420
rect 35716 7404 35768 7410
rect 35716 7346 35768 7352
rect 34796 7268 34848 7274
rect 35452 7262 35664 7290
rect 34796 7210 34848 7216
rect 34704 6724 34756 6730
rect 34704 6666 34756 6672
rect 34808 6390 34836 7210
rect 35440 7200 35492 7206
rect 35440 7142 35492 7148
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34888 6656 34940 6662
rect 34888 6598 34940 6604
rect 34796 6384 34848 6390
rect 34796 6326 34848 6332
rect 34900 6202 34928 6598
rect 34808 6174 34928 6202
rect 34612 5908 34664 5914
rect 34612 5850 34664 5856
rect 34428 5840 34480 5846
rect 34428 5782 34480 5788
rect 34060 5772 34112 5778
rect 34060 5714 34112 5720
rect 34152 5704 34204 5710
rect 34152 5646 34204 5652
rect 33968 4616 34020 4622
rect 33968 4558 34020 4564
rect 33980 3398 34008 4558
rect 33968 3392 34020 3398
rect 33968 3334 34020 3340
rect 34164 3194 34192 5646
rect 34440 5030 34468 5782
rect 34612 5636 34664 5642
rect 34612 5578 34664 5584
rect 34520 5568 34572 5574
rect 34520 5510 34572 5516
rect 34532 5370 34560 5510
rect 34520 5364 34572 5370
rect 34520 5306 34572 5312
rect 34624 5302 34652 5578
rect 34808 5574 34836 6174
rect 35348 6112 35400 6118
rect 35348 6054 35400 6060
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 35360 5642 35388 6054
rect 35348 5636 35400 5642
rect 35348 5578 35400 5584
rect 34796 5568 34848 5574
rect 34796 5510 34848 5516
rect 34612 5296 34664 5302
rect 34612 5238 34664 5244
rect 34520 5160 34572 5166
rect 34520 5102 34572 5108
rect 34428 5024 34480 5030
rect 34428 4966 34480 4972
rect 34440 4758 34468 4966
rect 34428 4752 34480 4758
rect 34428 4694 34480 4700
rect 34336 4548 34388 4554
rect 34336 4490 34388 4496
rect 34348 3398 34376 4490
rect 34428 4072 34480 4078
rect 34428 4014 34480 4020
rect 34440 3602 34468 4014
rect 34532 3738 34560 5102
rect 34624 4865 34652 5238
rect 34796 5228 34848 5234
rect 34796 5170 34848 5176
rect 35348 5228 35400 5234
rect 35348 5170 35400 5176
rect 34704 5092 34756 5098
rect 34704 5034 34756 5040
rect 34610 4856 34666 4865
rect 34610 4791 34666 4800
rect 34612 4752 34664 4758
rect 34612 4694 34664 4700
rect 34520 3732 34572 3738
rect 34520 3674 34572 3680
rect 34624 3670 34652 4694
rect 34612 3664 34664 3670
rect 34612 3606 34664 3612
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 34336 3392 34388 3398
rect 34336 3334 34388 3340
rect 33876 3188 33928 3194
rect 33876 3130 33928 3136
rect 34152 3188 34204 3194
rect 34152 3130 34204 3136
rect 33784 2916 33836 2922
rect 33784 2858 33836 2864
rect 33428 2746 33640 2774
rect 33428 2446 33456 2746
rect 33232 2440 33284 2446
rect 33232 2382 33284 2388
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 33140 2304 33192 2310
rect 33140 2246 33192 2252
rect 33152 1442 33180 2246
rect 33060 1414 33180 1442
rect 33060 800 33088 1414
rect 33796 800 33824 2858
rect 34612 2576 34664 2582
rect 34612 2518 34664 2524
rect 34624 800 34652 2518
rect 34716 2446 34744 5034
rect 34808 4282 34836 5170
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 35360 4758 35388 5170
rect 35348 4752 35400 4758
rect 34886 4720 34942 4729
rect 35348 4694 35400 4700
rect 34886 4655 34942 4664
rect 34900 4486 34928 4655
rect 34888 4480 34940 4486
rect 34888 4422 34940 4428
rect 34796 4276 34848 4282
rect 34796 4218 34848 4224
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 35452 3534 35480 7142
rect 35532 5568 35584 5574
rect 35532 5510 35584 5516
rect 35440 3528 35492 3534
rect 35440 3470 35492 3476
rect 35348 3392 35400 3398
rect 35348 3334 35400 3340
rect 35360 3126 35388 3334
rect 35348 3120 35400 3126
rect 35348 3062 35400 3068
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35544 2514 35572 5510
rect 35636 3466 35664 7262
rect 35728 4826 35756 7346
rect 35808 6792 35860 6798
rect 35808 6734 35860 6740
rect 35820 5914 35848 6734
rect 35900 6384 35952 6390
rect 35900 6326 35952 6332
rect 35808 5908 35860 5914
rect 35808 5850 35860 5856
rect 35808 5772 35860 5778
rect 35808 5714 35860 5720
rect 35716 4820 35768 4826
rect 35716 4762 35768 4768
rect 35820 4758 35848 5714
rect 35912 5302 35940 6326
rect 35992 6112 36044 6118
rect 35992 6054 36044 6060
rect 36004 5846 36032 6054
rect 35992 5840 36044 5846
rect 35992 5782 36044 5788
rect 35900 5296 35952 5302
rect 35900 5238 35952 5244
rect 35900 5024 35952 5030
rect 35900 4966 35952 4972
rect 35808 4752 35860 4758
rect 35808 4694 35860 4700
rect 35716 4616 35768 4622
rect 35714 4584 35716 4593
rect 35768 4584 35770 4593
rect 35714 4519 35770 4528
rect 35808 4276 35860 4282
rect 35808 4218 35860 4224
rect 35624 3460 35676 3466
rect 35624 3402 35676 3408
rect 35820 3126 35848 4218
rect 35808 3120 35860 3126
rect 35808 3062 35860 3068
rect 35532 2508 35584 2514
rect 35532 2450 35584 2456
rect 35912 2446 35940 4966
rect 36096 4214 36124 7482
rect 36452 7404 36504 7410
rect 36452 7346 36504 7352
rect 36464 6458 36492 7346
rect 37556 6860 37608 6866
rect 37556 6802 37608 6808
rect 36452 6452 36504 6458
rect 36452 6394 36504 6400
rect 37280 6316 37332 6322
rect 37280 6258 37332 6264
rect 36912 5704 36964 5710
rect 36912 5646 36964 5652
rect 37096 5704 37148 5710
rect 37096 5646 37148 5652
rect 36268 5228 36320 5234
rect 36268 5170 36320 5176
rect 36176 4480 36228 4486
rect 36176 4422 36228 4428
rect 36084 4208 36136 4214
rect 36084 4150 36136 4156
rect 36188 2922 36216 4422
rect 36280 3194 36308 5170
rect 36452 4480 36504 4486
rect 36452 4422 36504 4428
rect 36360 4208 36412 4214
rect 36360 4150 36412 4156
rect 36372 3398 36400 4150
rect 36464 3942 36492 4422
rect 36452 3936 36504 3942
rect 36452 3878 36504 3884
rect 36464 3738 36492 3878
rect 36924 3738 36952 5646
rect 36452 3732 36504 3738
rect 36452 3674 36504 3680
rect 36912 3732 36964 3738
rect 36912 3674 36964 3680
rect 36360 3392 36412 3398
rect 36360 3334 36412 3340
rect 36268 3188 36320 3194
rect 36268 3130 36320 3136
rect 36372 3126 36400 3334
rect 36360 3120 36412 3126
rect 36360 3062 36412 3068
rect 36176 2916 36228 2922
rect 36176 2858 36228 2864
rect 36464 2854 36492 3674
rect 37108 3194 37136 5646
rect 37292 5370 37320 6258
rect 37372 5840 37424 5846
rect 37372 5782 37424 5788
rect 37280 5364 37332 5370
rect 37280 5306 37332 5312
rect 37280 5024 37332 5030
rect 37280 4966 37332 4972
rect 37096 3188 37148 3194
rect 37096 3130 37148 3136
rect 36452 2848 36504 2854
rect 36452 2790 36504 2796
rect 36820 2848 36872 2854
rect 36820 2790 36872 2796
rect 36084 2576 36136 2582
rect 36084 2518 36136 2524
rect 34704 2440 34756 2446
rect 34704 2382 34756 2388
rect 35900 2440 35952 2446
rect 35900 2382 35952 2388
rect 35348 2372 35400 2378
rect 35348 2314 35400 2320
rect 35360 800 35388 2314
rect 36096 800 36124 2518
rect 36832 800 36860 2790
rect 37292 2446 37320 4966
rect 37384 3058 37412 5782
rect 37464 5568 37516 5574
rect 37464 5510 37516 5516
rect 37476 3534 37504 5510
rect 37568 4622 37596 6802
rect 37648 6656 37700 6662
rect 37648 6598 37700 6604
rect 37660 5234 37688 6598
rect 37924 6112 37976 6118
rect 37924 6054 37976 6060
rect 37740 5704 37792 5710
rect 37740 5646 37792 5652
rect 37648 5228 37700 5234
rect 37648 5170 37700 5176
rect 37556 4616 37608 4622
rect 37556 4558 37608 4564
rect 37752 4010 37780 5646
rect 37832 5568 37884 5574
rect 37832 5510 37884 5516
rect 37844 4146 37872 5510
rect 37832 4140 37884 4146
rect 37832 4082 37884 4088
rect 37936 4078 37964 6054
rect 39764 5024 39816 5030
rect 39764 4966 39816 4972
rect 39028 4480 39080 4486
rect 39028 4422 39080 4428
rect 37924 4072 37976 4078
rect 37924 4014 37976 4020
rect 37740 4004 37792 4010
rect 37740 3946 37792 3952
rect 38292 3936 38344 3942
rect 38292 3878 38344 3884
rect 37464 3528 37516 3534
rect 37464 3470 37516 3476
rect 37556 3392 37608 3398
rect 37556 3334 37608 3340
rect 37372 3052 37424 3058
rect 37372 2994 37424 3000
rect 37280 2440 37332 2446
rect 37280 2382 37332 2388
rect 37568 800 37596 3334
rect 38304 800 38332 3878
rect 39040 800 39068 4422
rect 39776 800 39804 4966
rect 26804 734 27016 762
rect 27066 0 27122 800
rect 27434 0 27490 800
rect 27802 0 27858 800
rect 28170 0 28226 800
rect 28538 0 28594 800
rect 28998 0 29054 800
rect 29366 0 29422 800
rect 29734 0 29790 800
rect 30102 0 30158 800
rect 30470 0 30526 800
rect 30838 0 30894 800
rect 31206 0 31262 800
rect 31574 0 31630 800
rect 31942 0 31998 800
rect 32310 0 32366 800
rect 32678 0 32734 800
rect 33046 0 33102 800
rect 33414 0 33470 800
rect 33782 0 33838 800
rect 34150 0 34206 800
rect 34610 0 34666 800
rect 34978 0 35034 800
rect 35346 0 35402 800
rect 35714 0 35770 800
rect 36082 0 36138 800
rect 36450 0 36506 800
rect 36818 0 36874 800
rect 37186 0 37242 800
rect 37554 0 37610 800
rect 37922 0 37978 800
rect 38290 0 38346 800
rect 38658 0 38714 800
rect 39026 0 39082 800
rect 39394 0 39450 800
rect 39762 0 39818 800
<< via2 >>
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 2962 6840 3018 6896
rect 2410 5344 2466 5400
rect 2686 5616 2742 5672
rect 3054 6704 3110 6760
rect 3054 6160 3110 6216
rect 2962 5752 3018 5808
rect 2870 5616 2926 5672
rect 2778 5480 2834 5536
rect 2870 5244 2872 5264
rect 2872 5244 2924 5264
rect 2924 5244 2926 5264
rect 2870 5208 2926 5244
rect 2594 4392 2650 4448
rect 2962 3304 3018 3360
rect 2870 3168 2926 3224
rect 3054 2488 3110 2544
rect 3238 7792 3294 7848
rect 3238 3440 3294 3496
rect 3422 2896 3478 2952
rect 3606 5616 3662 5672
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4618 8064 4674 8120
rect 4894 7384 4950 7440
rect 4710 7248 4766 7304
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4618 5364 4674 5400
rect 4618 5344 4620 5364
rect 4620 5344 4672 5364
rect 4672 5344 4674 5364
rect 3606 4256 3662 4312
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4158 4700 4160 4720
rect 4160 4700 4212 4720
rect 4212 4700 4214 4720
rect 4158 4664 4214 4700
rect 3882 4564 3884 4584
rect 3884 4564 3936 4584
rect 3936 4564 3938 4584
rect 3882 4528 3938 4564
rect 3698 4156 3700 4176
rect 3700 4156 3752 4176
rect 3752 4156 3754 4176
rect 3698 4120 3754 4156
rect 3790 4020 3792 4040
rect 3792 4020 3844 4040
rect 3844 4020 3846 4040
rect 3790 3984 3846 4020
rect 3698 3576 3754 3632
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4250 3032 4306 3088
rect 4618 2760 4674 2816
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 5078 8372 5080 8392
rect 5080 8372 5132 8392
rect 5132 8372 5134 8392
rect 5078 8336 5134 8372
rect 5078 6296 5134 6352
rect 4894 4256 4950 4312
rect 5262 5752 5318 5808
rect 5630 8492 5686 8528
rect 5630 8472 5632 8492
rect 5632 8472 5684 8492
rect 5684 8472 5686 8492
rect 5446 7656 5502 7712
rect 5262 3612 5264 3632
rect 5264 3612 5316 3632
rect 5316 3612 5318 3632
rect 5262 3576 5318 3612
rect 5538 6432 5594 6488
rect 5998 6704 6054 6760
rect 6458 8236 6460 8256
rect 6460 8236 6512 8256
rect 6512 8236 6514 8256
rect 6458 8200 6514 8236
rect 8850 11872 8906 11928
rect 6550 6704 6606 6760
rect 6458 6432 6514 6488
rect 5814 5208 5870 5264
rect 7378 6332 7380 6352
rect 7380 6332 7432 6352
rect 7432 6332 7434 6352
rect 6550 5208 6606 5264
rect 7378 6296 7434 6332
rect 7562 6704 7618 6760
rect 6918 2624 6974 2680
rect 8390 8200 8446 8256
rect 8022 5888 8078 5944
rect 8022 5364 8078 5400
rect 8022 5344 8024 5364
rect 8024 5344 8076 5364
rect 8076 5344 8078 5364
rect 8482 6432 8538 6488
rect 8206 6024 8262 6080
rect 8206 5616 8262 5672
rect 8298 3576 8354 3632
rect 8206 2896 8262 2952
rect 8666 6316 8722 6352
rect 8666 6296 8668 6316
rect 8668 6296 8720 6316
rect 8720 6296 8722 6316
rect 9034 6976 9090 7032
rect 8942 5752 8998 5808
rect 12346 26188 12348 26208
rect 12348 26188 12400 26208
rect 12400 26188 12402 26208
rect 12346 26152 12402 26188
rect 11978 23568 12034 23624
rect 12990 23568 13046 23624
rect 12806 23024 12862 23080
rect 12714 22480 12770 22536
rect 11794 15816 11850 15872
rect 9494 8608 9550 8664
rect 9402 7828 9404 7848
rect 9404 7828 9456 7848
rect 9456 7828 9458 7848
rect 9402 7792 9458 7828
rect 9586 7692 9588 7712
rect 9588 7692 9640 7712
rect 9640 7692 9642 7712
rect 9586 7656 9642 7692
rect 9402 7268 9458 7304
rect 9402 7248 9404 7268
rect 9404 7248 9456 7268
rect 9456 7248 9458 7268
rect 9402 6996 9458 7032
rect 9402 6976 9404 6996
rect 9404 6976 9456 6996
rect 9456 6976 9458 6996
rect 9402 6840 9458 6896
rect 9494 6568 9550 6624
rect 10046 9424 10102 9480
rect 10138 8608 10194 8664
rect 12438 15428 12494 15464
rect 12438 15408 12440 15428
rect 12440 15408 12492 15428
rect 12492 15408 12494 15428
rect 12254 13096 12310 13152
rect 12346 11872 12402 11928
rect 12254 11192 12310 11248
rect 12530 11212 12586 11248
rect 12530 11192 12532 11212
rect 12532 11192 12584 11212
rect 12584 11192 12586 11212
rect 11794 9596 11796 9616
rect 11796 9596 11848 9616
rect 11848 9596 11850 9616
rect 11794 9560 11850 9596
rect 10782 8608 10838 8664
rect 10046 7692 10048 7712
rect 10048 7692 10100 7712
rect 10100 7692 10102 7712
rect 10046 7656 10102 7692
rect 9770 5752 9826 5808
rect 10506 7828 10508 7848
rect 10508 7828 10560 7848
rect 10560 7828 10562 7848
rect 10506 7792 10562 7828
rect 9862 5616 9918 5672
rect 9770 5364 9826 5400
rect 9770 5344 9772 5364
rect 9772 5344 9824 5364
rect 9824 5344 9826 5364
rect 8758 2488 8814 2544
rect 8206 2388 8208 2408
rect 8208 2388 8260 2408
rect 8260 2388 8262 2408
rect 8206 2352 8262 2388
rect 9678 4936 9734 4992
rect 10322 5752 10378 5808
rect 10414 5480 10470 5536
rect 10322 4936 10378 4992
rect 9494 4800 9550 4856
rect 9954 4800 10010 4856
rect 10230 4800 10286 4856
rect 9310 4256 9366 4312
rect 9310 3984 9366 4040
rect 10874 6160 10930 6216
rect 10506 5344 10562 5400
rect 10690 5344 10746 5400
rect 10966 5364 11022 5400
rect 10966 5344 10968 5364
rect 10968 5344 11020 5364
rect 11020 5344 11022 5364
rect 9402 3576 9458 3632
rect 10414 3440 10470 3496
rect 9586 3032 9642 3088
rect 9310 2352 9366 2408
rect 10046 3052 10102 3088
rect 10046 3032 10048 3052
rect 10048 3032 10100 3052
rect 10100 3032 10102 3052
rect 10230 2760 10286 2816
rect 10874 4528 10930 4584
rect 10782 4392 10838 4448
rect 10966 3304 11022 3360
rect 10782 2624 10838 2680
rect 13542 22092 13598 22128
rect 13542 22072 13544 22092
rect 13544 22072 13596 22092
rect 13596 22072 13598 22092
rect 13174 17720 13230 17776
rect 13358 15272 13414 15328
rect 12714 9424 12770 9480
rect 11702 8608 11758 8664
rect 12254 8064 12310 8120
rect 11242 5752 11298 5808
rect 12346 7420 12348 7440
rect 12348 7420 12400 7440
rect 12400 7420 12402 7440
rect 12346 7384 12402 7420
rect 11426 5344 11482 5400
rect 11334 5208 11390 5264
rect 11518 4120 11574 4176
rect 12346 6876 12348 6896
rect 12348 6876 12400 6896
rect 12400 6876 12402 6896
rect 12346 6840 12402 6876
rect 12346 6316 12402 6352
rect 12346 6296 12348 6316
rect 12348 6296 12400 6316
rect 12400 6296 12402 6316
rect 12438 6160 12494 6216
rect 12346 6024 12402 6080
rect 14370 26152 14426 26208
rect 14554 22072 14610 22128
rect 14186 18128 14242 18184
rect 14922 19388 14924 19408
rect 14924 19388 14976 19408
rect 14976 19388 14978 19408
rect 14922 19352 14978 19388
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 15842 26424 15898 26480
rect 15566 26288 15622 26344
rect 15934 26288 15990 26344
rect 14922 18708 14924 18728
rect 14924 18708 14976 18728
rect 14976 18708 14978 18728
rect 14922 18672 14978 18708
rect 14462 15544 14518 15600
rect 13542 9560 13598 9616
rect 13634 8472 13690 8528
rect 13082 7656 13138 7712
rect 13450 6840 13506 6896
rect 12530 5616 12586 5672
rect 11886 5480 11942 5536
rect 12714 5480 12770 5536
rect 11978 5072 12034 5128
rect 11702 4664 11758 4720
rect 12254 4800 12310 4856
rect 12530 4800 12586 4856
rect 12162 3340 12164 3360
rect 12164 3340 12216 3360
rect 12216 3340 12218 3360
rect 12162 3304 12218 3340
rect 12162 3168 12218 3224
rect 13358 5344 13414 5400
rect 13082 3576 13138 3632
rect 14186 6296 14242 6352
rect 14002 5636 14058 5672
rect 14002 5616 14004 5636
rect 14004 5616 14056 5636
rect 14056 5616 14058 5636
rect 13910 4256 13966 4312
rect 13910 3032 13966 3088
rect 16302 26424 16358 26480
rect 15658 17448 15714 17504
rect 16118 17448 16174 17504
rect 17038 26308 17094 26344
rect 17038 26288 17040 26308
rect 17040 26288 17092 26308
rect 17092 26288 17094 26308
rect 16670 26152 16726 26208
rect 16578 18944 16634 19000
rect 16578 14068 16634 14104
rect 16578 14048 16580 14068
rect 16580 14048 16632 14068
rect 16632 14048 16634 14068
rect 16854 15816 16910 15872
rect 16946 15408 17002 15464
rect 17406 18944 17462 19000
rect 17498 18808 17554 18864
rect 17130 18128 17186 18184
rect 17866 19372 17922 19408
rect 17866 19352 17868 19372
rect 17868 19352 17920 19372
rect 17920 19352 17922 19372
rect 17866 18964 17922 19000
rect 17866 18944 17868 18964
rect 17868 18944 17920 18964
rect 17920 18944 17922 18964
rect 17958 17876 18014 17912
rect 17958 17856 17960 17876
rect 17960 17856 18012 17876
rect 18012 17856 18014 17876
rect 18326 18708 18328 18728
rect 18328 18708 18380 18728
rect 18380 18708 18382 18728
rect 18326 18672 18382 18708
rect 17958 17620 17960 17640
rect 17960 17620 18012 17640
rect 18012 17620 18014 17640
rect 17958 17584 18014 17620
rect 18234 17720 18290 17776
rect 17498 15952 17554 16008
rect 17222 14884 17278 14920
rect 17222 14864 17224 14884
rect 17224 14864 17276 14884
rect 17276 14864 17278 14884
rect 17314 14612 17370 14648
rect 17314 14592 17316 14612
rect 17316 14592 17368 14612
rect 17368 14592 17370 14612
rect 18510 18828 18566 18864
rect 18510 18808 18512 18828
rect 18512 18808 18564 18828
rect 18564 18808 18566 18828
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 20074 27820 20076 27840
rect 20076 27820 20128 27840
rect 20128 27820 20130 27840
rect 20074 27784 20130 27820
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 18602 14864 18658 14920
rect 14370 4664 14426 4720
rect 15014 6160 15070 6216
rect 15934 5616 15990 5672
rect 15382 3304 15438 3360
rect 17498 9424 17554 9480
rect 18694 9696 18750 9752
rect 17222 6432 17278 6488
rect 17130 5888 17186 5944
rect 19706 19760 19762 19816
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19430 19352 19486 19408
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19154 17720 19210 17776
rect 17774 5888 17830 5944
rect 17774 5208 17830 5264
rect 18510 4800 18566 4856
rect 17958 3052 18014 3088
rect 17958 3032 17960 3052
rect 17960 3032 18012 3052
rect 18012 3032 18014 3052
rect 18234 3068 18236 3088
rect 18236 3068 18288 3088
rect 18288 3068 18290 3088
rect 18234 3032 18290 3068
rect 19246 17620 19248 17640
rect 19248 17620 19300 17640
rect 19300 17620 19302 17640
rect 19246 17584 19302 17620
rect 19706 17620 19708 17640
rect 19708 17620 19760 17640
rect 19760 17620 19762 17640
rect 19706 17584 19762 17620
rect 19246 14900 19248 14920
rect 19248 14900 19300 14920
rect 19300 14900 19302 14920
rect 19246 14864 19302 14900
rect 19338 14048 19394 14104
rect 19246 13096 19302 13152
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19798 17176 19854 17232
rect 19614 17040 19670 17096
rect 19706 16904 19762 16960
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 20810 29008 20866 29064
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 20074 17584 20130 17640
rect 20442 16904 20498 16960
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19522 15680 19578 15736
rect 19522 15428 19578 15464
rect 19522 15408 19524 15428
rect 19524 15408 19576 15428
rect 19576 15408 19578 15428
rect 19982 15408 20038 15464
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19614 10648 19670 10704
rect 19890 10512 19946 10568
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19430 9696 19486 9752
rect 19798 9580 19854 9616
rect 19798 9560 19800 9580
rect 19800 9560 19852 9580
rect 19852 9560 19854 9580
rect 20350 14592 20406 14648
rect 22190 29008 22246 29064
rect 20258 11872 20314 11928
rect 20166 10376 20222 10432
rect 20074 9424 20130 9480
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 20350 9580 20406 9616
rect 20350 9560 20352 9580
rect 20352 9560 20404 9580
rect 20404 9560 20406 9580
rect 20258 8508 20260 8528
rect 20260 8508 20312 8528
rect 20312 8508 20314 8528
rect 20258 8472 20314 8508
rect 19246 6196 19248 6216
rect 19248 6196 19300 6216
rect 19300 6196 19302 6216
rect 19246 6160 19302 6196
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19982 6024 20038 6080
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19246 4936 19302 4992
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19430 3984 19486 4040
rect 19522 3848 19578 3904
rect 19982 3984 20038 4040
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20718 17584 20774 17640
rect 20902 17856 20958 17912
rect 20442 6160 20498 6216
rect 20350 5072 20406 5128
rect 20442 3848 20498 3904
rect 21178 11736 21234 11792
rect 22098 21972 22100 21992
rect 22100 21972 22152 21992
rect 22152 21972 22154 21992
rect 22098 21936 22154 21972
rect 22006 21800 22062 21856
rect 22098 21664 22154 21720
rect 22742 27784 22798 27840
rect 22466 24812 22522 24848
rect 22466 24792 22468 24812
rect 22468 24792 22520 24812
rect 22520 24792 22522 24812
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 22742 21936 22798 21992
rect 22834 21800 22890 21856
rect 21730 17312 21786 17368
rect 22190 17212 22192 17232
rect 22192 17212 22244 17232
rect 22244 17212 22246 17232
rect 22190 17176 22246 17212
rect 21822 17076 21824 17096
rect 21824 17076 21876 17096
rect 21876 17076 21878 17096
rect 21822 17040 21878 17076
rect 21454 4256 21510 4312
rect 21914 9424 21970 9480
rect 21822 9152 21878 9208
rect 21914 5752 21970 5808
rect 21914 3848 21970 3904
rect 22190 11500 22192 11520
rect 22192 11500 22244 11520
rect 22244 11500 22246 11520
rect 22190 11464 22246 11500
rect 22098 9460 22100 9480
rect 22100 9460 22152 9480
rect 22152 9460 22154 9480
rect 22098 9424 22154 9460
rect 22374 5888 22430 5944
rect 22098 3884 22100 3904
rect 22100 3884 22152 3904
rect 22152 3884 22154 3904
rect 22098 3848 22154 3884
rect 23662 18128 23718 18184
rect 23478 17176 23534 17232
rect 23478 15680 23534 15736
rect 22650 6296 22706 6352
rect 23386 6024 23442 6080
rect 24030 15544 24086 15600
rect 23754 11464 23810 11520
rect 24858 17040 24914 17096
rect 24674 15544 24730 15600
rect 24490 10240 24546 10296
rect 26146 24792 26202 24848
rect 25318 10240 25374 10296
rect 24766 9580 24822 9616
rect 24766 9560 24768 9580
rect 24768 9560 24820 9580
rect 24820 9560 24822 9580
rect 24674 9460 24676 9480
rect 24676 9460 24728 9480
rect 24728 9460 24730 9480
rect 24674 9424 24730 9460
rect 24766 9016 24822 9072
rect 26238 21664 26294 21720
rect 25962 19352 26018 19408
rect 26238 19372 26294 19408
rect 26238 19352 26240 19372
rect 26240 19352 26292 19372
rect 26292 19352 26294 19372
rect 25962 17312 26018 17368
rect 26146 18164 26148 18184
rect 26148 18164 26200 18184
rect 26200 18164 26202 18184
rect 26146 18128 26202 18164
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 24766 6740 24768 6760
rect 24768 6740 24820 6760
rect 24820 6740 24822 6760
rect 24766 6704 24822 6740
rect 24766 5888 24822 5944
rect 24766 5480 24822 5536
rect 24490 3032 24546 3088
rect 25502 6160 25558 6216
rect 25410 5480 25466 5536
rect 25318 3984 25374 4040
rect 26054 9424 26110 9480
rect 26238 10412 26240 10432
rect 26240 10412 26292 10432
rect 26292 10412 26294 10432
rect 26238 10376 26294 10412
rect 26238 9052 26240 9072
rect 26240 9052 26292 9072
rect 26292 9052 26294 9072
rect 26238 9016 26294 9052
rect 27434 19352 27490 19408
rect 25870 6160 25926 6216
rect 27342 17076 27344 17096
rect 27344 17076 27396 17096
rect 27396 17076 27398 17096
rect 27342 17040 27398 17076
rect 26974 8200 27030 8256
rect 26882 6976 26938 7032
rect 26882 5908 26938 5944
rect 26882 5888 26884 5908
rect 26884 5888 26936 5908
rect 26936 5888 26938 5908
rect 27158 10240 27214 10296
rect 27250 9560 27306 9616
rect 27434 10668 27490 10704
rect 27434 10648 27436 10668
rect 27436 10648 27488 10668
rect 27488 10648 27490 10668
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 27618 9152 27674 9208
rect 27158 8336 27214 8392
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 27710 8472 27766 8528
rect 27250 6704 27306 6760
rect 28998 11756 29054 11792
rect 28998 11736 29000 11756
rect 29000 11736 29052 11756
rect 29052 11736 29054 11756
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 28446 10376 28502 10432
rect 28262 8236 28264 8256
rect 28264 8236 28316 8256
rect 28316 8236 28318 8256
rect 28262 8200 28318 8236
rect 28722 10532 28778 10568
rect 28722 10512 28724 10532
rect 28724 10512 28776 10532
rect 28776 10512 28778 10532
rect 28354 5772 28410 5808
rect 28354 5752 28356 5772
rect 28356 5752 28408 5772
rect 28408 5752 28410 5772
rect 29182 10140 29184 10160
rect 29184 10140 29236 10160
rect 29236 10140 29238 10160
rect 29182 10104 29238 10140
rect 29182 7792 29238 7848
rect 28814 5072 28870 5128
rect 29734 11092 29736 11112
rect 29736 11092 29788 11112
rect 29788 11092 29790 11112
rect 29734 11056 29790 11092
rect 30194 9968 30250 10024
rect 29734 9696 29790 9752
rect 29734 5752 29790 5808
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 31022 9868 31024 9888
rect 31024 9868 31076 9888
rect 31076 9868 31078 9888
rect 31022 9832 31078 9868
rect 30654 9696 30710 9752
rect 31206 9016 31262 9072
rect 31206 8336 31262 8392
rect 30930 5616 30986 5672
rect 31666 6024 31722 6080
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 32770 5752 32826 5808
rect 32770 4528 32826 4584
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34610 4800 34666 4856
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34886 4664 34942 4720
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35714 4564 35716 4584
rect 35716 4564 35768 4584
rect 35768 4564 35770 4584
rect 35714 4528 35770 4564
<< metal3 >>
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 20805 29066 20871 29069
rect 22185 29066 22251 29069
rect 20805 29064 22251 29066
rect 20805 29008 20810 29064
rect 20866 29008 22190 29064
rect 22246 29008 22251 29064
rect 20805 29006 22251 29008
rect 20805 29003 20871 29006
rect 22185 29003 22251 29006
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 20069 27842 20135 27845
rect 22737 27842 22803 27845
rect 20069 27840 22803 27842
rect 20069 27784 20074 27840
rect 20130 27784 22742 27840
rect 22798 27784 22803 27840
rect 20069 27782 22803 27784
rect 20069 27779 20135 27782
rect 22737 27779 22803 27782
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 15837 26482 15903 26485
rect 16297 26482 16363 26485
rect 15837 26480 16363 26482
rect 15837 26424 15842 26480
rect 15898 26424 16302 26480
rect 16358 26424 16363 26480
rect 15837 26422 16363 26424
rect 15837 26419 15903 26422
rect 16297 26419 16363 26422
rect 15561 26346 15627 26349
rect 15929 26346 15995 26349
rect 17033 26346 17099 26349
rect 15561 26344 17099 26346
rect 15561 26288 15566 26344
rect 15622 26288 15934 26344
rect 15990 26288 17038 26344
rect 17094 26288 17099 26344
rect 15561 26286 17099 26288
rect 15561 26283 15627 26286
rect 15929 26283 15995 26286
rect 17033 26283 17099 26286
rect 12341 26210 12407 26213
rect 14365 26210 14431 26213
rect 16665 26210 16731 26213
rect 12341 26208 16731 26210
rect 12341 26152 12346 26208
rect 12402 26152 14370 26208
rect 14426 26152 16670 26208
rect 16726 26152 16731 26208
rect 12341 26150 16731 26152
rect 12341 26147 12407 26150
rect 14365 26147 14431 26150
rect 16665 26147 16731 26150
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 22461 24850 22527 24853
rect 26141 24850 26207 24853
rect 22461 24848 26207 24850
rect 22461 24792 22466 24848
rect 22522 24792 26146 24848
rect 26202 24792 26207 24848
rect 22461 24790 26207 24792
rect 22461 24787 22527 24790
rect 26141 24787 26207 24790
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 11973 23626 12039 23629
rect 12985 23626 13051 23629
rect 11973 23624 13051 23626
rect 11973 23568 11978 23624
rect 12034 23568 12990 23624
rect 13046 23568 13051 23624
rect 11973 23566 13051 23568
rect 11973 23563 12039 23566
rect 12985 23563 13051 23566
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 12801 23082 12867 23085
rect 12758 23080 12867 23082
rect 12758 23024 12806 23080
rect 12862 23024 12867 23080
rect 12758 23019 12867 23024
rect 12758 22541 12818 23019
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 12709 22536 12818 22541
rect 12709 22480 12714 22536
rect 12770 22480 12818 22536
rect 12709 22478 12818 22480
rect 12709 22475 12775 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 13537 22130 13603 22133
rect 14549 22130 14615 22133
rect 13537 22128 14615 22130
rect 13537 22072 13542 22128
rect 13598 22072 14554 22128
rect 14610 22072 14615 22128
rect 13537 22070 14615 22072
rect 13537 22067 13603 22070
rect 14549 22067 14615 22070
rect 22093 21994 22159 21997
rect 22737 21994 22803 21997
rect 22093 21992 22803 21994
rect 22093 21936 22098 21992
rect 22154 21936 22742 21992
rect 22798 21936 22803 21992
rect 22093 21934 22803 21936
rect 22093 21931 22159 21934
rect 22737 21931 22803 21934
rect 22001 21858 22067 21861
rect 22829 21858 22895 21861
rect 22001 21856 22895 21858
rect 22001 21800 22006 21856
rect 22062 21800 22834 21856
rect 22890 21800 22895 21856
rect 22001 21798 22895 21800
rect 22001 21795 22067 21798
rect 22829 21795 22895 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 22093 21722 22159 21725
rect 26233 21722 26299 21725
rect 22093 21720 26299 21722
rect 22093 21664 22098 21720
rect 22154 21664 26238 21720
rect 26294 21664 26299 21720
rect 22093 21662 26299 21664
rect 22093 21659 22159 21662
rect 26233 21659 26299 21662
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 19374 19756 19380 19820
rect 19444 19818 19450 19820
rect 19701 19818 19767 19821
rect 19444 19816 19767 19818
rect 19444 19760 19706 19816
rect 19762 19760 19767 19816
rect 19444 19758 19767 19760
rect 19444 19756 19450 19758
rect 19701 19755 19767 19758
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 14917 19410 14983 19413
rect 17861 19410 17927 19413
rect 14917 19408 17927 19410
rect 14917 19352 14922 19408
rect 14978 19352 17866 19408
rect 17922 19352 17927 19408
rect 14917 19350 17927 19352
rect 14917 19347 14983 19350
rect 17861 19347 17927 19350
rect 19425 19410 19491 19413
rect 25957 19410 26023 19413
rect 26233 19410 26299 19413
rect 27429 19410 27495 19413
rect 19425 19408 27495 19410
rect 19425 19352 19430 19408
rect 19486 19352 25962 19408
rect 26018 19352 26238 19408
rect 26294 19352 27434 19408
rect 27490 19352 27495 19408
rect 19425 19350 27495 19352
rect 19425 19347 19491 19350
rect 25957 19347 26023 19350
rect 26233 19347 26299 19350
rect 27429 19347 27495 19350
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 16573 19002 16639 19005
rect 17401 19002 17467 19005
rect 17861 19002 17927 19005
rect 16573 19000 17927 19002
rect 16573 18944 16578 19000
rect 16634 18944 17406 19000
rect 17462 18944 17866 19000
rect 17922 18944 17927 19000
rect 16573 18942 17927 18944
rect 16573 18939 16639 18942
rect 17401 18939 17467 18942
rect 17861 18939 17927 18942
rect 17493 18866 17559 18869
rect 18505 18866 18571 18869
rect 17493 18864 18571 18866
rect 17493 18808 17498 18864
rect 17554 18808 18510 18864
rect 18566 18808 18571 18864
rect 17493 18806 18571 18808
rect 17493 18803 17559 18806
rect 18505 18803 18571 18806
rect 14917 18730 14983 18733
rect 18321 18730 18387 18733
rect 14917 18728 18387 18730
rect 14917 18672 14922 18728
rect 14978 18672 18326 18728
rect 18382 18672 18387 18728
rect 14917 18670 18387 18672
rect 14917 18667 14983 18670
rect 18321 18667 18387 18670
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 14181 18186 14247 18189
rect 17125 18186 17191 18189
rect 14181 18184 17191 18186
rect 14181 18128 14186 18184
rect 14242 18128 17130 18184
rect 17186 18128 17191 18184
rect 14181 18126 17191 18128
rect 14181 18123 14247 18126
rect 17125 18123 17191 18126
rect 23657 18186 23723 18189
rect 26141 18186 26207 18189
rect 23657 18184 26207 18186
rect 23657 18128 23662 18184
rect 23718 18128 26146 18184
rect 26202 18128 26207 18184
rect 23657 18126 26207 18128
rect 23657 18123 23723 18126
rect 26141 18123 26207 18126
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 17953 17914 18019 17917
rect 20897 17914 20963 17917
rect 17953 17912 20963 17914
rect 17953 17856 17958 17912
rect 18014 17856 20902 17912
rect 20958 17856 20963 17912
rect 17953 17854 20963 17856
rect 17953 17851 18019 17854
rect 20897 17851 20963 17854
rect 13169 17778 13235 17781
rect 18229 17778 18295 17781
rect 19149 17778 19215 17781
rect 13169 17776 19215 17778
rect 13169 17720 13174 17776
rect 13230 17720 18234 17776
rect 18290 17720 19154 17776
rect 19210 17720 19215 17776
rect 13169 17718 19215 17720
rect 13169 17715 13235 17718
rect 18229 17715 18295 17718
rect 19149 17715 19215 17718
rect 17953 17642 18019 17645
rect 19241 17642 19307 17645
rect 19701 17642 19767 17645
rect 17953 17640 19307 17642
rect 17953 17584 17958 17640
rect 18014 17584 19246 17640
rect 19302 17584 19307 17640
rect 17953 17582 19307 17584
rect 17953 17579 18019 17582
rect 19241 17579 19307 17582
rect 19428 17640 19767 17642
rect 19428 17584 19706 17640
rect 19762 17584 19767 17640
rect 19428 17582 19767 17584
rect 15653 17506 15719 17509
rect 16113 17506 16179 17509
rect 15653 17504 16179 17506
rect 15653 17448 15658 17504
rect 15714 17448 16118 17504
rect 16174 17448 16179 17504
rect 15653 17446 16179 17448
rect 15653 17443 15719 17446
rect 16113 17443 16179 17446
rect 19428 17234 19488 17582
rect 19701 17579 19767 17582
rect 20069 17642 20135 17645
rect 20713 17642 20779 17645
rect 20069 17640 20779 17642
rect 20069 17584 20074 17640
rect 20130 17584 20718 17640
rect 20774 17584 20779 17640
rect 20069 17582 20779 17584
rect 20069 17579 20135 17582
rect 20713 17579 20779 17582
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 21725 17370 21791 17373
rect 25957 17370 26023 17373
rect 21725 17368 26023 17370
rect 21725 17312 21730 17368
rect 21786 17312 25962 17368
rect 26018 17312 26023 17368
rect 21725 17310 26023 17312
rect 21725 17307 21791 17310
rect 25957 17307 26023 17310
rect 19793 17234 19859 17237
rect 19428 17232 19859 17234
rect 19428 17176 19798 17232
rect 19854 17176 19859 17232
rect 19428 17174 19859 17176
rect 19793 17171 19859 17174
rect 22185 17234 22251 17237
rect 23473 17234 23539 17237
rect 22185 17232 23539 17234
rect 22185 17176 22190 17232
rect 22246 17176 23478 17232
rect 23534 17176 23539 17232
rect 22185 17174 23539 17176
rect 22185 17171 22251 17174
rect 23473 17171 23539 17174
rect 19609 17098 19675 17101
rect 21817 17098 21883 17101
rect 24853 17098 24919 17101
rect 27337 17098 27403 17101
rect 19609 17096 27403 17098
rect 19609 17040 19614 17096
rect 19670 17040 21822 17096
rect 21878 17040 24858 17096
rect 24914 17040 27342 17096
rect 27398 17040 27403 17096
rect 19609 17038 27403 17040
rect 19609 17035 19675 17038
rect 21817 17035 21883 17038
rect 24853 17035 24919 17038
rect 27337 17035 27403 17038
rect 19701 16962 19767 16965
rect 20294 16962 20300 16964
rect 19701 16960 20300 16962
rect 19701 16904 19706 16960
rect 19762 16904 20300 16960
rect 19701 16902 20300 16904
rect 19701 16899 19767 16902
rect 20294 16900 20300 16902
rect 20364 16962 20370 16964
rect 20437 16962 20503 16965
rect 20364 16960 20503 16962
rect 20364 16904 20442 16960
rect 20498 16904 20503 16960
rect 20364 16902 20503 16904
rect 20364 16900 20370 16902
rect 20437 16899 20503 16902
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 17493 16012 17559 16013
rect 17493 16010 17540 16012
rect 17448 16008 17540 16010
rect 17448 15952 17498 16008
rect 17448 15950 17540 15952
rect 17493 15948 17540 15950
rect 17604 15948 17610 16012
rect 17493 15947 17559 15948
rect 11789 15874 11855 15877
rect 16849 15874 16915 15877
rect 11789 15872 16915 15874
rect 11789 15816 11794 15872
rect 11850 15816 16854 15872
rect 16910 15816 16915 15872
rect 11789 15814 16915 15816
rect 11789 15811 11855 15814
rect 16849 15811 16915 15814
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 19517 15738 19583 15741
rect 23473 15738 23539 15741
rect 19517 15736 23539 15738
rect 19517 15680 19522 15736
rect 19578 15680 23478 15736
rect 23534 15680 23539 15736
rect 19517 15678 23539 15680
rect 19517 15675 19583 15678
rect 23473 15675 23539 15678
rect 14457 15602 14523 15605
rect 24025 15602 24091 15605
rect 24669 15602 24735 15605
rect 14457 15600 24735 15602
rect 14457 15544 14462 15600
rect 14518 15544 24030 15600
rect 24086 15544 24674 15600
rect 24730 15544 24735 15600
rect 14457 15542 24735 15544
rect 14457 15539 14523 15542
rect 24025 15539 24091 15542
rect 24669 15539 24735 15542
rect 12433 15466 12499 15469
rect 16941 15466 17007 15469
rect 12433 15464 17007 15466
rect 12433 15408 12438 15464
rect 12494 15408 16946 15464
rect 17002 15408 17007 15464
rect 12433 15406 17007 15408
rect 12433 15403 12499 15406
rect 16941 15403 17007 15406
rect 19517 15466 19583 15469
rect 19977 15466 20043 15469
rect 19517 15464 20043 15466
rect 19517 15408 19522 15464
rect 19578 15408 19982 15464
rect 20038 15408 20043 15464
rect 19517 15406 20043 15408
rect 19517 15403 19583 15406
rect 19977 15403 20043 15406
rect 13353 15330 13419 15333
rect 19374 15330 19380 15332
rect 13353 15328 19380 15330
rect 13353 15272 13358 15328
rect 13414 15272 19380 15328
rect 13353 15270 19380 15272
rect 13353 15267 13419 15270
rect 19374 15268 19380 15270
rect 19444 15268 19450 15332
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 17217 14922 17283 14925
rect 18597 14922 18663 14925
rect 19241 14922 19307 14925
rect 17217 14920 19307 14922
rect 17217 14864 17222 14920
rect 17278 14864 18602 14920
rect 18658 14864 19246 14920
rect 19302 14864 19307 14920
rect 17217 14862 19307 14864
rect 17217 14859 17283 14862
rect 18597 14859 18663 14862
rect 19241 14859 19307 14862
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 17309 14650 17375 14653
rect 20345 14650 20411 14653
rect 17309 14648 20411 14650
rect 17309 14592 17314 14648
rect 17370 14592 20350 14648
rect 20406 14592 20411 14648
rect 17309 14590 20411 14592
rect 17309 14587 17375 14590
rect 20345 14587 20411 14590
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 16573 14106 16639 14109
rect 19333 14106 19399 14109
rect 16573 14104 19399 14106
rect 16573 14048 16578 14104
rect 16634 14048 19338 14104
rect 19394 14048 19399 14104
rect 16573 14046 19399 14048
rect 16573 14043 16639 14046
rect 19333 14043 19399 14046
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 12249 13154 12315 13157
rect 19241 13154 19307 13157
rect 12249 13152 19307 13154
rect 12249 13096 12254 13152
rect 12310 13096 19246 13152
rect 19302 13096 19307 13152
rect 12249 13094 19307 13096
rect 12249 13091 12315 13094
rect 19241 13091 19307 13094
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 8845 11930 8911 11933
rect 12341 11930 12407 11933
rect 8845 11928 12407 11930
rect 8845 11872 8850 11928
rect 8906 11872 12346 11928
rect 12402 11872 12407 11928
rect 8845 11870 12407 11872
rect 8845 11867 8911 11870
rect 12341 11867 12407 11870
rect 20253 11932 20319 11933
rect 20253 11928 20300 11932
rect 20364 11930 20370 11932
rect 20253 11872 20258 11928
rect 20253 11868 20300 11872
rect 20364 11870 20410 11930
rect 20364 11868 20370 11870
rect 20253 11867 20319 11868
rect 21173 11794 21239 11797
rect 28993 11794 29059 11797
rect 21173 11792 29059 11794
rect 21173 11736 21178 11792
rect 21234 11736 28998 11792
rect 29054 11736 29059 11792
rect 21173 11734 29059 11736
rect 21173 11731 21239 11734
rect 28993 11731 29059 11734
rect 22185 11522 22251 11525
rect 23749 11522 23815 11525
rect 22185 11520 23815 11522
rect 22185 11464 22190 11520
rect 22246 11464 23754 11520
rect 23810 11464 23815 11520
rect 22185 11462 23815 11464
rect 22185 11459 22251 11462
rect 23749 11459 23815 11462
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 12249 11250 12315 11253
rect 12525 11250 12591 11253
rect 12249 11248 12591 11250
rect 12249 11192 12254 11248
rect 12310 11192 12530 11248
rect 12586 11192 12591 11248
rect 12249 11190 12591 11192
rect 12249 11187 12315 11190
rect 12525 11187 12591 11190
rect 25814 11052 25820 11116
rect 25884 11114 25890 11116
rect 29729 11114 29795 11117
rect 25884 11112 29795 11114
rect 25884 11056 29734 11112
rect 29790 11056 29795 11112
rect 25884 11054 29795 11056
rect 25884 11052 25890 11054
rect 29729 11051 29795 11054
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 19609 10706 19675 10709
rect 27429 10706 27495 10709
rect 19609 10704 27495 10706
rect 19609 10648 19614 10704
rect 19670 10648 27434 10704
rect 27490 10648 27495 10704
rect 19609 10646 27495 10648
rect 19609 10643 19675 10646
rect 27429 10643 27495 10646
rect 19885 10570 19951 10573
rect 28717 10570 28783 10573
rect 19885 10568 28783 10570
rect 19885 10512 19890 10568
rect 19946 10512 28722 10568
rect 28778 10512 28783 10568
rect 19885 10510 28783 10512
rect 19885 10507 19951 10510
rect 28717 10507 28783 10510
rect 20161 10434 20227 10437
rect 26233 10434 26299 10437
rect 28441 10434 28507 10437
rect 20161 10432 28507 10434
rect 20161 10376 20166 10432
rect 20222 10376 26238 10432
rect 26294 10376 28446 10432
rect 28502 10376 28507 10432
rect 20161 10374 28507 10376
rect 20161 10371 20227 10374
rect 26233 10371 26299 10374
rect 28441 10371 28507 10374
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 24485 10298 24551 10301
rect 25313 10298 25379 10301
rect 27153 10298 27219 10301
rect 24485 10296 27219 10298
rect 24485 10240 24490 10296
rect 24546 10240 25318 10296
rect 25374 10240 27158 10296
rect 27214 10240 27219 10296
rect 24485 10238 27219 10240
rect 24485 10235 24551 10238
rect 25313 10235 25379 10238
rect 27153 10235 27219 10238
rect 29177 10164 29243 10165
rect 29126 10162 29132 10164
rect 29086 10102 29132 10162
rect 29196 10160 29243 10164
rect 29238 10104 29243 10160
rect 29126 10100 29132 10102
rect 29196 10100 29243 10104
rect 29177 10099 29243 10100
rect 28942 9964 28948 10028
rect 29012 10026 29018 10028
rect 30189 10026 30255 10029
rect 29012 10024 30255 10026
rect 29012 9968 30194 10024
rect 30250 9968 30255 10024
rect 29012 9966 30255 9968
rect 29012 9964 29018 9966
rect 30189 9963 30255 9966
rect 24710 9828 24716 9892
rect 24780 9890 24786 9892
rect 31017 9890 31083 9893
rect 24780 9888 31083 9890
rect 24780 9832 31022 9888
rect 31078 9832 31083 9888
rect 24780 9830 31083 9832
rect 24780 9828 24786 9830
rect 31017 9827 31083 9830
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 18689 9754 18755 9757
rect 19425 9754 19491 9757
rect 18689 9752 19491 9754
rect 18689 9696 18694 9752
rect 18750 9696 19430 9752
rect 19486 9696 19491 9752
rect 18689 9694 19491 9696
rect 18689 9691 18755 9694
rect 19425 9691 19491 9694
rect 27654 9692 27660 9756
rect 27724 9754 27730 9756
rect 29729 9754 29795 9757
rect 27724 9752 29795 9754
rect 27724 9696 29734 9752
rect 29790 9696 29795 9752
rect 27724 9694 29795 9696
rect 27724 9692 27730 9694
rect 29729 9691 29795 9694
rect 30414 9692 30420 9756
rect 30484 9754 30490 9756
rect 30649 9754 30715 9757
rect 30484 9752 30715 9754
rect 30484 9696 30654 9752
rect 30710 9696 30715 9752
rect 30484 9694 30715 9696
rect 30484 9692 30490 9694
rect 30649 9691 30715 9694
rect 11789 9618 11855 9621
rect 13537 9618 13603 9621
rect 11789 9616 13603 9618
rect 11789 9560 11794 9616
rect 11850 9560 13542 9616
rect 13598 9560 13603 9616
rect 11789 9558 13603 9560
rect 11789 9555 11855 9558
rect 13537 9555 13603 9558
rect 19793 9618 19859 9621
rect 20345 9618 20411 9621
rect 19793 9616 20411 9618
rect 19793 9560 19798 9616
rect 19854 9560 20350 9616
rect 20406 9560 20411 9616
rect 19793 9558 20411 9560
rect 19793 9555 19859 9558
rect 20345 9555 20411 9558
rect 24761 9618 24827 9621
rect 27245 9618 27311 9621
rect 24761 9616 27311 9618
rect 24761 9560 24766 9616
rect 24822 9560 27250 9616
rect 27306 9560 27311 9616
rect 24761 9558 27311 9560
rect 24761 9555 24827 9558
rect 27245 9555 27311 9558
rect 10041 9482 10107 9485
rect 12709 9482 12775 9485
rect 17493 9482 17559 9485
rect 10041 9480 17559 9482
rect 10041 9424 10046 9480
rect 10102 9424 12714 9480
rect 12770 9424 17498 9480
rect 17554 9424 17559 9480
rect 10041 9422 17559 9424
rect 10041 9419 10107 9422
rect 12709 9419 12775 9422
rect 17493 9419 17559 9422
rect 19374 9420 19380 9484
rect 19444 9482 19450 9484
rect 20069 9482 20135 9485
rect 19444 9480 20135 9482
rect 19444 9424 20074 9480
rect 20130 9424 20135 9480
rect 19444 9422 20135 9424
rect 19444 9420 19450 9422
rect 20069 9419 20135 9422
rect 21909 9482 21975 9485
rect 22093 9482 22159 9485
rect 21909 9480 22159 9482
rect 21909 9424 21914 9480
rect 21970 9424 22098 9480
rect 22154 9424 22159 9480
rect 21909 9422 22159 9424
rect 21909 9419 21975 9422
rect 22093 9419 22159 9422
rect 24669 9482 24735 9485
rect 26049 9482 26115 9485
rect 24669 9480 26115 9482
rect 24669 9424 24674 9480
rect 24730 9424 26054 9480
rect 26110 9424 26115 9480
rect 24669 9422 26115 9424
rect 24669 9419 24735 9422
rect 26049 9419 26115 9422
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 21817 9210 21883 9213
rect 27613 9210 27679 9213
rect 21817 9208 27679 9210
rect 21817 9152 21822 9208
rect 21878 9152 27618 9208
rect 27674 9152 27679 9208
rect 21817 9150 27679 9152
rect 21817 9147 21883 9150
rect 27613 9147 27679 9150
rect 24761 9074 24827 9077
rect 26233 9074 26299 9077
rect 24761 9072 26299 9074
rect 24761 9016 24766 9072
rect 24822 9016 26238 9072
rect 26294 9016 26299 9072
rect 24761 9014 26299 9016
rect 24761 9011 24827 9014
rect 26233 9011 26299 9014
rect 30598 9012 30604 9076
rect 30668 9074 30674 9076
rect 31201 9074 31267 9077
rect 30668 9072 31267 9074
rect 30668 9016 31206 9072
rect 31262 9016 31267 9072
rect 30668 9014 31267 9016
rect 30668 9012 30674 9014
rect 31201 9011 31267 9014
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 9489 8668 9555 8669
rect 9438 8666 9444 8668
rect 9398 8606 9444 8666
rect 9508 8664 9555 8668
rect 9550 8608 9555 8664
rect 9438 8604 9444 8606
rect 9508 8604 9555 8608
rect 9489 8603 9555 8604
rect 10133 8666 10199 8669
rect 10777 8666 10843 8669
rect 11697 8666 11763 8669
rect 10133 8664 11763 8666
rect 10133 8608 10138 8664
rect 10194 8608 10782 8664
rect 10838 8608 11702 8664
rect 11758 8608 11763 8664
rect 10133 8606 11763 8608
rect 10133 8603 10199 8606
rect 10777 8603 10843 8606
rect 11697 8603 11763 8606
rect 5625 8530 5691 8533
rect 13629 8530 13695 8533
rect 5625 8528 13695 8530
rect 5625 8472 5630 8528
rect 5686 8472 13634 8528
rect 13690 8472 13695 8528
rect 5625 8470 13695 8472
rect 5625 8467 5691 8470
rect 13629 8467 13695 8470
rect 20253 8530 20319 8533
rect 27705 8530 27771 8533
rect 20253 8528 27771 8530
rect 20253 8472 20258 8528
rect 20314 8472 27710 8528
rect 27766 8472 27771 8528
rect 20253 8470 27771 8472
rect 20253 8467 20319 8470
rect 27705 8467 27771 8470
rect 5073 8394 5139 8397
rect 27153 8394 27219 8397
rect 31201 8394 31267 8397
rect 5073 8392 12450 8394
rect 5073 8336 5078 8392
rect 5134 8336 12450 8392
rect 5073 8334 12450 8336
rect 5073 8331 5139 8334
rect 6453 8258 6519 8261
rect 8385 8258 8451 8261
rect 6453 8256 8451 8258
rect 6453 8200 6458 8256
rect 6514 8200 8390 8256
rect 8446 8200 8451 8256
rect 6453 8198 8451 8200
rect 6453 8195 6519 8198
rect 8385 8195 8451 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 4613 8122 4679 8125
rect 12249 8122 12315 8125
rect 4613 8120 12315 8122
rect 4613 8064 4618 8120
rect 4674 8064 12254 8120
rect 12310 8064 12315 8120
rect 4613 8062 12315 8064
rect 4613 8059 4679 8062
rect 12249 8059 12315 8062
rect 3233 7850 3299 7853
rect 9397 7850 9463 7853
rect 3233 7848 9463 7850
rect 3233 7792 3238 7848
rect 3294 7792 9402 7848
rect 9458 7792 9463 7848
rect 3233 7790 9463 7792
rect 3233 7787 3299 7790
rect 9397 7787 9463 7790
rect 10358 7788 10364 7852
rect 10428 7850 10434 7852
rect 10501 7850 10567 7853
rect 10428 7848 10567 7850
rect 10428 7792 10506 7848
rect 10562 7792 10567 7848
rect 10428 7790 10567 7792
rect 12390 7850 12450 8334
rect 27153 8392 31267 8394
rect 27153 8336 27158 8392
rect 27214 8336 31206 8392
rect 31262 8336 31267 8392
rect 27153 8334 31267 8336
rect 27153 8331 27219 8334
rect 31201 8331 31267 8334
rect 26969 8258 27035 8261
rect 28257 8258 28323 8261
rect 26969 8256 28323 8258
rect 26969 8200 26974 8256
rect 27030 8200 28262 8256
rect 28318 8200 28323 8256
rect 26969 8198 28323 8200
rect 26969 8195 27035 8198
rect 28257 8195 28323 8198
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 29177 7850 29243 7853
rect 12390 7848 29243 7850
rect 12390 7792 29182 7848
rect 29238 7792 29243 7848
rect 12390 7790 29243 7792
rect 10428 7788 10434 7790
rect 10501 7787 10567 7790
rect 29177 7787 29243 7790
rect 5441 7714 5507 7717
rect 9581 7714 9647 7717
rect 5441 7712 9647 7714
rect 5441 7656 5446 7712
rect 5502 7656 9586 7712
rect 9642 7656 9647 7712
rect 5441 7654 9647 7656
rect 5441 7651 5507 7654
rect 9581 7651 9647 7654
rect 10041 7714 10107 7717
rect 13077 7714 13143 7717
rect 10041 7712 13143 7714
rect 10041 7656 10046 7712
rect 10102 7656 13082 7712
rect 13138 7656 13143 7712
rect 10041 7654 13143 7656
rect 10041 7651 10107 7654
rect 13077 7651 13143 7654
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 4889 7442 4955 7445
rect 12341 7442 12407 7445
rect 4889 7440 12407 7442
rect 4889 7384 4894 7440
rect 4950 7384 12346 7440
rect 12402 7384 12407 7440
rect 4889 7382 12407 7384
rect 4889 7379 4955 7382
rect 12341 7379 12407 7382
rect 4705 7306 4771 7309
rect 9397 7306 9463 7309
rect 4705 7304 9463 7306
rect 4705 7248 4710 7304
rect 4766 7248 9402 7304
rect 9458 7248 9463 7304
rect 4705 7246 9463 7248
rect 4705 7243 4771 7246
rect 9397 7243 9463 7246
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 9029 7034 9095 7037
rect 9397 7034 9463 7037
rect 9029 7032 9463 7034
rect 9029 6976 9034 7032
rect 9090 6976 9402 7032
rect 9458 6976 9463 7032
rect 9029 6974 9463 6976
rect 9029 6971 9095 6974
rect 9397 6971 9463 6974
rect 20110 6972 20116 7036
rect 20180 7034 20186 7036
rect 26877 7034 26943 7037
rect 20180 7032 26943 7034
rect 20180 6976 26882 7032
rect 26938 6976 26943 7032
rect 20180 6974 26943 6976
rect 20180 6972 20186 6974
rect 26877 6971 26943 6974
rect 2957 6898 3023 6901
rect 9397 6898 9463 6901
rect 2957 6896 9463 6898
rect 2957 6840 2962 6896
rect 3018 6840 9402 6896
rect 9458 6840 9463 6896
rect 2957 6838 9463 6840
rect 2957 6835 3023 6838
rect 9397 6835 9463 6838
rect 12341 6898 12407 6901
rect 13445 6898 13511 6901
rect 12341 6896 13511 6898
rect 12341 6840 12346 6896
rect 12402 6840 13450 6896
rect 13506 6840 13511 6896
rect 12341 6838 13511 6840
rect 12341 6835 12407 6838
rect 13445 6835 13511 6838
rect 3049 6762 3115 6765
rect 5993 6762 6059 6765
rect 3049 6760 6059 6762
rect 3049 6704 3054 6760
rect 3110 6704 5998 6760
rect 6054 6704 6059 6760
rect 3049 6702 6059 6704
rect 3049 6699 3115 6702
rect 5993 6699 6059 6702
rect 6545 6762 6611 6765
rect 7557 6762 7623 6765
rect 6545 6760 7623 6762
rect 6545 6704 6550 6760
rect 6606 6704 7562 6760
rect 7618 6704 7623 6760
rect 6545 6702 7623 6704
rect 6545 6699 6611 6702
rect 7557 6699 7623 6702
rect 24761 6762 24827 6765
rect 27245 6762 27311 6765
rect 24761 6760 27311 6762
rect 24761 6704 24766 6760
rect 24822 6704 27250 6760
rect 27306 6704 27311 6760
rect 24761 6702 27311 6704
rect 24761 6699 24827 6702
rect 27245 6699 27311 6702
rect 9489 6628 9555 6629
rect 9438 6564 9444 6628
rect 9508 6626 9555 6628
rect 9508 6624 9600 6626
rect 9550 6568 9600 6624
rect 9508 6566 9600 6568
rect 9508 6564 9555 6566
rect 9489 6563 9555 6564
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 5533 6490 5599 6493
rect 6453 6490 6519 6493
rect 5533 6488 6519 6490
rect 5533 6432 5538 6488
rect 5594 6432 6458 6488
rect 6514 6432 6519 6488
rect 5533 6430 6519 6432
rect 5533 6427 5599 6430
rect 6453 6427 6519 6430
rect 8477 6490 8543 6493
rect 17217 6490 17283 6493
rect 8477 6488 17283 6490
rect 8477 6432 8482 6488
rect 8538 6432 17222 6488
rect 17278 6432 17283 6488
rect 8477 6430 17283 6432
rect 8477 6427 8543 6430
rect 17217 6427 17283 6430
rect 5073 6354 5139 6357
rect 7373 6354 7439 6357
rect 5073 6352 7439 6354
rect 5073 6296 5078 6352
rect 5134 6296 7378 6352
rect 7434 6296 7439 6352
rect 5073 6294 7439 6296
rect 5073 6291 5139 6294
rect 7373 6291 7439 6294
rect 8661 6354 8727 6357
rect 12341 6354 12407 6357
rect 14181 6354 14247 6357
rect 8661 6352 11162 6354
rect 8661 6296 8666 6352
rect 8722 6296 11162 6352
rect 8661 6294 11162 6296
rect 8661 6291 8727 6294
rect 3049 6218 3115 6221
rect 10869 6218 10935 6221
rect 3049 6216 10935 6218
rect 3049 6160 3054 6216
rect 3110 6160 10874 6216
rect 10930 6160 10935 6216
rect 3049 6158 10935 6160
rect 11102 6218 11162 6294
rect 12341 6352 14247 6354
rect 12341 6296 12346 6352
rect 12402 6296 14186 6352
rect 14242 6296 14247 6352
rect 12341 6294 14247 6296
rect 12341 6291 12407 6294
rect 14181 6291 14247 6294
rect 22645 6354 22711 6357
rect 30414 6354 30420 6356
rect 22645 6352 30420 6354
rect 22645 6296 22650 6352
rect 22706 6296 30420 6352
rect 22645 6294 30420 6296
rect 22645 6291 22711 6294
rect 30414 6292 30420 6294
rect 30484 6292 30490 6356
rect 12433 6218 12499 6221
rect 11102 6216 12499 6218
rect 11102 6160 12438 6216
rect 12494 6160 12499 6216
rect 11102 6158 12499 6160
rect 3049 6155 3115 6158
rect 10869 6155 10935 6158
rect 12433 6155 12499 6158
rect 15009 6218 15075 6221
rect 19241 6218 19307 6221
rect 15009 6216 19307 6218
rect 15009 6160 15014 6216
rect 15070 6160 19246 6216
rect 19302 6160 19307 6216
rect 15009 6158 19307 6160
rect 15009 6155 15075 6158
rect 19241 6155 19307 6158
rect 20437 6218 20503 6221
rect 24710 6218 24716 6220
rect 20437 6216 24716 6218
rect 20437 6160 20442 6216
rect 20498 6160 24716 6216
rect 20437 6158 24716 6160
rect 20437 6155 20503 6158
rect 24710 6156 24716 6158
rect 24780 6156 24786 6220
rect 25497 6218 25563 6221
rect 25865 6218 25931 6221
rect 25497 6216 25931 6218
rect 25497 6160 25502 6216
rect 25558 6160 25870 6216
rect 25926 6160 25931 6216
rect 25497 6158 25931 6160
rect 25497 6155 25563 6158
rect 25865 6155 25931 6158
rect 8201 6082 8267 6085
rect 12341 6082 12407 6085
rect 8201 6080 12407 6082
rect 8201 6024 8206 6080
rect 8262 6024 12346 6080
rect 12402 6024 12407 6080
rect 8201 6022 12407 6024
rect 8201 6019 8267 6022
rect 12341 6019 12407 6022
rect 19977 6082 20043 6085
rect 23381 6082 23447 6085
rect 19977 6080 23447 6082
rect 19977 6024 19982 6080
rect 20038 6024 23386 6080
rect 23442 6024 23447 6080
rect 19977 6022 23447 6024
rect 19977 6019 20043 6022
rect 23381 6019 23447 6022
rect 24526 6020 24532 6084
rect 24596 6082 24602 6084
rect 31661 6082 31727 6085
rect 24596 6080 31727 6082
rect 24596 6024 31666 6080
rect 31722 6024 31727 6080
rect 24596 6022 31727 6024
rect 24596 6020 24602 6022
rect 31661 6019 31727 6022
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 8017 5946 8083 5949
rect 17125 5946 17191 5949
rect 8017 5944 17191 5946
rect 8017 5888 8022 5944
rect 8078 5888 17130 5944
rect 17186 5888 17191 5944
rect 8017 5886 17191 5888
rect 8017 5883 8083 5886
rect 17125 5883 17191 5886
rect 17769 5946 17835 5949
rect 22369 5946 22435 5949
rect 17769 5944 22435 5946
rect 17769 5888 17774 5944
rect 17830 5888 22374 5944
rect 22430 5888 22435 5944
rect 17769 5886 22435 5888
rect 17769 5883 17835 5886
rect 22369 5883 22435 5886
rect 24761 5946 24827 5949
rect 26877 5946 26943 5949
rect 24761 5944 26943 5946
rect 24761 5888 24766 5944
rect 24822 5888 26882 5944
rect 26938 5888 26943 5944
rect 24761 5886 26943 5888
rect 24761 5883 24827 5886
rect 26877 5883 26943 5886
rect 2957 5810 3023 5813
rect 5257 5810 5323 5813
rect 2957 5808 5323 5810
rect 2957 5752 2962 5808
rect 3018 5752 5262 5808
rect 5318 5752 5323 5808
rect 2957 5750 5323 5752
rect 2957 5747 3023 5750
rect 5257 5747 5323 5750
rect 8937 5810 9003 5813
rect 9765 5810 9831 5813
rect 8937 5808 9831 5810
rect 8937 5752 8942 5808
rect 8998 5752 9770 5808
rect 9826 5752 9831 5808
rect 8937 5750 9831 5752
rect 8937 5747 9003 5750
rect 9765 5747 9831 5750
rect 10317 5810 10383 5813
rect 11237 5810 11303 5813
rect 10317 5808 11303 5810
rect 10317 5752 10322 5808
rect 10378 5752 11242 5808
rect 11298 5752 11303 5808
rect 10317 5750 11303 5752
rect 10317 5747 10383 5750
rect 11237 5747 11303 5750
rect 21909 5810 21975 5813
rect 28349 5810 28415 5813
rect 21909 5808 28415 5810
rect 21909 5752 21914 5808
rect 21970 5752 28354 5808
rect 28410 5752 28415 5808
rect 21909 5750 28415 5752
rect 21909 5747 21975 5750
rect 28349 5747 28415 5750
rect 29729 5810 29795 5813
rect 32765 5810 32831 5813
rect 29729 5808 32831 5810
rect 29729 5752 29734 5808
rect 29790 5752 32770 5808
rect 32826 5752 32831 5808
rect 29729 5750 32831 5752
rect 29729 5747 29795 5750
rect 32765 5747 32831 5750
rect 2681 5674 2747 5677
rect 2865 5674 2931 5677
rect 2681 5672 2931 5674
rect 2681 5616 2686 5672
rect 2742 5616 2870 5672
rect 2926 5616 2931 5672
rect 2681 5614 2931 5616
rect 2681 5611 2747 5614
rect 2865 5611 2931 5614
rect 3601 5674 3667 5677
rect 8201 5674 8267 5677
rect 3601 5672 8267 5674
rect 3601 5616 3606 5672
rect 3662 5616 8206 5672
rect 8262 5616 8267 5672
rect 3601 5614 8267 5616
rect 3601 5611 3667 5614
rect 8201 5611 8267 5614
rect 9857 5674 9923 5677
rect 12525 5674 12591 5677
rect 9857 5672 12591 5674
rect 9857 5616 9862 5672
rect 9918 5616 12530 5672
rect 12586 5616 12591 5672
rect 9857 5614 12591 5616
rect 9857 5611 9923 5614
rect 12525 5611 12591 5614
rect 13997 5674 14063 5677
rect 15929 5674 15995 5677
rect 13997 5672 15995 5674
rect 13997 5616 14002 5672
rect 14058 5616 15934 5672
rect 15990 5616 15995 5672
rect 13997 5614 15995 5616
rect 13997 5611 14063 5614
rect 15929 5611 15995 5614
rect 25446 5612 25452 5676
rect 25516 5674 25522 5676
rect 30925 5674 30991 5677
rect 25516 5672 30991 5674
rect 25516 5616 30930 5672
rect 30986 5616 30991 5672
rect 25516 5614 30991 5616
rect 25516 5612 25522 5614
rect 30925 5611 30991 5614
rect 2773 5538 2839 5541
rect 10409 5538 10475 5541
rect 2773 5536 10475 5538
rect 2773 5480 2778 5536
rect 2834 5480 10414 5536
rect 10470 5480 10475 5536
rect 2773 5478 10475 5480
rect 2773 5475 2839 5478
rect 10409 5475 10475 5478
rect 11881 5538 11947 5541
rect 12709 5538 12775 5541
rect 11881 5536 12775 5538
rect 11881 5480 11886 5536
rect 11942 5480 12714 5536
rect 12770 5480 12775 5536
rect 11881 5478 12775 5480
rect 11881 5475 11947 5478
rect 12709 5475 12775 5478
rect 24761 5538 24827 5541
rect 25405 5538 25471 5541
rect 24761 5536 25471 5538
rect 24761 5480 24766 5536
rect 24822 5480 25410 5536
rect 25466 5480 25471 5536
rect 24761 5478 25471 5480
rect 24761 5475 24827 5478
rect 25405 5475 25471 5478
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 2405 5402 2471 5405
rect 4613 5402 4679 5405
rect 8017 5402 8083 5405
rect 2405 5400 2790 5402
rect 2405 5344 2410 5400
rect 2466 5344 2790 5400
rect 2405 5342 2790 5344
rect 2405 5339 2471 5342
rect 2730 5130 2790 5342
rect 4613 5400 8083 5402
rect 4613 5344 4618 5400
rect 4674 5344 8022 5400
rect 8078 5344 8083 5400
rect 4613 5342 8083 5344
rect 4613 5339 4679 5342
rect 8017 5339 8083 5342
rect 9765 5402 9831 5405
rect 10501 5402 10567 5405
rect 9765 5400 10567 5402
rect 9765 5344 9770 5400
rect 9826 5344 10506 5400
rect 10562 5344 10567 5400
rect 9765 5342 10567 5344
rect 9765 5339 9831 5342
rect 10501 5339 10567 5342
rect 10685 5402 10751 5405
rect 10961 5402 11027 5405
rect 10685 5400 11027 5402
rect 10685 5344 10690 5400
rect 10746 5344 10966 5400
rect 11022 5344 11027 5400
rect 10685 5342 11027 5344
rect 10685 5339 10751 5342
rect 10961 5339 11027 5342
rect 11421 5402 11487 5405
rect 13353 5402 13419 5405
rect 11421 5400 13419 5402
rect 11421 5344 11426 5400
rect 11482 5344 13358 5400
rect 13414 5344 13419 5400
rect 11421 5342 13419 5344
rect 11421 5339 11487 5342
rect 13353 5339 13419 5342
rect 2865 5266 2931 5269
rect 5809 5266 5875 5269
rect 2865 5264 5875 5266
rect 2865 5208 2870 5264
rect 2926 5208 5814 5264
rect 5870 5208 5875 5264
rect 2865 5206 5875 5208
rect 2865 5203 2931 5206
rect 5809 5203 5875 5206
rect 6545 5266 6611 5269
rect 11329 5266 11395 5269
rect 6545 5264 11395 5266
rect 6545 5208 6550 5264
rect 6606 5208 11334 5264
rect 11390 5208 11395 5264
rect 6545 5206 11395 5208
rect 6545 5203 6611 5206
rect 11329 5203 11395 5206
rect 17769 5266 17835 5269
rect 27654 5266 27660 5268
rect 17769 5264 27660 5266
rect 17769 5208 17774 5264
rect 17830 5208 27660 5264
rect 17769 5206 27660 5208
rect 17769 5203 17835 5206
rect 27654 5204 27660 5206
rect 27724 5204 27730 5268
rect 11973 5130 12039 5133
rect 2730 5128 12039 5130
rect 2730 5072 11978 5128
rect 12034 5072 12039 5128
rect 2730 5070 12039 5072
rect 11973 5067 12039 5070
rect 20345 5130 20411 5133
rect 28809 5130 28875 5133
rect 20345 5128 28875 5130
rect 20345 5072 20350 5128
rect 20406 5072 28814 5128
rect 28870 5072 28875 5128
rect 20345 5070 28875 5072
rect 20345 5067 20411 5070
rect 28809 5067 28875 5070
rect 9673 4994 9739 4997
rect 10317 4994 10383 4997
rect 9673 4992 10383 4994
rect 9673 4936 9678 4992
rect 9734 4936 10322 4992
rect 10378 4936 10383 4992
rect 9673 4934 10383 4936
rect 9673 4931 9739 4934
rect 10317 4931 10383 4934
rect 19241 4994 19307 4997
rect 28942 4994 28948 4996
rect 19241 4992 28948 4994
rect 19241 4936 19246 4992
rect 19302 4936 28948 4992
rect 19241 4934 28948 4936
rect 19241 4931 19307 4934
rect 28942 4932 28948 4934
rect 29012 4932 29018 4996
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 9489 4858 9555 4861
rect 9949 4858 10015 4861
rect 9489 4856 10015 4858
rect 9489 4800 9494 4856
rect 9550 4800 9954 4856
rect 10010 4800 10015 4856
rect 9489 4798 10015 4800
rect 9489 4795 9555 4798
rect 9949 4795 10015 4798
rect 10225 4858 10291 4861
rect 12249 4858 12315 4861
rect 12525 4858 12591 4861
rect 10225 4856 12082 4858
rect 10225 4800 10230 4856
rect 10286 4800 12082 4856
rect 10225 4798 12082 4800
rect 10225 4795 10291 4798
rect 4153 4722 4219 4725
rect 11697 4722 11763 4725
rect 4153 4720 11763 4722
rect 4153 4664 4158 4720
rect 4214 4664 11702 4720
rect 11758 4664 11763 4720
rect 4153 4662 11763 4664
rect 12022 4722 12082 4798
rect 12249 4856 12591 4858
rect 12249 4800 12254 4856
rect 12310 4800 12530 4856
rect 12586 4800 12591 4856
rect 12249 4798 12591 4800
rect 12249 4795 12315 4798
rect 12525 4795 12591 4798
rect 18505 4858 18571 4861
rect 30598 4858 30604 4860
rect 18505 4856 30604 4858
rect 18505 4800 18510 4856
rect 18566 4800 30604 4856
rect 18505 4798 30604 4800
rect 18505 4795 18571 4798
rect 30598 4796 30604 4798
rect 30668 4796 30674 4860
rect 34605 4858 34671 4861
rect 34605 4856 34714 4858
rect 34605 4800 34610 4856
rect 34666 4800 34714 4856
rect 34605 4795 34714 4800
rect 14365 4722 14431 4725
rect 12022 4720 14431 4722
rect 12022 4664 14370 4720
rect 14426 4664 14431 4720
rect 12022 4662 14431 4664
rect 34654 4722 34714 4795
rect 34881 4722 34947 4725
rect 34654 4720 34947 4722
rect 34654 4664 34886 4720
rect 34942 4664 34947 4720
rect 34654 4662 34947 4664
rect 4153 4659 4219 4662
rect 11697 4659 11763 4662
rect 14365 4659 14431 4662
rect 34881 4659 34947 4662
rect 3877 4586 3943 4589
rect 10869 4586 10935 4589
rect 3877 4584 10935 4586
rect 3877 4528 3882 4584
rect 3938 4528 10874 4584
rect 10930 4528 10935 4584
rect 3877 4526 10935 4528
rect 3877 4523 3943 4526
rect 10869 4523 10935 4526
rect 32765 4586 32831 4589
rect 35709 4586 35775 4589
rect 32765 4584 35775 4586
rect 32765 4528 32770 4584
rect 32826 4528 35714 4584
rect 35770 4528 35775 4584
rect 32765 4526 35775 4528
rect 32765 4523 32831 4526
rect 35709 4523 35775 4526
rect 2589 4450 2655 4453
rect 10777 4450 10843 4453
rect 2589 4448 10843 4450
rect 2589 4392 2594 4448
rect 2650 4392 10782 4448
rect 10838 4392 10843 4448
rect 2589 4390 10843 4392
rect 2589 4387 2655 4390
rect 10777 4387 10843 4390
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 3601 4314 3667 4317
rect 4889 4314 4955 4317
rect 3601 4312 4955 4314
rect 3601 4256 3606 4312
rect 3662 4256 4894 4312
rect 4950 4256 4955 4312
rect 3601 4254 4955 4256
rect 3601 4251 3667 4254
rect 4889 4251 4955 4254
rect 9305 4314 9371 4317
rect 13905 4314 13971 4317
rect 9305 4312 13971 4314
rect 9305 4256 9310 4312
rect 9366 4256 13910 4312
rect 13966 4256 13971 4312
rect 9305 4254 13971 4256
rect 9305 4251 9371 4254
rect 13905 4251 13971 4254
rect 21449 4314 21515 4317
rect 25814 4314 25820 4316
rect 21449 4312 25820 4314
rect 21449 4256 21454 4312
rect 21510 4256 25820 4312
rect 21449 4254 25820 4256
rect 21449 4251 21515 4254
rect 25814 4252 25820 4254
rect 25884 4252 25890 4316
rect 3693 4178 3759 4181
rect 11513 4178 11579 4181
rect 3693 4176 11579 4178
rect 3693 4120 3698 4176
rect 3754 4120 11518 4176
rect 11574 4120 11579 4176
rect 3693 4118 11579 4120
rect 3693 4115 3759 4118
rect 11513 4115 11579 4118
rect 3785 4042 3851 4045
rect 9305 4042 9371 4045
rect 19425 4044 19491 4045
rect 19374 4042 19380 4044
rect 3785 4040 9371 4042
rect 3785 3984 3790 4040
rect 3846 3984 9310 4040
rect 9366 3984 9371 4040
rect 3785 3982 9371 3984
rect 19334 3982 19380 4042
rect 19444 4040 19491 4044
rect 19486 3984 19491 4040
rect 3785 3979 3851 3982
rect 9305 3979 9371 3982
rect 19374 3980 19380 3982
rect 19444 3980 19491 3984
rect 19425 3979 19491 3980
rect 19977 4042 20043 4045
rect 20110 4042 20116 4044
rect 19977 4040 20116 4042
rect 19977 3984 19982 4040
rect 20038 3984 20116 4040
rect 19977 3982 20116 3984
rect 19977 3979 20043 3982
rect 20110 3980 20116 3982
rect 20180 3980 20186 4044
rect 25313 4042 25379 4045
rect 25446 4042 25452 4044
rect 25313 4040 25452 4042
rect 25313 3984 25318 4040
rect 25374 3984 25452 4040
rect 25313 3982 25452 3984
rect 25313 3979 25379 3982
rect 25446 3980 25452 3982
rect 25516 3980 25522 4044
rect 19517 3906 19583 3909
rect 20437 3906 20503 3909
rect 19517 3904 20503 3906
rect 19517 3848 19522 3904
rect 19578 3848 20442 3904
rect 20498 3848 20503 3904
rect 19517 3846 20503 3848
rect 19517 3843 19583 3846
rect 20437 3843 20503 3846
rect 21909 3906 21975 3909
rect 22093 3906 22159 3909
rect 21909 3904 22159 3906
rect 21909 3848 21914 3904
rect 21970 3848 22098 3904
rect 22154 3848 22159 3904
rect 21909 3846 22159 3848
rect 21909 3843 21975 3846
rect 22093 3843 22159 3846
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 10358 3770 10364 3772
rect 4662 3710 10364 3770
rect 3693 3634 3759 3637
rect 4662 3634 4722 3710
rect 10358 3708 10364 3710
rect 10428 3708 10434 3772
rect 3693 3632 4722 3634
rect 3693 3576 3698 3632
rect 3754 3576 4722 3632
rect 3693 3574 4722 3576
rect 5257 3634 5323 3637
rect 8293 3634 8359 3637
rect 5257 3632 8359 3634
rect 5257 3576 5262 3632
rect 5318 3576 8298 3632
rect 8354 3576 8359 3632
rect 5257 3574 8359 3576
rect 3693 3571 3759 3574
rect 5257 3571 5323 3574
rect 8293 3571 8359 3574
rect 9397 3634 9463 3637
rect 13077 3634 13143 3637
rect 9397 3632 13143 3634
rect 9397 3576 9402 3632
rect 9458 3576 13082 3632
rect 13138 3576 13143 3632
rect 9397 3574 13143 3576
rect 9397 3571 9463 3574
rect 13077 3571 13143 3574
rect 3233 3498 3299 3501
rect 10409 3498 10475 3501
rect 3233 3496 10475 3498
rect 3233 3440 3238 3496
rect 3294 3440 10414 3496
rect 10470 3440 10475 3496
rect 3233 3438 10475 3440
rect 3233 3435 3299 3438
rect 10409 3435 10475 3438
rect 2957 3362 3023 3365
rect 10961 3362 11027 3365
rect 2957 3360 11027 3362
rect 2957 3304 2962 3360
rect 3018 3304 10966 3360
rect 11022 3304 11027 3360
rect 2957 3302 11027 3304
rect 2957 3299 3023 3302
rect 10961 3299 11027 3302
rect 12157 3362 12223 3365
rect 15377 3362 15443 3365
rect 12157 3360 15443 3362
rect 12157 3304 12162 3360
rect 12218 3304 15382 3360
rect 15438 3304 15443 3360
rect 12157 3302 15443 3304
rect 12157 3299 12223 3302
rect 15377 3299 15443 3302
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 2865 3226 2931 3229
rect 12157 3226 12223 3229
rect 29126 3226 29132 3228
rect 2865 3224 12223 3226
rect 2865 3168 2870 3224
rect 2926 3168 12162 3224
rect 12218 3168 12223 3224
rect 2865 3166 12223 3168
rect 2865 3163 2931 3166
rect 12157 3163 12223 3166
rect 22050 3166 29132 3226
rect 4245 3090 4311 3093
rect 9581 3090 9647 3093
rect 4245 3088 9647 3090
rect 4245 3032 4250 3088
rect 4306 3032 9586 3088
rect 9642 3032 9647 3088
rect 4245 3030 9647 3032
rect 4245 3027 4311 3030
rect 9581 3027 9647 3030
rect 10041 3090 10107 3093
rect 13905 3090 13971 3093
rect 10041 3088 13971 3090
rect 10041 3032 10046 3088
rect 10102 3032 13910 3088
rect 13966 3032 13971 3088
rect 10041 3030 13971 3032
rect 10041 3027 10107 3030
rect 13905 3027 13971 3030
rect 17534 3028 17540 3092
rect 17604 3090 17610 3092
rect 17953 3090 18019 3093
rect 17604 3088 18019 3090
rect 17604 3032 17958 3088
rect 18014 3032 18019 3088
rect 17604 3030 18019 3032
rect 17604 3028 17610 3030
rect 17953 3027 18019 3030
rect 18229 3090 18295 3093
rect 22050 3090 22110 3166
rect 29126 3164 29132 3166
rect 29196 3164 29202 3228
rect 24485 3092 24551 3093
rect 24485 3090 24532 3092
rect 18229 3088 22110 3090
rect 18229 3032 18234 3088
rect 18290 3032 22110 3088
rect 18229 3030 22110 3032
rect 24440 3088 24532 3090
rect 24440 3032 24490 3088
rect 24440 3030 24532 3032
rect 18229 3027 18295 3030
rect 24485 3028 24532 3030
rect 24596 3028 24602 3092
rect 24485 3027 24551 3028
rect 3417 2954 3483 2957
rect 8201 2954 8267 2957
rect 3417 2952 8267 2954
rect 3417 2896 3422 2952
rect 3478 2896 8206 2952
rect 8262 2896 8267 2952
rect 3417 2894 8267 2896
rect 3417 2891 3483 2894
rect 8201 2891 8267 2894
rect 4613 2818 4679 2821
rect 10225 2818 10291 2821
rect 4613 2816 10291 2818
rect 4613 2760 4618 2816
rect 4674 2760 10230 2816
rect 10286 2760 10291 2816
rect 4613 2758 10291 2760
rect 4613 2755 4679 2758
rect 10225 2755 10291 2758
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 6913 2682 6979 2685
rect 10777 2682 10843 2685
rect 6913 2680 10843 2682
rect 6913 2624 6918 2680
rect 6974 2624 10782 2680
rect 10838 2624 10843 2680
rect 6913 2622 10843 2624
rect 6913 2619 6979 2622
rect 10777 2619 10843 2622
rect 3049 2546 3115 2549
rect 8753 2546 8819 2549
rect 3049 2544 8819 2546
rect 3049 2488 3054 2544
rect 3110 2488 8758 2544
rect 8814 2488 8819 2544
rect 3049 2486 8819 2488
rect 3049 2483 3115 2486
rect 8753 2483 8819 2486
rect 8201 2410 8267 2413
rect 9305 2410 9371 2413
rect 8201 2408 9371 2410
rect 8201 2352 8206 2408
rect 8262 2352 9310 2408
rect 9366 2352 9371 2408
rect 8201 2350 9371 2352
rect 8201 2347 8267 2350
rect 9305 2347 9371 2350
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19380 19756 19444 19820
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 20300 16900 20364 16964
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 17540 16008 17604 16012
rect 17540 15952 17554 16008
rect 17554 15952 17604 16008
rect 17540 15948 17604 15952
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19380 15268 19444 15332
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 20300 11928 20364 11932
rect 20300 11872 20314 11928
rect 20314 11872 20364 11928
rect 20300 11868 20364 11872
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 25820 11052 25884 11116
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 29132 10160 29196 10164
rect 29132 10104 29182 10160
rect 29182 10104 29196 10160
rect 29132 10100 29196 10104
rect 28948 9964 29012 10028
rect 24716 9828 24780 9892
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 27660 9692 27724 9756
rect 30420 9692 30484 9756
rect 19380 9420 19444 9484
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 30604 9012 30668 9076
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 9444 8664 9508 8668
rect 9444 8608 9494 8664
rect 9494 8608 9508 8664
rect 9444 8604 9508 8608
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 10364 7788 10428 7852
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 20116 6972 20180 7036
rect 9444 6624 9508 6628
rect 9444 6568 9494 6624
rect 9494 6568 9508 6624
rect 9444 6564 9508 6568
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 30420 6292 30484 6356
rect 24716 6156 24780 6220
rect 24532 6020 24596 6084
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 25452 5612 25516 5676
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 27660 5204 27724 5268
rect 28948 4932 29012 4996
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 30604 4796 30668 4860
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 25820 4252 25884 4316
rect 19380 4040 19444 4044
rect 19380 3984 19430 4040
rect 19430 3984 19444 4040
rect 19380 3980 19444 3984
rect 20116 3980 20180 4044
rect 25452 3980 25516 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 10364 3708 10428 3772
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 17540 3028 17604 3092
rect 29132 3164 29196 3228
rect 24532 3088 24596 3092
rect 24532 3032 24546 3088
rect 24546 3032 24596 3088
rect 24532 3028 24596 3032
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19379 19820 19445 19821
rect 19379 19756 19380 19820
rect 19444 19756 19445 19820
rect 19379 19755 19445 19756
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 17539 16012 17605 16013
rect 17539 15948 17540 16012
rect 17604 15948 17605 16012
rect 17539 15947 17605 15948
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 9443 8668 9509 8669
rect 9443 8604 9444 8668
rect 9508 8604 9509 8668
rect 9443 8603 9509 8604
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 9446 6629 9506 8603
rect 10363 7852 10429 7853
rect 10363 7788 10364 7852
rect 10428 7788 10429 7852
rect 10363 7787 10429 7788
rect 9443 6628 9509 6629
rect 9443 6564 9444 6628
rect 9508 6564 9509 6628
rect 9443 6563 9509 6564
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 10366 3773 10426 7787
rect 10363 3772 10429 3773
rect 10363 3708 10364 3772
rect 10428 3708 10429 3772
rect 10363 3707 10429 3708
rect 17542 3093 17602 15947
rect 19382 15333 19442 19755
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 20299 16964 20365 16965
rect 20299 16900 20300 16964
rect 20364 16900 20365 16964
rect 20299 16899 20365 16900
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19379 15332 19445 15333
rect 19379 15268 19380 15332
rect 19444 15268 19445 15332
rect 19379 15267 19445 15268
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 20302 11933 20362 16899
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 20299 11932 20365 11933
rect 20299 11868 20300 11932
rect 20364 11868 20365 11932
rect 20299 11867 20365 11868
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 25819 11116 25885 11117
rect 25819 11052 25820 11116
rect 25884 11052 25885 11116
rect 25819 11051 25885 11052
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 24715 9892 24781 9893
rect 24715 9828 24716 9892
rect 24780 9828 24781 9892
rect 24715 9827 24781 9828
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19379 9484 19445 9485
rect 19379 9420 19380 9484
rect 19444 9420 19445 9484
rect 19379 9419 19445 9420
rect 19382 4045 19442 9419
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 20115 7036 20181 7037
rect 20115 6972 20116 7036
rect 20180 6972 20181 7036
rect 20115 6971 20181 6972
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19379 4044 19445 4045
rect 19379 3980 19380 4044
rect 19444 3980 19445 4044
rect 19379 3979 19445 3980
rect 19568 3296 19888 4320
rect 20118 4045 20178 6971
rect 24718 6221 24778 9827
rect 24715 6220 24781 6221
rect 24715 6156 24716 6220
rect 24780 6156 24781 6220
rect 24715 6155 24781 6156
rect 24531 6084 24597 6085
rect 24531 6020 24532 6084
rect 24596 6020 24597 6084
rect 24531 6019 24597 6020
rect 20115 4044 20181 4045
rect 20115 3980 20116 4044
rect 20180 3980 20181 4044
rect 20115 3979 20181 3980
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 17539 3092 17605 3093
rect 17539 3028 17540 3092
rect 17604 3028 17605 3092
rect 17539 3027 17605 3028
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 2208 19888 3232
rect 24534 3093 24594 6019
rect 25451 5676 25517 5677
rect 25451 5612 25452 5676
rect 25516 5612 25517 5676
rect 25451 5611 25517 5612
rect 25454 4045 25514 5611
rect 25822 4317 25882 11051
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 29131 10164 29197 10165
rect 29131 10100 29132 10164
rect 29196 10100 29197 10164
rect 29131 10099 29197 10100
rect 28947 10028 29013 10029
rect 28947 9964 28948 10028
rect 29012 9964 29013 10028
rect 28947 9963 29013 9964
rect 27659 9756 27725 9757
rect 27659 9692 27660 9756
rect 27724 9692 27725 9756
rect 27659 9691 27725 9692
rect 27662 5269 27722 9691
rect 27659 5268 27725 5269
rect 27659 5204 27660 5268
rect 27724 5204 27725 5268
rect 27659 5203 27725 5204
rect 28950 4997 29010 9963
rect 28947 4996 29013 4997
rect 28947 4932 28948 4996
rect 29012 4932 29013 4996
rect 28947 4931 29013 4932
rect 25819 4316 25885 4317
rect 25819 4252 25820 4316
rect 25884 4252 25885 4316
rect 25819 4251 25885 4252
rect 25451 4044 25517 4045
rect 25451 3980 25452 4044
rect 25516 3980 25517 4044
rect 25451 3979 25517 3980
rect 29134 3229 29194 10099
rect 30419 9756 30485 9757
rect 30419 9692 30420 9756
rect 30484 9692 30485 9756
rect 30419 9691 30485 9692
rect 30422 6357 30482 9691
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 30603 9076 30669 9077
rect 30603 9012 30604 9076
rect 30668 9012 30669 9076
rect 30603 9011 30669 9012
rect 30419 6356 30485 6357
rect 30419 6292 30420 6356
rect 30484 6292 30485 6356
rect 30419 6291 30485 6292
rect 30606 4861 30666 9011
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 30603 4860 30669 4861
rect 30603 4796 30604 4860
rect 30668 4796 30669 4860
rect 30603 4795 30669 4796
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 29131 3228 29197 3229
rect 29131 3164 29132 3228
rect 29196 3164 29197 3228
rect 29131 3163 29197 3164
rect 24531 3092 24597 3093
rect 24531 3028 24532 3092
rect 24596 3028 24597 3092
rect 24531 3027 24597 3028
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 2852 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform -1 0 2300 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform -1 0 2208 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform 1 0 17756 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 2576 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2300 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33
timestamp 1644511149
transform 1 0 4140 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49
timestamp 1644511149
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1644511149
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64
timestamp 1644511149
transform 1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71
timestamp 1644511149
transform 1 0 7636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_92
timestamp 1644511149
transform 1 0 9568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101
timestamp 1644511149
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1644511149
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1644511149
transform 1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_124
timestamp 1644511149
transform 1 0 12512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_130 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13064 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp 1644511149
transform 1 0 14996 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_162
timestamp 1644511149
transform 1 0 16008 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_186
timestamp 1644511149
transform 1 0 18216 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1644511149
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_201
timestamp 1644511149
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1644511149
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_236
timestamp 1644511149
transform 1 0 22816 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1644511149
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_257
timestamp 1644511149
transform 1 0 24748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_263
timestamp 1644511149
transform 1 0 25300 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_269
timestamp 1644511149
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1644511149
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_285
timestamp 1644511149
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_292
timestamp 1644511149
transform 1 0 27968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1644511149
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1644511149
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_313
timestamp 1644511149
transform 1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_329
timestamp 1644511149
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1644511149
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_341
timestamp 1644511149
transform 1 0 32476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1644511149
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1644511149
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_369
timestamp 1644511149
transform 1 0 35052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1644511149
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_397
timestamp 1644511149
transform 1 0 37628 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1644511149
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_10
timestamp 1644511149
transform 1 0 2024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_17
timestamp 1644511149
transform 1 0 2668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_24
timestamp 1644511149
transform 1 0 3312 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_31
timestamp 1644511149
transform 1 0 3956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_38
timestamp 1644511149
transform 1 0 4600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45
timestamp 1644511149
transform 1 0 5244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_76
timestamp 1644511149
transform 1 0 8096 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_94
timestamp 1644511149
transform 1 0 9752 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1644511149
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_129
timestamp 1644511149
transform 1 0 12972 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_140
timestamp 1644511149
transform 1 0 13984 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_146
timestamp 1644511149
transform 1 0 14536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_157
timestamp 1644511149
transform 1 0 15548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1644511149
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_179
timestamp 1644511149
transform 1 0 17572 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_190
timestamp 1644511149
transform 1 0 18584 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_198
timestamp 1644511149
transform 1 0 19320 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_205
timestamp 1644511149
transform 1 0 19964 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_214
timestamp 1644511149
transform 1 0 20792 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1644511149
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_232
timestamp 1644511149
transform 1 0 22448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_241
timestamp 1644511149
transform 1 0 23276 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_255
timestamp 1644511149
transform 1 0 24564 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_269
timestamp 1644511149
transform 1 0 25852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_291
timestamp 1644511149
transform 1 0 27876 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_302
timestamp 1644511149
transform 1 0 28888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_311
timestamp 1644511149
transform 1 0 29716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_331
timestamp 1644511149
transform 1 0 31556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_341
timestamp 1644511149
transform 1 0 32476 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_349
timestamp 1644511149
transform 1 0 33212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_360
timestamp 1644511149
transform 1 0 34224 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_368
timestamp 1644511149
transform 1 0 34960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_377
timestamp 1644511149
transform 1 0 35788 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_386
timestamp 1644511149
transform 1 0 36616 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_397
timestamp 1644511149
transform 1 0 37628 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_10
timestamp 1644511149
transform 1 0 2024 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_17
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_61
timestamp 1644511149
transform 1 0 6716 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_72
timestamp 1644511149
transform 1 0 7728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_76
timestamp 1644511149
transform 1 0 8096 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1644511149
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_108
timestamp 1644511149
transform 1 0 11040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_119
timestamp 1644511149
transform 1 0 12052 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_127
timestamp 1644511149
transform 1 0 12788 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1644511149
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_145
timestamp 1644511149
transform 1 0 14444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_165
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_172
timestamp 1644511149
transform 1 0 16928 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1644511149
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_202
timestamp 1644511149
transform 1 0 19688 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_210
timestamp 1644511149
transform 1 0 20424 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_218
timestamp 1644511149
transform 1 0 21160 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_222
timestamp 1644511149
transform 1 0 21528 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_228
timestamp 1644511149
transform 1 0 22080 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1644511149
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_258
timestamp 1644511149
transform 1 0 24840 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_264
timestamp 1644511149
transform 1 0 25392 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_271
timestamp 1644511149
transform 1 0 26036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_279
timestamp 1644511149
transform 1 0 26772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_299
timestamp 1644511149
transform 1 0 28612 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_327
timestamp 1644511149
transform 1 0 31188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_336
timestamp 1644511149
transform 1 0 32016 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_354
timestamp 1644511149
transform 1 0 33672 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_362
timestamp 1644511149
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_381
timestamp 1644511149
transform 1 0 36156 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_390
timestamp 1644511149
transform 1 0 36984 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_396
timestamp 1644511149
transform 1 0 37536 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_12
timestamp 1644511149
transform 1 0 2208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_19
timestamp 1644511149
transform 1 0 2852 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_26
timestamp 1644511149
transform 1 0 3496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_46
timestamp 1644511149
transform 1 0 5336 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1644511149
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_64
timestamp 1644511149
transform 1 0 6992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_84
timestamp 1644511149
transform 1 0 8832 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1644511149
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1644511149
transform 1 0 13248 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_152
timestamp 1644511149
transform 1 0 15088 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_163
timestamp 1644511149
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_190
timestamp 1644511149
transform 1 0 18584 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_196
timestamp 1644511149
transform 1 0 19136 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_204
timestamp 1644511149
transform 1 0 19872 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_213
timestamp 1644511149
transform 1 0 20700 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1644511149
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_241
timestamp 1644511149
transform 1 0 23276 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_253
timestamp 1644511149
transform 1 0 24380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_259
timestamp 1644511149
transform 1 0 24932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_266
timestamp 1644511149
transform 1 0 25576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_275
timestamp 1644511149
transform 1 0 26404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_297
timestamp 1644511149
transform 1 0 28428 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_311
timestamp 1644511149
transform 1 0 29716 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_321
timestamp 1644511149
transform 1 0 30636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_331
timestamp 1644511149
transform 1 0 31556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_353
timestamp 1644511149
transform 1 0 33580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_378
timestamp 1644511149
transform 1 0 35880 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_387
timestamp 1644511149
transform 1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_403
timestamp 1644511149
transform 1 0 38180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_10
timestamp 1644511149
transform 1 0 2024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_17
timestamp 1644511149
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1644511149
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_36
timestamp 1644511149
transform 1 0 4416 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_47
timestamp 1644511149
transform 1 0 5428 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_67
timestamp 1644511149
transform 1 0 7268 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_78
timestamp 1644511149
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_90
timestamp 1644511149
transform 1 0 9384 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_117
timestamp 1644511149
transform 1 0 11868 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_124
timestamp 1644511149
transform 1 0 12512 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1644511149
transform 1 0 14720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_168
timestamp 1644511149
transform 1 0 16560 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_182
timestamp 1644511149
transform 1 0 17848 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_191
timestamp 1644511149
transform 1 0 18676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_205
timestamp 1644511149
transform 1 0 19964 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_213
timestamp 1644511149
transform 1 0 20700 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_228
timestamp 1644511149
transform 1 0 22080 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_236
timestamp 1644511149
transform 1 0 22816 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_244
timestamp 1644511149
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_257
timestamp 1644511149
transform 1 0 24748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_278
timestamp 1644511149
transform 1 0 26680 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_286
timestamp 1644511149
transform 1 0 27416 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_294
timestamp 1644511149
transform 1 0 28152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1644511149
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_314
timestamp 1644511149
transform 1 0 29992 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_332
timestamp 1644511149
transform 1 0 31648 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_341
timestamp 1644511149
transform 1 0 32476 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_350
timestamp 1644511149
transform 1 0 33304 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_370
timestamp 1644511149
transform 1 0 35144 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_384
timestamp 1644511149
transform 1 0 36432 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_391
timestamp 1644511149
transform 1 0 37076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_403
timestamp 1644511149
transform 1 0 38180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_9
timestamp 1644511149
transform 1 0 1932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_16
timestamp 1644511149
transform 1 0 2576 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_23
timestamp 1644511149
transform 1 0 3220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_43
timestamp 1644511149
transform 1 0 5060 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_50
timestamp 1644511149
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_62
timestamp 1644511149
transform 1 0 6808 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_74
timestamp 1644511149
transform 1 0 7912 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_85
timestamp 1644511149
transform 1 0 8924 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_96
timestamp 1644511149
transform 1 0 9936 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp 1644511149
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_118
timestamp 1644511149
transform 1 0 11960 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_126
timestamp 1644511149
transform 1 0 12696 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_130
timestamp 1644511149
transform 1 0 13064 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_139
timestamp 1644511149
transform 1 0 13892 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_147
timestamp 1644511149
transform 1 0 14628 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_154
timestamp 1644511149
transform 1 0 15272 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_163
timestamp 1644511149
transform 1 0 16100 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_178
timestamp 1644511149
transform 1 0 17480 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_184
timestamp 1644511149
transform 1 0 18032 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_190
timestamp 1644511149
transform 1 0 18584 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_215
timestamp 1644511149
transform 1 0 20884 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_229
timestamp 1644511149
transform 1 0 22172 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_257
timestamp 1644511149
transform 1 0 24748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_268
timestamp 1644511149
transform 1 0 25760 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_275
timestamp 1644511149
transform 1 0 26404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_284
timestamp 1644511149
transform 1 0 27232 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_291
timestamp 1644511149
transform 1 0 27876 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_299
timestamp 1644511149
transform 1 0 28612 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_306
timestamp 1644511149
transform 1 0 29256 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_313
timestamp 1644511149
transform 1 0 29900 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_324
timestamp 1644511149
transform 1 0 30912 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_331
timestamp 1644511149
transform 1 0 31556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_341
timestamp 1644511149
transform 1 0 32476 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_346
timestamp 1644511149
transform 1 0 32936 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_353
timestamp 1644511149
transform 1 0 33580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_367
timestamp 1644511149
transform 1 0 34868 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_374
timestamp 1644511149
transform 1 0 35512 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_381
timestamp 1644511149
transform 1 0 36156 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1644511149
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_403
timestamp 1644511149
transform 1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_8
timestamp 1644511149
transform 1 0 1840 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_12
timestamp 1644511149
transform 1 0 2208 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_17
timestamp 1644511149
transform 1 0 2668 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1644511149
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_38
timestamp 1644511149
transform 1 0 4600 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_46
timestamp 1644511149
transform 1 0 5336 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_51
timestamp 1644511149
transform 1 0 5796 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_60
timestamp 1644511149
transform 1 0 6624 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_64
timestamp 1644511149
transform 1 0 6992 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_69
timestamp 1644511149
transform 1 0 7452 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_104
timestamp 1644511149
transform 1 0 10672 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_111
timestamp 1644511149
transform 1 0 11316 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_125
timestamp 1644511149
transform 1 0 12604 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_129
timestamp 1644511149
transform 1 0 12972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1644511149
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_146
timestamp 1644511149
transform 1 0 14536 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1644511149
transform 1 0 15088 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_159
timestamp 1644511149
transform 1 0 15732 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_163
timestamp 1644511149
transform 1 0 16100 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_170
timestamp 1644511149
transform 1 0 16744 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_179
timestamp 1644511149
transform 1 0 17572 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_183
timestamp 1644511149
transform 1 0 17940 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1644511149
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_205
timestamp 1644511149
transform 1 0 19964 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_212
timestamp 1644511149
transform 1 0 20608 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_223
timestamp 1644511149
transform 1 0 21620 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_227
timestamp 1644511149
transform 1 0 21988 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_235
timestamp 1644511149
transform 1 0 22724 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp 1644511149
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_258
timestamp 1644511149
transform 1 0 24840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_278
timestamp 1644511149
transform 1 0 26680 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_286
timestamp 1644511149
transform 1 0 27416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_297
timestamp 1644511149
transform 1 0 28428 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_304
timestamp 1644511149
transform 1 0 29072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_331
timestamp 1644511149
transform 1 0 31556 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_354
timestamp 1644511149
transform 1 0 33672 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1644511149
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_370
timestamp 1644511149
transform 1 0 35144 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_381
timestamp 1644511149
transform 1 0 36156 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_385
timestamp 1644511149
transform 1 0 36524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_392
timestamp 1644511149
transform 1 0 37168 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_399
timestamp 1644511149
transform 1 0 37812 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_10
timestamp 1644511149
transform 1 0 2024 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_19
timestamp 1644511149
transform 1 0 2852 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_24
timestamp 1644511149
transform 1 0 3312 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_31
timestamp 1644511149
transform 1 0 3956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_42
timestamp 1644511149
transform 1 0 4968 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_46
timestamp 1644511149
transform 1 0 5336 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1644511149
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_64
timestamp 1644511149
transform 1 0 6992 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_72
timestamp 1644511149
transform 1 0 7728 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_80
timestamp 1644511149
transform 1 0 8464 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_86
timestamp 1644511149
transform 1 0 9016 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_99
timestamp 1644511149
transform 1 0 10212 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_106
timestamp 1644511149
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_119
timestamp 1644511149
transform 1 0 12052 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_134
timestamp 1644511149
transform 1 0 13432 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_144
timestamp 1644511149
transform 1 0 14352 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1644511149
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_179
timestamp 1644511149
transform 1 0 17572 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_201
timestamp 1644511149
transform 1 0 19596 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_209
timestamp 1644511149
transform 1 0 20332 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1644511149
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_229
timestamp 1644511149
transform 1 0 22172 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_246
timestamp 1644511149
transform 1 0 23736 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_255
timestamp 1644511149
transform 1 0 24564 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1644511149
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_285
timestamp 1644511149
transform 1 0 27324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_302
timestamp 1644511149
transform 1 0 28888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_322
timestamp 1644511149
transform 1 0 30728 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_353
timestamp 1644511149
transform 1 0 33580 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_382
timestamp 1644511149
transform 1 0 36248 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_390
timestamp 1644511149
transform 1 0 36984 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_396
timestamp 1644511149
transform 1 0 37536 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_404
timestamp 1644511149
transform 1 0 38272 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_10
timestamp 1644511149
transform 1 0 2024 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_17
timestamp 1644511149
transform 1 0 2668 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1644511149
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_45
timestamp 1644511149
transform 1 0 5244 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_56
timestamp 1644511149
transform 1 0 6256 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_62
timestamp 1644511149
transform 1 0 6808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_73
timestamp 1644511149
transform 1 0 7820 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1644511149
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_92
timestamp 1644511149
transform 1 0 9568 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_116
timestamp 1644511149
transform 1 0 11776 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_124
timestamp 1644511149
transform 1 0 12512 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_157
timestamp 1644511149
transform 1 0 15548 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_168
timestamp 1644511149
transform 1 0 16560 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_172
timestamp 1644511149
transform 1 0 16928 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_200
timestamp 1644511149
transform 1 0 19504 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_241
timestamp 1644511149
transform 1 0 23276 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1644511149
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_260
timestamp 1644511149
transform 1 0 25024 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_267
timestamp 1644511149
transform 1 0 25668 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_274
timestamp 1644511149
transform 1 0 26312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_281
timestamp 1644511149
transform 1 0 26956 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_294
timestamp 1644511149
transform 1 0 28152 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_303
timestamp 1644511149
transform 1 0 28980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_327
timestamp 1644511149
transform 1 0 31188 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_334
timestamp 1644511149
transform 1 0 31832 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_341
timestamp 1644511149
transform 1 0 32476 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_352
timestamp 1644511149
transform 1 0 33488 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_359
timestamp 1644511149
transform 1 0 34132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_370
timestamp 1644511149
transform 1 0 35144 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_374
timestamp 1644511149
transform 1 0 35512 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_378
timestamp 1644511149
transform 1 0 35880 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_385 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 36524 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_397
timestamp 1644511149
transform 1 0 37628 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_405
timestamp 1644511149
transform 1 0 38364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_6
timestamp 1644511149
transform 1 0 1656 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_12
timestamp 1644511149
transform 1 0 2208 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_16
timestamp 1644511149
transform 1 0 2576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_23
timestamp 1644511149
transform 1 0 3220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_43
timestamp 1644511149
transform 1 0 5060 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_50
timestamp 1644511149
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_73
timestamp 1644511149
transform 1 0 7820 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_107
timestamp 1644511149
transform 1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_133
timestamp 1644511149
transform 1 0 13340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_141
timestamp 1644511149
transform 1 0 14076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_152
timestamp 1644511149
transform 1 0 15088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1644511149
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_182
timestamp 1644511149
transform 1 0 17848 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_189
timestamp 1644511149
transform 1 0 18492 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_207
timestamp 1644511149
transform 1 0 20148 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1644511149
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_232
timestamp 1644511149
transform 1 0 22448 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_239
timestamp 1644511149
transform 1 0 23092 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_246
timestamp 1644511149
transform 1 0 23736 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_257
timestamp 1644511149
transform 1 0 24748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_264
timestamp 1644511149
transform 1 0 25392 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_271
timestamp 1644511149
transform 1 0 26036 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_297
timestamp 1644511149
transform 1 0 28428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_315
timestamp 1644511149
transform 1 0 30084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_324
timestamp 1644511149
transform 1 0 30912 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_331
timestamp 1644511149
transform 1 0 31556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_341
timestamp 1644511149
transform 1 0 32476 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_351
timestamp 1644511149
transform 1 0 33396 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_371
timestamp 1644511149
transform 1 0 35236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_378
timestamp 1644511149
transform 1 0 35880 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_14
timestamp 1644511149
transform 1 0 2392 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_18
timestamp 1644511149
transform 1 0 2760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1644511149
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_33
timestamp 1644511149
transform 1 0 4140 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_39
timestamp 1644511149
transform 1 0 4692 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_48
timestamp 1644511149
transform 1 0 5520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_55
timestamp 1644511149
transform 1 0 6164 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_61
timestamp 1644511149
transform 1 0 6716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_79
timestamp 1644511149
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_92
timestamp 1644511149
transform 1 0 9568 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_103
timestamp 1644511149
transform 1 0 10580 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_114
timestamp 1644511149
transform 1 0 11592 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_125
timestamp 1644511149
transform 1 0 12604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1644511149
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_155
timestamp 1644511149
transform 1 0 15364 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_164
timestamp 1644511149
transform 1 0 16192 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_172
timestamp 1644511149
transform 1 0 16928 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_180
timestamp 1644511149
transform 1 0 17664 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_188
timestamp 1644511149
transform 1 0 18400 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_204
timestamp 1644511149
transform 1 0 19872 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_211
timestamp 1644511149
transform 1 0 20516 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_218
timestamp 1644511149
transform 1 0 21160 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_232
timestamp 1644511149
transform 1 0 22448 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_241
timestamp 1644511149
transform 1 0 23276 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_248
timestamp 1644511149
transform 1 0 23920 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_256
timestamp 1644511149
transform 1 0 24656 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_272
timestamp 1644511149
transform 1 0 26128 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_278
timestamp 1644511149
transform 1 0 26680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_297
timestamp 1644511149
transform 1 0 28428 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1644511149
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_312
timestamp 1644511149
transform 1 0 29808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_319
timestamp 1644511149
transform 1 0 30452 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_326
timestamp 1644511149
transform 1 0 31096 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_355
timestamp 1644511149
transform 1 0 33764 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_371
timestamp 1644511149
transform 1 0 35236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_381
timestamp 1644511149
transform 1 0 36156 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_393
timestamp 1644511149
transform 1 0 37260 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_405
timestamp 1644511149
transform 1 0 38364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_6
timestamp 1644511149
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_18
timestamp 1644511149
transform 1 0 2760 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_26
timestamp 1644511149
transform 1 0 3496 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_31
timestamp 1644511149
transform 1 0 3956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_38
timestamp 1644511149
transform 1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_45
timestamp 1644511149
transform 1 0 5244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1644511149
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_61
timestamp 1644511149
transform 1 0 6716 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_71
timestamp 1644511149
transform 1 0 7636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_75
timestamp 1644511149
transform 1 0 8004 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_79
timestamp 1644511149
transform 1 0 8372 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_92
timestamp 1644511149
transform 1 0 9568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_101
timestamp 1644511149
transform 1 0 10396 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1644511149
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_118
timestamp 1644511149
transform 1 0 11960 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_131
timestamp 1644511149
transform 1 0 13156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_140
timestamp 1644511149
transform 1 0 13984 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_152
timestamp 1644511149
transform 1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_156
timestamp 1644511149
transform 1 0 15456 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_162
timestamp 1644511149
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_178
timestamp 1644511149
transform 1 0 17480 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_198
timestamp 1644511149
transform 1 0 19320 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_209
timestamp 1644511149
transform 1 0 20332 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_216
timestamp 1644511149
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_241
timestamp 1644511149
transform 1 0 23276 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_247
timestamp 1644511149
transform 1 0 23828 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_255
timestamp 1644511149
transform 1 0 24564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1644511149
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_301
timestamp 1644511149
transform 1 0 28796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_308
timestamp 1644511149
transform 1 0 29440 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_315
timestamp 1644511149
transform 1 0 30084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_322
timestamp 1644511149
transform 1 0 30728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_342
timestamp 1644511149
transform 1 0 32568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_353
timestamp 1644511149
transform 1 0 33580 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_370
timestamp 1644511149
transform 1 0 35144 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_382
timestamp 1644511149
transform 1 0 36248 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_390
timestamp 1644511149
transform 1 0 36984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1644511149
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_38
timestamp 1644511149
transform 1 0 4600 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_42
timestamp 1644511149
transform 1 0 4968 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_64
timestamp 1644511149
transform 1 0 6992 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_68
timestamp 1644511149
transform 1 0 7360 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_76
timestamp 1644511149
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_95
timestamp 1644511149
transform 1 0 9844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_99
timestamp 1644511149
transform 1 0 10212 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_116
timestamp 1644511149
transform 1 0 11776 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1644511149
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_145
timestamp 1644511149
transform 1 0 14444 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_149
timestamp 1644511149
transform 1 0 14812 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_156
timestamp 1644511149
transform 1 0 15456 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_164
timestamp 1644511149
transform 1 0 16192 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_172
timestamp 1644511149
transform 1 0 16928 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1644511149
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_219
timestamp 1644511149
transform 1 0 21252 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_227
timestamp 1644511149
transform 1 0 21988 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_244
timestamp 1644511149
transform 1 0 23552 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_269
timestamp 1644511149
transform 1 0 25852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_280
timestamp 1644511149
transform 1 0 26864 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_288
timestamp 1644511149
transform 1 0 27600 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_300
timestamp 1644511149
transform 1 0 28704 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_314
timestamp 1644511149
transform 1 0 29992 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_328
timestamp 1644511149
transform 1 0 31280 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_335
timestamp 1644511149
transform 1 0 31924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_347
timestamp 1644511149
transform 1 0 33028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_359
timestamp 1644511149
transform 1 0 34132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_46
timestamp 1644511149
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1644511149
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_73
timestamp 1644511149
transform 1 0 7820 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_99
timestamp 1644511149
transform 1 0 10212 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1644511149
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_121
timestamp 1644511149
transform 1 0 12236 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_129
timestamp 1644511149
transform 1 0 12972 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_144
timestamp 1644511149
transform 1 0 14352 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_152
timestamp 1644511149
transform 1 0 15088 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1644511149
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_175
timestamp 1644511149
transform 1 0 17204 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_186
timestamp 1644511149
transform 1 0 18216 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_190
timestamp 1644511149
transform 1 0 18584 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_198
timestamp 1644511149
transform 1 0 19320 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_213
timestamp 1644511149
transform 1 0 20700 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1644511149
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_229
timestamp 1644511149
transform 1 0 22172 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_245
timestamp 1644511149
transform 1 0 23644 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_254
timestamp 1644511149
transform 1 0 24472 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_258
timestamp 1644511149
transform 1 0 24840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_266
timestamp 1644511149
transform 1 0 25576 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_284
timestamp 1644511149
transform 1 0 27232 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_300
timestamp 1644511149
transform 1 0 28704 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_307
timestamp 1644511149
transform 1 0 29348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_314
timestamp 1644511149
transform 1 0 29992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_321
timestamp 1644511149
transform 1 0 30636 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_328
timestamp 1644511149
transform 1 0 31280 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_47
timestamp 1644511149
transform 1 0 5428 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_58
timestamp 1644511149
transform 1 0 6440 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_64
timestamp 1644511149
transform 1 0 6992 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_72
timestamp 1644511149
transform 1 0 7728 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1644511149
transform 1 0 8372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_95
timestamp 1644511149
transform 1 0 9844 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_119
timestamp 1644511149
transform 1 0 12052 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_128
timestamp 1644511149
transform 1 0 12880 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1644511149
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_152
timestamp 1644511149
transform 1 0 15088 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_176
timestamp 1644511149
transform 1 0 17296 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1644511149
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_200
timestamp 1644511149
transform 1 0 19504 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1644511149
transform 1 0 20700 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_219
timestamp 1644511149
transform 1 0 21252 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_230
timestamp 1644511149
transform 1 0 22264 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_237
timestamp 1644511149
transform 1 0 22908 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_264
timestamp 1644511149
transform 1 0 25392 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_284
timestamp 1644511149
transform 1 0 27232 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1644511149
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_312
timestamp 1644511149
transform 1 0 29808 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_319
timestamp 1644511149
transform 1 0 30452 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_328
timestamp 1644511149
transform 1 0 31280 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_340
timestamp 1644511149
transform 1 0 32384 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_352
timestamp 1644511149
transform 1 0 33488 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_42
timestamp 1644511149
transform 1 0 4968 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_46
timestamp 1644511149
transform 1 0 5336 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1644511149
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_61
timestamp 1644511149
transform 1 0 6716 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_72
timestamp 1644511149
transform 1 0 7728 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_76
timestamp 1644511149
transform 1 0 8096 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_80
timestamp 1644511149
transform 1 0 8464 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_100
timestamp 1644511149
transform 1 0 10304 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1644511149
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_117
timestamp 1644511149
transform 1 0 11868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_122
timestamp 1644511149
transform 1 0 12328 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_130
timestamp 1644511149
transform 1 0 13064 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_147
timestamp 1644511149
transform 1 0 14628 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_155
timestamp 1644511149
transform 1 0 15364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_177
timestamp 1644511149
transform 1 0 17388 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_185
timestamp 1644511149
transform 1 0 18124 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_192
timestamp 1644511149
transform 1 0 18768 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_200
timestamp 1644511149
transform 1 0 19504 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_243
timestamp 1644511149
transform 1 0 23460 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_254
timestamp 1644511149
transform 1 0 24472 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_265
timestamp 1644511149
transform 1 0 25484 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_271
timestamp 1644511149
transform 1 0 26036 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1644511149
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_289
timestamp 1644511149
transform 1 0 27692 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_296
timestamp 1644511149
transform 1 0 28336 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_303
timestamp 1644511149
transform 1 0 28980 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_310
timestamp 1644511149
transform 1 0 29624 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_324
timestamp 1644511149
transform 1 0 30912 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_37
timestamp 1644511149
transform 1 0 4508 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_52
timestamp 1644511149
transform 1 0 5888 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_60
timestamp 1644511149
transform 1 0 6624 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_67
timestamp 1644511149
transform 1 0 7268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_76
timestamp 1644511149
transform 1 0 8096 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_90
timestamp 1644511149
transform 1 0 9384 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_98
timestamp 1644511149
transform 1 0 10120 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_102
timestamp 1644511149
transform 1 0 10488 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_110
timestamp 1644511149
transform 1 0 11224 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_120
timestamp 1644511149
transform 1 0 12144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_131
timestamp 1644511149
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_144
timestamp 1644511149
transform 1 0 14352 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_152
timestamp 1644511149
transform 1 0 15088 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_164
timestamp 1644511149
transform 1 0 16192 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_173
timestamp 1644511149
transform 1 0 17020 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_182
timestamp 1644511149
transform 1 0 17848 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_190
timestamp 1644511149
transform 1 0 18584 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_201
timestamp 1644511149
transform 1 0 19596 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_205
timestamp 1644511149
transform 1 0 19964 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_214
timestamp 1644511149
transform 1 0 20792 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_234
timestamp 1644511149
transform 1 0 22632 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1644511149
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_269
timestamp 1644511149
transform 1 0 25852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_283
timestamp 1644511149
transform 1 0 27140 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_291
timestamp 1644511149
transform 1 0 27876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_298
timestamp 1644511149
transform 1 0 28520 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1644511149
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_312
timestamp 1644511149
transform 1 0 29808 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_324
timestamp 1644511149
transform 1 0 30912 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_336
timestamp 1644511149
transform 1 0 32016 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_348
timestamp 1644511149
transform 1 0 33120 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_360
timestamp 1644511149
transform 1 0 34224 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_73
timestamp 1644511149
transform 1 0 7820 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_77
timestamp 1644511149
transform 1 0 8188 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_95
timestamp 1644511149
transform 1 0 9844 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_103
timestamp 1644511149
transform 1 0 10580 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1644511149
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_116
timestamp 1644511149
transform 1 0 11776 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_124
timestamp 1644511149
transform 1 0 12512 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_133
timestamp 1644511149
transform 1 0 13340 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_145
timestamp 1644511149
transform 1 0 14444 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_157
timestamp 1644511149
transform 1 0 15548 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1644511149
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_175
timestamp 1644511149
transform 1 0 17204 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_198
timestamp 1644511149
transform 1 0 19320 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_211
timestamp 1644511149
transform 1 0 20516 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1644511149
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_242
timestamp 1644511149
transform 1 0 23368 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_258
timestamp 1644511149
transform 1 0 24840 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_266
timestamp 1644511149
transform 1 0 25576 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_270
timestamp 1644511149
transform 1 0 25944 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_276
timestamp 1644511149
transform 1 0 26496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_297
timestamp 1644511149
transform 1 0 28428 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_304
timestamp 1644511149
transform 1 0 29072 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_316
timestamp 1644511149
transform 1 0 30176 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_328
timestamp 1644511149
transform 1 0 31280 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_69
timestamp 1644511149
transform 1 0 7452 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_73
timestamp 1644511149
transform 1 0 7820 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1644511149
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_90
timestamp 1644511149
transform 1 0 9384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_117
timestamp 1644511149
transform 1 0 11868 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_125
timestamp 1644511149
transform 1 0 12604 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_131
timestamp 1644511149
transform 1 0 13156 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1644511149
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_150
timestamp 1644511149
transform 1 0 14904 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_161
timestamp 1644511149
transform 1 0 15916 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_169
timestamp 1644511149
transform 1 0 16652 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_181
timestamp 1644511149
transform 1 0 17756 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_187
timestamp 1644511149
transform 1 0 18308 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1644511149
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_213
timestamp 1644511149
transform 1 0 20700 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_222
timestamp 1644511149
transform 1 0 21528 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_228
timestamp 1644511149
transform 1 0 22080 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_236
timestamp 1644511149
transform 1 0 22816 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1644511149
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_258
timestamp 1644511149
transform 1 0 24840 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_267
timestamp 1644511149
transform 1 0 25668 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_274
timestamp 1644511149
transform 1 0 26312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_288
timestamp 1644511149
transform 1 0 27600 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_299
timestamp 1644511149
transform 1 0 28612 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_76
timestamp 1644511149
transform 1 0 8096 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_96
timestamp 1644511149
transform 1 0 9936 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_118
timestamp 1644511149
transform 1 0 11960 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_126
timestamp 1644511149
transform 1 0 12696 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_132
timestamp 1644511149
transform 1 0 13248 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_150
timestamp 1644511149
transform 1 0 14904 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_158
timestamp 1644511149
transform 1 0 15640 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1644511149
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_179
timestamp 1644511149
transform 1 0 17572 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_195
timestamp 1644511149
transform 1 0 19044 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_203
timestamp 1644511149
transform 1 0 19780 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1644511149
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_229
timestamp 1644511149
transform 1 0 22172 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_235
timestamp 1644511149
transform 1 0 22724 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_244
timestamp 1644511149
transform 1 0 23552 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_253
timestamp 1644511149
transform 1 0 24380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_271
timestamp 1644511149
transform 1 0 26036 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_297
timestamp 1644511149
transform 1 0 28428 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_304
timestamp 1644511149
transform 1 0 29072 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_316
timestamp 1644511149
transform 1 0 30176 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_328
timestamp 1644511149
transform 1 0 31280 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1644511149
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_94
timestamp 1644511149
transform 1 0 9752 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_100
timestamp 1644511149
transform 1 0 10304 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_117
timestamp 1644511149
transform 1 0 11868 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_126
timestamp 1644511149
transform 1 0 12696 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1644511149
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_147
timestamp 1644511149
transform 1 0 14628 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_158
timestamp 1644511149
transform 1 0 15640 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_167
timestamp 1644511149
transform 1 0 16468 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_176
timestamp 1644511149
transform 1 0 17296 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_182
timestamp 1644511149
transform 1 0 17848 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_188
timestamp 1644511149
transform 1 0 18400 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_202
timestamp 1644511149
transform 1 0 19688 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1644511149
transform 1 0 20424 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_220
timestamp 1644511149
transform 1 0 21344 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_224
timestamp 1644511149
transform 1 0 21712 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_239
timestamp 1644511149
transform 1 0 23092 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1644511149
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_257
timestamp 1644511149
transform 1 0 24748 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_274
timestamp 1644511149
transform 1 0 26312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_282
timestamp 1644511149
transform 1 0 27048 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_290
timestamp 1644511149
transform 1 0 27784 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_297
timestamp 1644511149
transform 1 0 28428 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_305
timestamp 1644511149
transform 1 0 29164 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_89
timestamp 1644511149
transform 1 0 9292 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_97
timestamp 1644511149
transform 1 0 10028 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_102
timestamp 1644511149
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1644511149
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_118
timestamp 1644511149
transform 1 0 11960 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_124
timestamp 1644511149
transform 1 0 12512 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_128
timestamp 1644511149
transform 1 0 12880 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_136
timestamp 1644511149
transform 1 0 13616 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_142
timestamp 1644511149
transform 1 0 14168 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1644511149
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1644511149
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_174
timestamp 1644511149
transform 1 0 17112 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_183
timestamp 1644511149
transform 1 0 17940 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_190
timestamp 1644511149
transform 1 0 18584 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_201
timestamp 1644511149
transform 1 0 19596 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_210
timestamp 1644511149
transform 1 0 20424 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_219
timestamp 1644511149
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_241
timestamp 1644511149
transform 1 0 23276 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_265
timestamp 1644511149
transform 1 0 25484 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_274
timestamp 1644511149
transform 1 0 26312 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_284
timestamp 1644511149
transform 1 0 27232 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_296
timestamp 1644511149
transform 1 0 28336 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_308
timestamp 1644511149
transform 1 0 29440 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_320
timestamp 1644511149
transform 1 0 30544 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1644511149
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_69
timestamp 1644511149
transform 1 0 7452 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_73
timestamp 1644511149
transform 1 0 7820 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1644511149
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_90
timestamp 1644511149
transform 1 0 9384 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_117
timestamp 1644511149
transform 1 0 11868 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_123
timestamp 1644511149
transform 1 0 12420 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_127
timestamp 1644511149
transform 1 0 12788 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1644511149
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_157
timestamp 1644511149
transform 1 0 15548 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_164
timestamp 1644511149
transform 1 0 16192 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_176
timestamp 1644511149
transform 1 0 17296 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_185
timestamp 1644511149
transform 1 0 18124 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1644511149
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_213
timestamp 1644511149
transform 1 0 20700 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_228
timestamp 1644511149
transform 1 0 22080 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_237
timestamp 1644511149
transform 1 0 22908 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_257
timestamp 1644511149
transform 1 0 24748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_264
timestamp 1644511149
transform 1 0 25392 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_276
timestamp 1644511149
transform 1 0 26496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_294
timestamp 1644511149
transform 1 0 28152 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_306
timestamp 1644511149
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_65
timestamp 1644511149
transform 1 0 7084 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_89
timestamp 1644511149
transform 1 0 9292 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_98
timestamp 1644511149
transform 1 0 10120 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_104
timestamp 1644511149
transform 1 0 10672 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1644511149
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_118
timestamp 1644511149
transform 1 0 11960 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_142
timestamp 1644511149
transform 1 0 14168 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_163
timestamp 1644511149
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_173
timestamp 1644511149
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_182
timestamp 1644511149
transform 1 0 17848 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_186
timestamp 1644511149
transform 1 0 18216 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_195
timestamp 1644511149
transform 1 0 19044 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_199
timestamp 1644511149
transform 1 0 19412 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_210
timestamp 1644511149
transform 1 0 20424 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_235
timestamp 1644511149
transform 1 0 22724 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_244
timestamp 1644511149
transform 1 0 23552 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_251
timestamp 1644511149
transform 1 0 24196 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_271
timestamp 1644511149
transform 1 0 26036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_297
timestamp 1644511149
transform 1 0 28428 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_309
timestamp 1644511149
transform 1 0 29532 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_321
timestamp 1644511149
transform 1 0 30636 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_333
timestamp 1644511149
transform 1 0 31740 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_61
timestamp 1644511149
transform 1 0 6716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1644511149
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_90
timestamp 1644511149
transform 1 0 9384 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_98
timestamp 1644511149
transform 1 0 10120 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_116
timestamp 1644511149
transform 1 0 11776 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_122
timestamp 1644511149
transform 1 0 12328 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_128
timestamp 1644511149
transform 1 0 12880 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 1644511149
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_152
timestamp 1644511149
transform 1 0 15088 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_172
timestamp 1644511149
transform 1 0 16928 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_181
timestamp 1644511149
transform 1 0 17756 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_202
timestamp 1644511149
transform 1 0 19688 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_222
timestamp 1644511149
transform 1 0 21528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_229
timestamp 1644511149
transform 1 0 22172 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_239
timestamp 1644511149
transform 1 0 23092 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_246
timestamp 1644511149
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_262
timestamp 1644511149
transform 1 0 25208 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_270
timestamp 1644511149
transform 1 0 25944 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_282
timestamp 1644511149
transform 1 0 27048 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_292
timestamp 1644511149
transform 1 0 27968 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_302
timestamp 1644511149
transform 1 0 28888 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_65
timestamp 1644511149
transform 1 0 7084 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_89
timestamp 1644511149
transform 1 0 9292 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_98
timestamp 1644511149
transform 1 0 10120 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_104
timestamp 1644511149
transform 1 0 10672 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1644511149
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_129
timestamp 1644511149
transform 1 0 12972 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_143
timestamp 1644511149
transform 1 0 14260 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_155
timestamp 1644511149
transform 1 0 15364 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_162
timestamp 1644511149
transform 1 0 16008 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_172
timestamp 1644511149
transform 1 0 16928 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_190
timestamp 1644511149
transform 1 0 18584 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_194
timestamp 1644511149
transform 1 0 18952 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_201
timestamp 1644511149
transform 1 0 19596 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_215
timestamp 1644511149
transform 1 0 20884 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_247
timestamp 1644511149
transform 1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_275
timestamp 1644511149
transform 1 0 26404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_290
timestamp 1644511149
transform 1 0 27784 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_300
timestamp 1644511149
transform 1 0 28704 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_312
timestamp 1644511149
transform 1 0 29808 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_324
timestamp 1644511149
transform 1 0 30912 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1644511149
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_90
timestamp 1644511149
transform 1 0 9384 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_102
timestamp 1644511149
transform 1 0 10488 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_119
timestamp 1644511149
transform 1 0 12052 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_126
timestamp 1644511149
transform 1 0 12696 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_132
timestamp 1644511149
transform 1 0 13248 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1644511149
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_144
timestamp 1644511149
transform 1 0 14352 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_154
timestamp 1644511149
transform 1 0 15272 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_164
timestamp 1644511149
transform 1 0 16192 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_172
timestamp 1644511149
transform 1 0 16928 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1644511149
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_239
timestamp 1644511149
transform 1 0 23092 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_246
timestamp 1644511149
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_257
timestamp 1644511149
transform 1 0 24748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_268
timestamp 1644511149
transform 1 0 25760 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_281
timestamp 1644511149
transform 1 0 26956 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_287
timestamp 1644511149
transform 1 0 27508 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1644511149
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_89
timestamp 1644511149
transform 1 0 9292 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_97
timestamp 1644511149
transform 1 0 10028 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_103
timestamp 1644511149
transform 1 0 10580 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_120
timestamp 1644511149
transform 1 0 12144 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_127
timestamp 1644511149
transform 1 0 12788 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_141
timestamp 1644511149
transform 1 0 14076 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_155
timestamp 1644511149
transform 1 0 15364 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1644511149
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_183
timestamp 1644511149
transform 1 0 17940 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_191
timestamp 1644511149
transform 1 0 18676 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_203
timestamp 1644511149
transform 1 0 19780 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_216
timestamp 1644511149
transform 1 0 20976 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_235
timestamp 1644511149
transform 1 0 22724 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_244
timestamp 1644511149
transform 1 0 23552 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_264
timestamp 1644511149
transform 1 0 25392 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_274
timestamp 1644511149
transform 1 0 26312 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_290
timestamp 1644511149
transform 1 0 27784 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_300
timestamp 1644511149
transform 1 0 28704 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_312
timestamp 1644511149
transform 1 0 29808 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_324
timestamp 1644511149
transform 1 0 30912 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_101
timestamp 1644511149
transform 1 0 10396 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_110
timestamp 1644511149
transform 1 0 11224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_118
timestamp 1644511149
transform 1 0 11960 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_126
timestamp 1644511149
transform 1 0 12696 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1644511149
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_157
timestamp 1644511149
transform 1 0 15548 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_169
timestamp 1644511149
transform 1 0 16652 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_179
timestamp 1644511149
transform 1 0 17572 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1644511149
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_206
timestamp 1644511149
transform 1 0 20056 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_210
timestamp 1644511149
transform 1 0 20424 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_231
timestamp 1644511149
transform 1 0 22356 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_262
timestamp 1644511149
transform 1 0 25208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_266
timestamp 1644511149
transform 1 0 25576 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_276
timestamp 1644511149
transform 1 0 26496 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_284
timestamp 1644511149
transform 1 0 27232 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_302
timestamp 1644511149
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1644511149
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_98
timestamp 1644511149
transform 1 0 10120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_106
timestamp 1644511149
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_117
timestamp 1644511149
transform 1 0 11868 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_135
timestamp 1644511149
transform 1 0 13524 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_147
timestamp 1644511149
transform 1 0 14628 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1644511149
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_191
timestamp 1644511149
transform 1 0 18676 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_219
timestamp 1644511149
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_235
timestamp 1644511149
transform 1 0 22724 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_248
timestamp 1644511149
transform 1 0 23920 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_261
timestamp 1644511149
transform 1 0 25116 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1644511149
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_297
timestamp 1644511149
transform 1 0 28428 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_307
timestamp 1644511149
transform 1 0 29348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_319
timestamp 1644511149
transform 1 0 30452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_331
timestamp 1644511149
transform 1 0 31556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_111
timestamp 1644511149
transform 1 0 11316 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_122
timestamp 1644511149
transform 1 0 12328 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_126
timestamp 1644511149
transform 1 0 12696 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_135
timestamp 1644511149
transform 1 0 13524 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_151
timestamp 1644511149
transform 1 0 14996 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_164
timestamp 1644511149
transform 1 0 16192 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_176
timestamp 1644511149
transform 1 0 17296 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_188
timestamp 1644511149
transform 1 0 18400 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_229
timestamp 1644511149
transform 1 0 22172 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1644511149
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_271
timestamp 1644511149
transform 1 0 26036 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_279
timestamp 1644511149
transform 1 0 26772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_299
timestamp 1644511149
transform 1 0 28612 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_87
timestamp 1644511149
transform 1 0 9108 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_95
timestamp 1644511149
transform 1 0 9844 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1644511149
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_120
timestamp 1644511149
transform 1 0 12144 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_128
timestamp 1644511149
transform 1 0 12880 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_132
timestamp 1644511149
transform 1 0 13248 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_145
timestamp 1644511149
transform 1 0 14444 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_153
timestamp 1644511149
transform 1 0 15180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1644511149
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_175
timestamp 1644511149
transform 1 0 17204 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_189
timestamp 1644511149
transform 1 0 18492 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_195
timestamp 1644511149
transform 1 0 19044 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_206
timestamp 1644511149
transform 1 0 20056 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_210
timestamp 1644511149
transform 1 0 20424 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1644511149
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_235
timestamp 1644511149
transform 1 0 22724 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_243
timestamp 1644511149
transform 1 0 23460 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_255
timestamp 1644511149
transform 1 0 24564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_275
timestamp 1644511149
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_287
timestamp 1644511149
transform 1 0 27508 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_304
timestamp 1644511149
transform 1 0 29072 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_316
timestamp 1644511149
transform 1 0 30176 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_328
timestamp 1644511149
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_361
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1644511149
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_92
timestamp 1644511149
transform 1 0 9568 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_100
timestamp 1644511149
transform 1 0 10304 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_113
timestamp 1644511149
transform 1 0 11500 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_123
timestamp 1644511149
transform 1 0 12420 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_132
timestamp 1644511149
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_144
timestamp 1644511149
transform 1 0 14352 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_156
timestamp 1644511149
transform 1 0 15456 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_173
timestamp 1644511149
transform 1 0 17020 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_179
timestamp 1644511149
transform 1 0 17572 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1644511149
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_206
timestamp 1644511149
transform 1 0 20056 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_216
timestamp 1644511149
transform 1 0 20976 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_238
timestamp 1644511149
transform 1 0 23000 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1644511149
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_273
timestamp 1644511149
transform 1 0 26220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_281
timestamp 1644511149
transform 1 0 26956 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_285
timestamp 1644511149
transform 1 0 27324 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_302
timestamp 1644511149
transform 1 0 28888 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_333
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_345
timestamp 1644511149
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1644511149
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_76
timestamp 1644511149
transform 1 0 8096 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_96
timestamp 1644511149
transform 1 0 9936 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_102
timestamp 1644511149
transform 1 0 10488 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_107
timestamp 1644511149
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_124
timestamp 1644511149
transform 1 0 12512 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_132
timestamp 1644511149
transform 1 0 13248 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_140
timestamp 1644511149
transform 1 0 13984 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_158
timestamp 1644511149
transform 1 0 15640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1644511149
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_173
timestamp 1644511149
transform 1 0 17020 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_182
timestamp 1644511149
transform 1 0 17848 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_186
timestamp 1644511149
transform 1 0 18216 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_213
timestamp 1644511149
transform 1 0 20700 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_221
timestamp 1644511149
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_241
timestamp 1644511149
transform 1 0 23276 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_289
timestamp 1644511149
transform 1 0 27692 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_297
timestamp 1644511149
transform 1 0 28428 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_309
timestamp 1644511149
transform 1 0 29532 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_321
timestamp 1644511149
transform 1 0 30636 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_333
timestamp 1644511149
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_71
timestamp 1644511149
transform 1 0 7636 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1644511149
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_98
timestamp 1644511149
transform 1 0 10120 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_112
timestamp 1644511149
transform 1 0 11408 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_120
timestamp 1644511149
transform 1 0 12144 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_129
timestamp 1644511149
transform 1 0 12972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1644511149
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1644511149
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_162
timestamp 1644511149
transform 1 0 16008 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_170
timestamp 1644511149
transform 1 0 16744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_187
timestamp 1644511149
transform 1 0 18308 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_203
timestamp 1644511149
transform 1 0 19780 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_223
timestamp 1644511149
transform 1 0 21620 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_235
timestamp 1644511149
transform 1 0 22724 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_239
timestamp 1644511149
transform 1 0 23092 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_248
timestamp 1644511149
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_263
timestamp 1644511149
transform 1 0 25300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_283
timestamp 1644511149
transform 1 0 27140 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_296
timestamp 1644511149
transform 1 0 28336 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1644511149
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1644511149
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1644511149
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_121
timestamp 1644511149
transform 1 0 12236 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_144
timestamp 1644511149
transform 1 0 14352 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_155
timestamp 1644511149
transform 1 0 15364 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_159
timestamp 1644511149
transform 1 0 15732 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1644511149
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_177
timestamp 1644511149
transform 1 0 17388 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_184
timestamp 1644511149
transform 1 0 18032 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_192
timestamp 1644511149
transform 1 0 18768 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_211
timestamp 1644511149
transform 1 0 20516 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_215
timestamp 1644511149
transform 1 0 20884 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1644511149
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_233
timestamp 1644511149
transform 1 0 22540 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_244
timestamp 1644511149
transform 1 0 23552 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_253
timestamp 1644511149
transform 1 0 24380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_261
timestamp 1644511149
transform 1 0 25116 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_269
timestamp 1644511149
transform 1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1644511149
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_290
timestamp 1644511149
transform 1 0 27784 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_297
timestamp 1644511149
transform 1 0 28428 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_317
timestamp 1644511149
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1644511149
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_73
timestamp 1644511149
transform 1 0 7820 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1644511149
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_94
timestamp 1644511149
transform 1 0 9752 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_110
timestamp 1644511149
transform 1 0 11224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_117
timestamp 1644511149
transform 1 0 11868 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_128
timestamp 1644511149
transform 1 0 12880 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1644511149
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_144
timestamp 1644511149
transform 1 0 14352 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_157
timestamp 1644511149
transform 1 0 15548 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_171
timestamp 1644511149
transform 1 0 16836 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_191
timestamp 1644511149
transform 1 0 18676 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_215
timestamp 1644511149
transform 1 0 20884 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_223
timestamp 1644511149
transform 1 0 21620 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_235
timestamp 1644511149
transform 1 0 22724 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_246
timestamp 1644511149
transform 1 0 23736 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_263
timestamp 1644511149
transform 1 0 25300 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_271
timestamp 1644511149
transform 1 0 26036 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_283
timestamp 1644511149
transform 1 0 27140 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_294
timestamp 1644511149
transform 1 0 28152 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_303
timestamp 1644511149
transform 1 0 28980 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_314
timestamp 1644511149
transform 1 0 29992 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_326
timestamp 1644511149
transform 1 0 31096 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_338
timestamp 1644511149
transform 1 0 32200 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_350
timestamp 1644511149
transform 1 0 33304 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1644511149
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_66
timestamp 1644511149
transform 1 0 7176 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_73
timestamp 1644511149
transform 1 0 7820 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_83
timestamp 1644511149
transform 1 0 8740 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_91
timestamp 1644511149
transform 1 0 9476 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_100
timestamp 1644511149
transform 1 0 10304 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1644511149
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_117
timestamp 1644511149
transform 1 0 11868 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_130
timestamp 1644511149
transform 1 0 13064 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_134
timestamp 1644511149
transform 1 0 13432 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_140
timestamp 1644511149
transform 1 0 13984 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_151
timestamp 1644511149
transform 1 0 14996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_159
timestamp 1644511149
transform 1 0 15732 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_173
timestamp 1644511149
transform 1 0 17020 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_183
timestamp 1644511149
transform 1 0 17940 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_192
timestamp 1644511149
transform 1 0 18768 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_202
timestamp 1644511149
transform 1 0 19688 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_216
timestamp 1644511149
transform 1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_234
timestamp 1644511149
transform 1 0 22632 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_249
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_253
timestamp 1644511149
transform 1 0 24380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_270
timestamp 1644511149
transform 1 0 25944 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1644511149
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_294
timestamp 1644511149
transform 1 0 28152 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_314
timestamp 1644511149
transform 1 0 29992 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_326
timestamp 1644511149
transform 1 0 31096 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1644511149
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_73
timestamp 1644511149
transform 1 0 7820 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1644511149
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_93
timestamp 1644511149
transform 1 0 9660 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_101
timestamp 1644511149
transform 1 0 10396 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_119
timestamp 1644511149
transform 1 0 12052 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_144
timestamp 1644511149
transform 1 0 14352 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_156
timestamp 1644511149
transform 1 0 15456 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_162
timestamp 1644511149
transform 1 0 16008 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_179
timestamp 1644511149
transform 1 0 17572 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_188
timestamp 1644511149
transform 1 0 18400 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_228
timestamp 1644511149
transform 1 0 22080 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_241
timestamp 1644511149
transform 1 0 23276 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1644511149
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_260
timestamp 1644511149
transform 1 0 25024 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_267
timestamp 1644511149
transform 1 0 25668 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_275
timestamp 1644511149
transform 1 0 26404 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_286
timestamp 1644511149
transform 1 0 27416 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_294
timestamp 1644511149
transform 1 0 28152 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_300
timestamp 1644511149
transform 1 0 28704 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_325
timestamp 1644511149
transform 1 0 31004 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_337
timestamp 1644511149
transform 1 0 32108 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_349
timestamp 1644511149
transform 1 0 33212 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_361
timestamp 1644511149
transform 1 0 34316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_65
timestamp 1644511149
transform 1 0 7084 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_83
timestamp 1644511149
transform 1 0 8740 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_91
timestamp 1644511149
transform 1 0 9476 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_97
timestamp 1644511149
transform 1 0 10028 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1644511149
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_116
timestamp 1644511149
transform 1 0 11776 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_128
timestamp 1644511149
transform 1 0 12880 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_138
timestamp 1644511149
transform 1 0 13800 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_145
timestamp 1644511149
transform 1 0 14444 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_156
timestamp 1644511149
transform 1 0 15456 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1644511149
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_178
timestamp 1644511149
transform 1 0 17480 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_202
timestamp 1644511149
transform 1 0 19688 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_214
timestamp 1644511149
transform 1 0 20792 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1644511149
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_234
timestamp 1644511149
transform 1 0 22632 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_258
timestamp 1644511149
transform 1 0 24840 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_266
timestamp 1644511149
transform 1 0 25576 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_290
timestamp 1644511149
transform 1 0 27784 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_299
timestamp 1644511149
transform 1 0 28612 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_306
timestamp 1644511149
transform 1 0 29256 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_313
timestamp 1644511149
transform 1 0 29900 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_325
timestamp 1644511149
transform 1 0 31004 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_333
timestamp 1644511149
transform 1 0 31740 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_94
timestamp 1644511149
transform 1 0 9752 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_107
timestamp 1644511149
transform 1 0 10948 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_117
timestamp 1644511149
transform 1 0 11868 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_124
timestamp 1644511149
transform 1 0 12512 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_135
timestamp 1644511149
transform 1 0 13524 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_145
timestamp 1644511149
transform 1 0 14444 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_155
timestamp 1644511149
transform 1 0 15364 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_166
timestamp 1644511149
transform 1 0 16376 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_174
timestamp 1644511149
transform 1 0 17112 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_188
timestamp 1644511149
transform 1 0 18400 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_205
timestamp 1644511149
transform 1 0 19964 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_213
timestamp 1644511149
transform 1 0 20700 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_224
timestamp 1644511149
transform 1 0 21712 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_235
timestamp 1644511149
transform 1 0 22724 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1644511149
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_272
timestamp 1644511149
transform 1 0 26128 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_285
timestamp 1644511149
transform 1 0 27324 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_293
timestamp 1644511149
transform 1 0 28060 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_300
timestamp 1644511149
transform 1 0 28704 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1644511149
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_78
timestamp 1644511149
transform 1 0 8280 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_82
timestamp 1644511149
transform 1 0 8648 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_92
timestamp 1644511149
transform 1 0 9568 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_118
timestamp 1644511149
transform 1 0 11960 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_126
timestamp 1644511149
transform 1 0 12696 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_136
timestamp 1644511149
transform 1 0 13616 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_145
timestamp 1644511149
transform 1 0 14444 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_153
timestamp 1644511149
transform 1 0 15180 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_174
timestamp 1644511149
transform 1 0 17112 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_182
timestamp 1644511149
transform 1 0 17848 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_187
timestamp 1644511149
transform 1 0 18308 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_204
timestamp 1644511149
transform 1 0 19872 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_212
timestamp 1644511149
transform 1 0 20608 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1644511149
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_274
timestamp 1644511149
transform 1 0 26312 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_303
timestamp 1644511149
transform 1 0 28980 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_315
timestamp 1644511149
transform 1 0 30084 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_327
timestamp 1644511149
transform 1 0 31188 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_61
timestamp 1644511149
transform 1 0 6716 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_80
timestamp 1644511149
transform 1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_93
timestamp 1644511149
transform 1 0 9660 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_100
timestamp 1644511149
transform 1 0 10304 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_110
timestamp 1644511149
transform 1 0 11224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_114
timestamp 1644511149
transform 1 0 11592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_120
timestamp 1644511149
transform 1 0 12144 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_130
timestamp 1644511149
transform 1 0 13064 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1644511149
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_148
timestamp 1644511149
transform 1 0 14720 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_160
timestamp 1644511149
transform 1 0 15824 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_166
timestamp 1644511149
transform 1 0 16376 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_171
timestamp 1644511149
transform 1 0 16836 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_180
timestamp 1644511149
transform 1 0 17664 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1644511149
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_202
timestamp 1644511149
transform 1 0 19688 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_214
timestamp 1644511149
transform 1 0 20792 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_225
timestamp 1644511149
transform 1 0 21804 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_231
timestamp 1644511149
transform 1 0 22356 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_240
timestamp 1644511149
transform 1 0 23184 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_244
timestamp 1644511149
transform 1 0 23552 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_258
timestamp 1644511149
transform 1 0 24840 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_266
timestamp 1644511149
transform 1 0 25576 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_273
timestamp 1644511149
transform 1 0 26220 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_279
timestamp 1644511149
transform 1 0 26772 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_283
timestamp 1644511149
transform 1 0 27140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_295
timestamp 1644511149
transform 1 0 28244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1644511149
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_68
timestamp 1644511149
transform 1 0 7360 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_87
timestamp 1644511149
transform 1 0 9108 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_97
timestamp 1644511149
transform 1 0 10028 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_103
timestamp 1644511149
transform 1 0 10580 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1644511149
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_117
timestamp 1644511149
transform 1 0 11868 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_122
timestamp 1644511149
transform 1 0 12328 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_133
timestamp 1644511149
transform 1 0 13340 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_157
timestamp 1644511149
transform 1 0 15548 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1644511149
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_178
timestamp 1644511149
transform 1 0 17480 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_185
timestamp 1644511149
transform 1 0 18124 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_198
timestamp 1644511149
transform 1 0 19320 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_202
timestamp 1644511149
transform 1 0 19688 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_206
timestamp 1644511149
transform 1 0 20056 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1644511149
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_232
timestamp 1644511149
transform 1 0 22448 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_239
timestamp 1644511149
transform 1 0 23092 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_246
timestamp 1644511149
transform 1 0 23736 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_253
timestamp 1644511149
transform 1 0 24380 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_261
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_267
timestamp 1644511149
transform 1 0 25668 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_274
timestamp 1644511149
transform 1 0 26312 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_299
timestamp 1644511149
transform 1 0 28612 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_311
timestamp 1644511149
transform 1 0 29716 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_323
timestamp 1644511149
transform 1 0 30820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_73
timestamp 1644511149
transform 1 0 7820 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1644511149
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_91
timestamp 1644511149
transform 1 0 9476 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_95
timestamp 1644511149
transform 1 0 9844 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_105
timestamp 1644511149
transform 1 0 10764 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_115
timestamp 1644511149
transform 1 0 11684 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_127
timestamp 1644511149
transform 1 0 12788 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_135
timestamp 1644511149
transform 1 0 13524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_145
timestamp 1644511149
transform 1 0 14444 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_157
timestamp 1644511149
transform 1 0 15548 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_169
timestamp 1644511149
transform 1 0 16652 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_179
timestamp 1644511149
transform 1 0 17572 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_188
timestamp 1644511149
transform 1 0 18400 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_200
timestamp 1644511149
transform 1 0 19504 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_206
timestamp 1644511149
transform 1 0 20056 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_210
timestamp 1644511149
transform 1 0 20424 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_219
timestamp 1644511149
transform 1 0 21252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_230
timestamp 1644511149
transform 1 0 22264 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_237
timestamp 1644511149
transform 1 0 22908 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_244
timestamp 1644511149
transform 1 0 23552 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_258
timestamp 1644511149
transform 1 0 24840 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_264
timestamp 1644511149
transform 1 0 25392 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_274
timestamp 1644511149
transform 1 0 26312 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_296
timestamp 1644511149
transform 1 0 28336 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_76
timestamp 1644511149
transform 1 0 8096 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_88
timestamp 1644511149
transform 1 0 9200 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_96
timestamp 1644511149
transform 1 0 9936 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1644511149
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_116
timestamp 1644511149
transform 1 0 11776 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_130
timestamp 1644511149
transform 1 0 13064 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_142
timestamp 1644511149
transform 1 0 14168 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_146
timestamp 1644511149
transform 1 0 14536 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_155
timestamp 1644511149
transform 1 0 15364 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1644511149
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_174
timestamp 1644511149
transform 1 0 17112 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_187
timestamp 1644511149
transform 1 0 18308 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_198
timestamp 1644511149
transform 1 0 19320 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_207
timestamp 1644511149
transform 1 0 20148 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_214
timestamp 1644511149
transform 1 0 20792 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1644511149
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_231
timestamp 1644511149
transform 1 0 22356 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_239
timestamp 1644511149
transform 1 0 23092 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_274
timestamp 1644511149
transform 1 0 26312 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_288
timestamp 1644511149
transform 1 0 27600 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_297
timestamp 1644511149
transform 1 0 28428 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_309
timestamp 1644511149
transform 1 0 29532 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_321
timestamp 1644511149
transform 1 0 30636 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_333
timestamp 1644511149
transform 1 0 31740 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_73
timestamp 1644511149
transform 1 0 7820 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1644511149
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_94
timestamp 1644511149
transform 1 0 9752 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_102
timestamp 1644511149
transform 1 0 10488 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_120
timestamp 1644511149
transform 1 0 12144 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1644511149
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_145
timestamp 1644511149
transform 1 0 14444 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_152
timestamp 1644511149
transform 1 0 15088 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_163
timestamp 1644511149
transform 1 0 16100 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_183
timestamp 1644511149
transform 1 0 17940 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1644511149
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_204
timestamp 1644511149
transform 1 0 19872 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_210
timestamp 1644511149
transform 1 0 20424 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_217
timestamp 1644511149
transform 1 0 21068 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_225
timestamp 1644511149
transform 1 0 21804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_242
timestamp 1644511149
transform 1 0 23368 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_250
timestamp 1644511149
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_260
timestamp 1644511149
transform 1 0 25024 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_266
timestamp 1644511149
transform 1 0 25576 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_274
timestamp 1644511149
transform 1 0 26312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_283
timestamp 1644511149
transform 1 0 27140 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_290
timestamp 1644511149
transform 1 0 27784 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_302
timestamp 1644511149
transform 1 0 28888 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1644511149
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_84
timestamp 1644511149
transform 1 0 8832 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_104
timestamp 1644511149
transform 1 0 10672 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_131
timestamp 1644511149
transform 1 0 13156 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_140
timestamp 1644511149
transform 1 0 13984 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_144
timestamp 1644511149
transform 1 0 14352 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_148
timestamp 1644511149
transform 1 0 14720 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_159
timestamp 1644511149
transform 1 0 15732 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_172
timestamp 1644511149
transform 1 0 16928 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_182
timestamp 1644511149
transform 1 0 17848 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_201
timestamp 1644511149
transform 1 0 19596 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_213
timestamp 1644511149
transform 1 0 20700 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1644511149
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_235
timestamp 1644511149
transform 1 0 22724 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_241
timestamp 1644511149
transform 1 0 23276 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_251
timestamp 1644511149
transform 1 0 24196 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_265
timestamp 1644511149
transform 1 0 25484 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1644511149
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_286
timestamp 1644511149
transform 1 0 27416 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_101
timestamp 1644511149
transform 1 0 10396 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_113
timestamp 1644511149
transform 1 0 11500 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_119
timestamp 1644511149
transform 1 0 12052 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1644511149
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_163
timestamp 1644511149
transform 1 0 16100 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_171
timestamp 1644511149
transform 1 0 16836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_183
timestamp 1644511149
transform 1 0 17940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_204
timestamp 1644511149
transform 1 0 19872 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_217
timestamp 1644511149
transform 1 0 21068 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_229
timestamp 1644511149
transform 1 0 22172 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_240
timestamp 1644511149
transform 1 0 23184 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_247
timestamp 1644511149
transform 1 0 23828 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_266
timestamp 1644511149
transform 1 0 25576 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_279
timestamp 1644511149
transform 1 0 26772 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_299
timestamp 1644511149
transform 1 0 28612 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_129
timestamp 1644511149
transform 1 0 12972 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_133
timestamp 1644511149
transform 1 0 13340 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_141
timestamp 1644511149
transform 1 0 14076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_159
timestamp 1644511149
transform 1 0 15732 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_173
timestamp 1644511149
transform 1 0 17020 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_185
timestamp 1644511149
transform 1 0 18124 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_189
timestamp 1644511149
transform 1 0 18492 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_199
timestamp 1644511149
transform 1 0 19412 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_203
timestamp 1644511149
transform 1 0 19780 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_207
timestamp 1644511149
transform 1 0 20148 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_215
timestamp 1644511149
transform 1 0 20884 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1644511149
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_230
timestamp 1644511149
transform 1 0 22264 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_239
timestamp 1644511149
transform 1 0 23092 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_248
timestamp 1644511149
transform 1 0 23920 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_262
timestamp 1644511149
transform 1 0 25208 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_275
timestamp 1644511149
transform 1 0 26404 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_288
timestamp 1644511149
transform 1 0 27600 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_300
timestamp 1644511149
transform 1 0 28704 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_312
timestamp 1644511149
transform 1 0 29808 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_324
timestamp 1644511149
transform 1 0 30912 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_147
timestamp 1644511149
transform 1 0 14628 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_151
timestamp 1644511149
transform 1 0 14996 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_159
timestamp 1644511149
transform 1 0 15732 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_182
timestamp 1644511149
transform 1 0 17848 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1644511149
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_206
timestamp 1644511149
transform 1 0 20056 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_210
timestamp 1644511149
transform 1 0 20424 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_220
timestamp 1644511149
transform 1 0 21344 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_229
timestamp 1644511149
transform 1 0 22172 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_238
timestamp 1644511149
transform 1 0 23000 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_273
timestamp 1644511149
transform 1 0 26220 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_291
timestamp 1644511149
transform 1 0 27876 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_298
timestamp 1644511149
transform 1 0 28520 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_306
timestamp 1644511149
transform 1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_157
timestamp 1644511149
transform 1 0 15548 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_164
timestamp 1644511149
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_185
timestamp 1644511149
transform 1 0 18124 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_199
timestamp 1644511149
transform 1 0 19412 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_212
timestamp 1644511149
transform 1 0 20608 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_228
timestamp 1644511149
transform 1 0 22080 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_245
timestamp 1644511149
transform 1 0 23644 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_252
timestamp 1644511149
transform 1 0 24288 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_258
timestamp 1644511149
transform 1 0 24840 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_266
timestamp 1644511149
transform 1 0 25576 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_275
timestamp 1644511149
transform 1 0 26404 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_286
timestamp 1644511149
transform 1 0 27416 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_298
timestamp 1644511149
transform 1 0 28520 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_310
timestamp 1644511149
transform 1 0 29624 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_322
timestamp 1644511149
transform 1 0 30728 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1644511149
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_169
timestamp 1644511149
transform 1 0 16652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_175
timestamp 1644511149
transform 1 0 17204 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_183
timestamp 1644511149
transform 1 0 17940 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1644511149
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_207
timestamp 1644511149
transform 1 0 20148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_229
timestamp 1644511149
transform 1 0 22172 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_237
timestamp 1644511149
transform 1 0 22908 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1644511149
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_256
timestamp 1644511149
transform 1 0 24656 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_276
timestamp 1644511149
transform 1 0 26496 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_288
timestamp 1644511149
transform 1 0 27600 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_300
timestamp 1644511149
transform 1 0 28704 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1644511149
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_172
timestamp 1644511149
transform 1 0 16928 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_180
timestamp 1644511149
transform 1 0 17664 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_190
timestamp 1644511149
transform 1 0 18584 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_203
timestamp 1644511149
transform 1 0 19780 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_207
timestamp 1644511149
transform 1 0 20148 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_234
timestamp 1644511149
transform 1 0 22632 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_247
timestamp 1644511149
transform 1 0 23828 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_258
timestamp 1644511149
transform 1 0 24840 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_267
timestamp 1644511149
transform 1 0 25668 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_274
timestamp 1644511149
transform 1 0 26312 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_173
timestamp 1644511149
transform 1 0 17020 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_181
timestamp 1644511149
transform 1 0 17756 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1644511149
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_204
timestamp 1644511149
transform 1 0 19872 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_212
timestamp 1644511149
transform 1 0 20608 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_222
timestamp 1644511149
transform 1 0 21528 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_235
timestamp 1644511149
transform 1 0 22724 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_246
timestamp 1644511149
transform 1 0 23736 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_269
timestamp 1644511149
transform 1 0 25852 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_281
timestamp 1644511149
transform 1 0 26956 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_293
timestamp 1644511149
transform 1 0 28060 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_305
timestamp 1644511149
transform 1 0 29164 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_188
timestamp 1644511149
transform 1 0 18400 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_55_203
timestamp 1644511149
transform 1 0 19780 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_211
timestamp 1644511149
transform 1 0 20516 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1644511149
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_235
timestamp 1644511149
transform 1 0 22724 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_241
timestamp 1644511149
transform 1 0 23276 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_258
timestamp 1644511149
transform 1 0 24840 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_265
timestamp 1644511149
transform 1 0 25484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_277
timestamp 1644511149
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_174
timestamp 1644511149
transform 1 0 17112 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_183
timestamp 1644511149
transform 1 0 17940 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1644511149
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_213
timestamp 1644511149
transform 1 0 20700 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_242
timestamp 1644511149
transform 1 0 23368 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1644511149
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_258
timestamp 1644511149
transform 1 0 24840 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_270
timestamp 1644511149
transform 1 0 25944 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_282
timestamp 1644511149
transform 1 0 27048 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_294
timestamp 1644511149
transform 1 0 28152 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_306
timestamp 1644511149
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_177
timestamp 1644511149
transform 1 0 17388 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_183
timestamp 1644511149
transform 1 0 17940 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_203
timestamp 1644511149
transform 1 0 19780 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_207
timestamp 1644511149
transform 1 0 20148 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_211
timestamp 1644511149
transform 1 0 20516 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1644511149
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_247
timestamp 1644511149
transform 1 0 23828 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_254
timestamp 1644511149
transform 1 0 24472 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_266
timestamp 1644511149
transform 1 0 25576 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1644511149
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_200
timestamp 1644511149
transform 1 0 19504 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_208
timestamp 1644511149
transform 1 0 20240 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_227
timestamp 1644511149
transform 1 0 21988 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_231
timestamp 1644511149
transform 1 0 22356 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_237
timestamp 1644511149
transform 1 0 22908 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_244
timestamp 1644511149
transform 1 0 23552 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1644511149
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_228
timestamp 1644511149
transform 1 0 22080 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_240
timestamp 1644511149
transform 1 0 23184 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_252
timestamp 1644511149
transform 1 0 24288 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_264
timestamp 1644511149
transform 1 0 25392 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_276
timestamp 1644511149
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1644511149
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1644511149
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1644511149
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1644511149
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_317
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_277
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_289
timestamp 1644511149
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1644511149
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_345
timestamp 1644511149
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1644511149
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1644511149
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_193
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_205
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1644511149
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1644511149
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_249
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_261
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1644511149
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1644511149
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_317
timestamp 1644511149
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1644511149
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1644511149
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_209
timestamp 1644511149
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_221
timestamp 1644511149
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1644511149
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1644511149
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_265
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_277
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_289
timestamp 1644511149
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1644511149
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1644511149
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1644511149
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1644511149
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_15
timestamp 1644511149
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_27
timestamp 1644511149
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_181
timestamp 1644511149
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_237
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_249
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_261
timestamp 1644511149
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1644511149
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_317
timestamp 1644511149
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1644511149
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_177
timestamp 1644511149
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1644511149
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1644511149
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_209
timestamp 1644511149
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_233
timestamp 1644511149
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1644511149
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_265
timestamp 1644511149
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_277
timestamp 1644511149
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_289
timestamp 1644511149
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1644511149
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1644511149
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_333
timestamp 1644511149
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_345
timestamp 1644511149
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1644511149
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1644511149
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_193
timestamp 1644511149
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_237
timestamp 1644511149
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_249
timestamp 1644511149
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_261
timestamp 1644511149
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_293
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_305
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1644511149
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_209
timestamp 1644511149
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1644511149
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_265
timestamp 1644511149
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_277
timestamp 1644511149
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_289
timestamp 1644511149
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1644511149
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1644511149
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1644511149
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1644511149
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1644511149
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_193
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_237
timestamp 1644511149
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_249
timestamp 1644511149
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_261
timestamp 1644511149
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1644511149
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1644511149
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1644511149
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1644511149
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_233
timestamp 1644511149
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1644511149
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1644511149
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_27
timestamp 1644511149
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1644511149
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1644511149
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_237
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1644511149
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_27
timestamp 1644511149
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_39
timestamp 1644511149
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1644511149
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_289
timestamp 1644511149
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1644511149
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1644511149
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1644511149
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1644511149
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1644511149
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_39
timestamp 1644511149
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1644511149
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1644511149
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1644511149
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1644511149
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1644511149
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1644511149
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_349
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_361
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_373
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1644511149
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1644511149
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_15
timestamp 1644511149
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1644511149
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1644511149
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1644511149
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1644511149
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_109
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_121
timestamp 1644511149
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1644511149
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1644511149
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_141
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_153
timestamp 1644511149
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_165
timestamp 1644511149
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_177
timestamp 1644511149
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1644511149
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1644511149
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_209
timestamp 1644511149
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_221
timestamp 1644511149
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_233
timestamp 1644511149
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1644511149
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1644511149
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_265
timestamp 1644511149
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_277
timestamp 1644511149
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_289
timestamp 1644511149
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1644511149
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_333
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_345
timestamp 1644511149
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1644511149
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1644511149
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_15
timestamp 1644511149
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1644511149
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_39
timestamp 1644511149
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1644511149
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1644511149
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1644511149
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_121
timestamp 1644511149
transform 1 0 12236 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_126
timestamp 1644511149
transform 1 0 12696 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_138
timestamp 1644511149
transform 1 0 13800 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_150
timestamp 1644511149
transform 1 0 14904 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_158
timestamp 1644511149
transform 1 0 15640 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_164
timestamp 1644511149
transform 1 0 16192 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_205
timestamp 1644511149
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1644511149
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1644511149
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_237
timestamp 1644511149
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_249
timestamp 1644511149
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_261
timestamp 1644511149
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1644511149
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1644511149
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_305
timestamp 1644511149
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_317
timestamp 1644511149
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1644511149
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_337
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_349
timestamp 1644511149
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_361
timestamp 1644511149
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_373
timestamp 1644511149
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1644511149
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1644511149
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_405
timestamp 1644511149
transform 1 0 38364 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_3
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_15
timestamp 1644511149
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1644511149
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_29
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_39
timestamp 1644511149
transform 1 0 4692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_51
timestamp 1644511149
transform 1 0 5796 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_55
timestamp 1644511149
transform 1 0 6164 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_57
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_69
timestamp 1644511149
transform 1 0 7452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_81
timestamp 1644511149
transform 1 0 8556 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_97
timestamp 1644511149
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_109
timestamp 1644511149
transform 1 0 11132 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_82_113
timestamp 1644511149
transform 1 0 11500 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_82_123
timestamp 1644511149
transform 1 0 12420 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_135
timestamp 1644511149
transform 1 0 13524 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1644511149
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_153
timestamp 1644511149
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_165
timestamp 1644511149
transform 1 0 16284 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_169
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_181
timestamp 1644511149
transform 1 0 17756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_193
timestamp 1644511149
transform 1 0 18860 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_205
timestamp 1644511149
transform 1 0 19964 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_210
timestamp 1644511149
transform 1 0 20424 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_222
timestamp 1644511149
transform 1 0 21528 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_225
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_237
timestamp 1644511149
transform 1 0 22908 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_249
timestamp 1644511149
transform 1 0 24012 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_265
timestamp 1644511149
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_277
timestamp 1644511149
transform 1 0 26588 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_281
timestamp 1644511149
transform 1 0 26956 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_297
timestamp 1644511149
transform 1 0 28428 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_305
timestamp 1644511149
transform 1 0 29164 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_321
timestamp 1644511149
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_333
timestamp 1644511149
transform 1 0 31740 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_337
timestamp 1644511149
transform 1 0 32108 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_349
timestamp 1644511149
transform 1 0 33212 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_361
timestamp 1644511149
transform 1 0 34316 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_82_386
timestamp 1644511149
transform 1 0 36616 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_82_393
timestamp 1644511149
transform 1 0 37260 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_405
timestamp 1644511149
transform 1 0 38364 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 38824 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 38824 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 38824 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 38824 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 38824 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 38824 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 38824 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 38824 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 38824 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 38824 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 38824 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 38824 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 38824 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 38824 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 38824 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 38824 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 38824 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 38824 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0826_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15916 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_2  _0827_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5060 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nand3_1  _0828_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12144 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0829_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7084 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0830_
timestamp 1644511149
transform 1 0 7360 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0831_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0832_
timestamp 1644511149
transform 1 0 13800 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0833_
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0834_
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0835_
timestamp 1644511149
transform 1 0 11684 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0836_
timestamp 1644511149
transform 1 0 12696 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _0837_
timestamp 1644511149
transform 1 0 13800 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0838_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0839_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14996 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0840_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15272 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _0841_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1644511149
transform 1 0 18216 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0843_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17480 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0844_
timestamp 1644511149
transform 1 0 17940 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0846_
timestamp 1644511149
transform 1 0 10396 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0847_
timestamp 1644511149
transform 1 0 10488 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0848_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10948 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0849_
timestamp 1644511149
transform 1 0 10580 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0850_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0851_
timestamp 1644511149
transform 1 0 10304 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _0852_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10212 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0853_
timestamp 1644511149
transform 1 0 11592 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0854_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_2  _0855_
timestamp 1644511149
transform 1 0 10672 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0856_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10120 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0857_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10304 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _0858_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11316 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _0859_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9200 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_1  _0860_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9568 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0861_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0862_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0863_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12788 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0864_
timestamp 1644511149
transform 1 0 12696 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__a22oi_1  _0865_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13248 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0866_
timestamp 1644511149
transform 1 0 11684 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _0867_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11868 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0868_
timestamp 1644511149
transform 1 0 9200 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o2bb2a_1  _0869_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10488 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0870_
timestamp 1644511149
transform 1 0 10488 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o2bb2a_1  _0871_
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0872_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12144 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0873_
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0874_
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a2111oi_1  _0875_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11776 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0876_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0877_
timestamp 1644511149
transform 1 0 11316 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0878_
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0879_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10396 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0880_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11592 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _0881_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12236 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_2  _0882_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12420 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__nand4_1  _0883_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13524 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0884_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14352 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0885_
timestamp 1644511149
transform 1 0 16744 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0886_
timestamp 1644511149
transform 1 0 16744 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _0887_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14720 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0888_
timestamp 1644511149
transform 1 0 15824 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0889_
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0890_
timestamp 1644511149
transform 1 0 14812 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0891_
timestamp 1644511149
transform 1 0 15916 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _0892_
timestamp 1644511149
transform 1 0 17940 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _0893_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16468 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _0894_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0895_
timestamp 1644511149
transform 1 0 16744 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0896_
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0897_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18676 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0898_
timestamp 1644511149
transform 1 0 19780 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0899_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18676 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _0900_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0901_
timestamp 1644511149
transform 1 0 27692 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0902_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22448 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0903_
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0904_
timestamp 1644511149
transform 1 0 18676 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0905_
timestamp 1644511149
transform 1 0 20884 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0906_
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0907_
timestamp 1644511149
transform 1 0 18308 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0908_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0909_
timestamp 1644511149
transform 1 0 20424 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0910_
timestamp 1644511149
transform 1 0 23092 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0911_
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0912_
timestamp 1644511149
transform 1 0 19228 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0913_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0914_
timestamp 1644511149
transform 1 0 19596 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0915_
timestamp 1644511149
transform 1 0 21252 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0916_
timestamp 1644511149
transform 1 0 22080 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0917_
timestamp 1644511149
transform 1 0 22172 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0918_
timestamp 1644511149
transform 1 0 16836 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0920_
timestamp 1644511149
transform 1 0 17480 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0921_
timestamp 1644511149
transform 1 0 18584 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0922_
timestamp 1644511149
transform 1 0 22724 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0923_
timestamp 1644511149
transform 1 0 21160 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0924_
timestamp 1644511149
transform 1 0 26496 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0925_
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0926_
timestamp 1644511149
transform 1 0 25484 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0927_
timestamp 1644511149
transform 1 0 25668 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0928_
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0929_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25760 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0930_
timestamp 1644511149
transform 1 0 22448 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0931_
timestamp 1644511149
transform 1 0 19688 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0932_
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _0933_
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_2  _0934_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20056 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0935_
timestamp 1644511149
transform 1 0 12420 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1644511149
transform 1 0 15732 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _0937_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14996 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _0938_
timestamp 1644511149
transform 1 0 15548 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0939_
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0940_
timestamp 1644511149
transform 1 0 12880 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _0941_
timestamp 1644511149
transform 1 0 12512 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0942_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _0943_
timestamp 1644511149
transform 1 0 15272 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0944_
timestamp 1644511149
transform 1 0 15272 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0945_
timestamp 1644511149
transform 1 0 18492 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0946_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15456 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0947_
timestamp 1644511149
transform 1 0 17020 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0948_
timestamp 1644511149
transform 1 0 32568 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0949_
timestamp 1644511149
transform 1 0 25300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0950_
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0951_
timestamp 1644511149
transform 1 0 13984 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0952_
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0953_
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0954_
timestamp 1644511149
transform 1 0 18308 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0955_
timestamp 1644511149
transform 1 0 16560 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0956_
timestamp 1644511149
transform 1 0 17020 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0957_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17112 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0958_
timestamp 1644511149
transform 1 0 18952 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0959_
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0960_
timestamp 1644511149
transform 1 0 16652 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0961_
timestamp 1644511149
transform 1 0 18400 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0962_
timestamp 1644511149
transform 1 0 20792 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0963_
timestamp 1644511149
transform 1 0 16836 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1644511149
transform 1 0 14076 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _0965_
timestamp 1644511149
transform 1 0 16560 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0966_
timestamp 1644511149
transform 1 0 20056 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0967_
timestamp 1644511149
transform 1 0 19504 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0968_
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0969_
timestamp 1644511149
transform 1 0 18216 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0970_
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0971_
timestamp 1644511149
transform 1 0 23552 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0972_
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0973_
timestamp 1644511149
transform 1 0 17940 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0974_
timestamp 1644511149
transform 1 0 20608 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0975_
timestamp 1644511149
transform 1 0 20240 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0976_
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0977_
timestamp 1644511149
transform 1 0 26680 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0978_
timestamp 1644511149
transform 1 0 17664 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0979_
timestamp 1644511149
transform 1 0 21804 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0980_
timestamp 1644511149
transform 1 0 21620 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0981_
timestamp 1644511149
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0982_
timestamp 1644511149
transform 1 0 16836 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0983_
timestamp 1644511149
transform 1 0 20056 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0984_
timestamp 1644511149
transform 1 0 20332 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0985_
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0986_
timestamp 1644511149
transform 1 0 26128 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0987_
timestamp 1644511149
transform 1 0 17480 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0988_
timestamp 1644511149
transform 1 0 23184 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0989_
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 1644511149
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0991_
timestamp 1644511149
transform 1 0 22448 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0992_
timestamp 1644511149
transform 1 0 18308 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0993_
timestamp 1644511149
transform 1 0 22264 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0994_
timestamp 1644511149
transform 1 0 22816 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0995_
timestamp 1644511149
transform 1 0 27692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0996_
timestamp 1644511149
transform 1 0 22264 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0997_
timestamp 1644511149
transform 1 0 18308 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0998_
timestamp 1644511149
transform 1 0 22172 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0999_
timestamp 1644511149
transform 1 0 22356 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1644511149
transform 1 0 22816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1001_
timestamp 1644511149
transform 1 0 27324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1002_
timestamp 1644511149
transform 1 0 25208 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_2  _1003_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26772 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1005_
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1644511149
transform 1 0 27600 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1007_
timestamp 1644511149
transform 1 0 24104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1008_
timestamp 1644511149
transform 1 0 24840 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1009_
timestamp 1644511149
transform 1 0 24104 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_2  _1011_
timestamp 1644511149
transform 1 0 27784 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _1012_
timestamp 1644511149
transform 1 0 25300 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1013_
timestamp 1644511149
transform 1 0 25392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1014_
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1015_
timestamp 1644511149
transform 1 0 25300 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1016_
timestamp 1644511149
transform 1 0 24472 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_2  _1018_
timestamp 1644511149
transform 1 0 27784 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1020_
timestamp 1644511149
transform 1 0 27324 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1644511149
transform 1 0 26036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1022_
timestamp 1644511149
transform 1 0 27968 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1023_
timestamp 1644511149
transform 1 0 25944 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1644511149
transform 1 0 26680 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1025_
timestamp 1644511149
transform 1 0 15732 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1026_
timestamp 1644511149
transform 1 0 23184 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1027_
timestamp 1644511149
transform 1 0 25392 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1028_
timestamp 1644511149
transform 1 0 29624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1029_
timestamp 1644511149
transform 1 0 17296 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1030_
timestamp 1644511149
transform 1 0 25576 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1031_
timestamp 1644511149
transform 1 0 26220 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 1644511149
transform 1 0 30360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1644511149
transform 1 0 31280 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1034_
timestamp 1644511149
transform 1 0 28428 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1644511149
transform 1 0 27876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1036_
timestamp 1644511149
transform 1 0 28336 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1644511149
transform 1 0 31096 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1038_
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1644511149
transform 1 0 33672 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1040_
timestamp 1644511149
transform 1 0 29256 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1644511149
transform 1 0 33304 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1042_
timestamp 1644511149
transform 1 0 31280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1043_
timestamp 1644511149
transform 1 0 35512 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1044_
timestamp 1644511149
transform 1 0 31188 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1045_
timestamp 1644511149
transform 1 0 31556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1046_
timestamp 1644511149
transform 1 0 31556 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1047_
timestamp 1644511149
transform 1 0 32200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1048_
timestamp 1644511149
transform 1 0 32384 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1049_
timestamp 1644511149
transform 1 0 35236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1050_
timestamp 1644511149
transform 1 0 32016 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1051_
timestamp 1644511149
transform 1 0 36156 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1052_
timestamp 1644511149
transform 1 0 33212 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1053_
timestamp 1644511149
transform 1 0 35880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1054_
timestamp 1644511149
transform 1 0 36800 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1055_
timestamp 1644511149
transform 1 0 33212 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1056_
timestamp 1644511149
transform 1 0 33764 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1057_
timestamp 1644511149
transform 1 0 35512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1058_
timestamp 1644511149
transform 1 0 35328 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1059_
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1060_
timestamp 1644511149
transform 1 0 36524 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1061_
timestamp 1644511149
transform 1 0 36248 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1062_
timestamp 1644511149
transform 1 0 36156 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1063_
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1064_
timestamp 1644511149
transform 1 0 36248 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1065_
timestamp 1644511149
transform 1 0 37536 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1066_
timestamp 1644511149
transform 1 0 33856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1067_
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1068_
timestamp 1644511149
transform 1 0 35604 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1069_
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1070_
timestamp 1644511149
transform 1 0 36248 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1071_
timestamp 1644511149
transform 1 0 18124 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1072_
timestamp 1644511149
transform 1 0 19320 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1073_
timestamp 1644511149
transform 1 0 14720 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1074_
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1075_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1076_
timestamp 1644511149
transform 1 0 13340 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1077_
timestamp 1644511149
transform 1 0 12420 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1078_
timestamp 1644511149
transform 1 0 12420 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1079_
timestamp 1644511149
transform 1 0 12880 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1080_
timestamp 1644511149
transform 1 0 12512 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1081_
timestamp 1644511149
transform 1 0 10488 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1082_
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1083_
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1084_
timestamp 1644511149
transform 1 0 21068 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1085_
timestamp 1644511149
transform 1 0 19504 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1086_
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1087_
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1088_
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1089_
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1090_
timestamp 1644511149
transform 1 0 13248 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1091_
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1092_
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1093_
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1094_
timestamp 1644511149
transform 1 0 7176 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1095_
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1096_
timestamp 1644511149
transform 1 0 9752 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1097_
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1098_
timestamp 1644511149
transform 1 0 7176 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1099_
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1100_
timestamp 1644511149
transform 1 0 7544 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1101_
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1102_
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1103_
timestamp 1644511149
transform 1 0 9292 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1104_
timestamp 1644511149
transform 1 0 9108 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1105_
timestamp 1644511149
transform 1 0 29624 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1106_
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_2  _1107_
timestamp 1644511149
transform 1 0 1564 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1108_
timestamp 1644511149
transform 1 0 14904 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1109_
timestamp 1644511149
transform 1 0 14720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1110_
timestamp 1644511149
transform 1 0 19228 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1111_
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1112_
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1113_
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1114_
timestamp 1644511149
transform 1 0 17848 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1115_
timestamp 1644511149
transform 1 0 16008 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1116_
timestamp 1644511149
transform 1 0 16560 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1117_
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1118_
timestamp 1644511149
transform 1 0 17572 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1119_
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1120_
timestamp 1644511149
transform 1 0 14352 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1121_
timestamp 1644511149
transform 1 0 13156 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1122_
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1123_
timestamp 1644511149
transform 1 0 13892 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1124_
timestamp 1644511149
transform 1 0 19780 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1125_
timestamp 1644511149
transform 1 0 20240 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1126_
timestamp 1644511149
transform 1 0 16560 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1127_
timestamp 1644511149
transform 1 0 17296 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1128_
timestamp 1644511149
transform 1 0 16928 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _1129_
timestamp 1644511149
transform 1 0 15548 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1130_
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1131_
timestamp 1644511149
transform 1 0 16744 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1132_
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1133_
timestamp 1644511149
transform 1 0 14168 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1134_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16192 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1135_
timestamp 1644511149
transform 1 0 16928 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1136_
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1137_
timestamp 1644511149
transform 1 0 14168 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1138_
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1139_
timestamp 1644511149
transform 1 0 16928 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1140_
timestamp 1644511149
transform 1 0 17020 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1141_
timestamp 1644511149
transform 1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1142_
timestamp 1644511149
transform 1 0 17940 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1143_
timestamp 1644511149
transform 1 0 18216 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1144_
timestamp 1644511149
transform 1 0 12788 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1145_
timestamp 1644511149
transform 1 0 18124 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1146_
timestamp 1644511149
transform 1 0 18124 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1147_
timestamp 1644511149
transform 1 0 20700 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1148_
timestamp 1644511149
transform 1 0 19228 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1149_
timestamp 1644511149
transform 1 0 19504 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1150_
timestamp 1644511149
transform 1 0 23460 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1151_
timestamp 1644511149
transform 1 0 19320 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1152_
timestamp 1644511149
transform 1 0 19412 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1153_
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1154_
timestamp 1644511149
transform 1 0 20516 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1155_
timestamp 1644511149
transform 1 0 20884 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1156_
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1157_
timestamp 1644511149
transform 1 0 20424 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1158_
timestamp 1644511149
transform 1 0 20976 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1159_
timestamp 1644511149
transform 1 0 20884 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1160_
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1161_
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1162_
timestamp 1644511149
transform 1 0 21620 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1163_
timestamp 1644511149
transform 1 0 25760 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1164_
timestamp 1644511149
transform 1 0 22080 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1165_
timestamp 1644511149
transform 1 0 21988 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1166_
timestamp 1644511149
transform 1 0 21988 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1167_
timestamp 1644511149
transform 1 0 13064 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1168_
timestamp 1644511149
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1169_
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1170_
timestamp 1644511149
transform 1 0 13248 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1171_
timestamp 1644511149
transform 1 0 23920 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1172_
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1173_
timestamp 1644511149
transform 1 0 25944 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1174_
timestamp 1644511149
transform 1 0 7360 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1175_
timestamp 1644511149
transform 1 0 7820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1176_
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1177_
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1178_
timestamp 1644511149
transform 1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1179_
timestamp 1644511149
transform 1 0 24932 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1180_
timestamp 1644511149
transform 1 0 24932 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1181_
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1182_
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1183_
timestamp 1644511149
transform 1 0 24104 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1184_
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1185_
timestamp 1644511149
transform 1 0 26220 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1186_
timestamp 1644511149
transform 1 0 25024 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1187_
timestamp 1644511149
transform 1 0 29072 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1188_
timestamp 1644511149
transform 1 0 24104 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1189_
timestamp 1644511149
transform 1 0 23460 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1190_
timestamp 1644511149
transform 1 0 22632 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1191_
timestamp 1644511149
transform 1 0 14444 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1192_
timestamp 1644511149
transform 1 0 13892 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1193_
timestamp 1644511149
transform 1 0 10212 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1194_
timestamp 1644511149
transform 1 0 6900 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1195_
timestamp 1644511149
transform 1 0 4324 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1196_
timestamp 1644511149
transform 1 0 4140 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1197_
timestamp 1644511149
transform 1 0 3680 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1198_
timestamp 1644511149
transform 1 0 11592 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1199_
timestamp 1644511149
transform 1 0 12420 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1200_
timestamp 1644511149
transform 1 0 8188 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1201_
timestamp 1644511149
transform 1 0 5612 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1202_
timestamp 1644511149
transform 1 0 4232 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1203_
timestamp 1644511149
transform 1 0 5428 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1204_
timestamp 1644511149
transform 1 0 8096 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1205_
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1206_
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1207_
timestamp 1644511149
transform 1 0 7084 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1208_
timestamp 1644511149
transform 1 0 7636 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1209_
timestamp 1644511149
transform 1 0 9752 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1210_
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1211_
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1212_
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1213_
timestamp 1644511149
transform 1 0 4416 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1214_
timestamp 1644511149
transform 1 0 4324 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1215_
timestamp 1644511149
transform 1 0 5796 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1216_
timestamp 1644511149
transform 1 0 5428 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1217_
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1218_
timestamp 1644511149
transform 1 0 4784 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1219_
timestamp 1644511149
transform 1 0 3956 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1220_
timestamp 1644511149
transform 1 0 5428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1221_
timestamp 1644511149
transform 1 0 6348 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1222_
timestamp 1644511149
transform 1 0 5428 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1223_
timestamp 1644511149
transform 1 0 4600 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1224_
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1225_
timestamp 1644511149
transform 1 0 5428 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1226_
timestamp 1644511149
transform 1 0 5888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1227_
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1228_
timestamp 1644511149
transform 1 0 6808 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1229_
timestamp 1644511149
transform 1 0 8096 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1230_
timestamp 1644511149
transform 1 0 7452 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1231_
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1232_
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1233_
timestamp 1644511149
transform 1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1234_
timestamp 1644511149
transform 1 0 7452 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1235_
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1236_
timestamp 1644511149
transform 1 0 6440 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1237_
timestamp 1644511149
transform 1 0 7636 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1238_
timestamp 1644511149
transform 1 0 6164 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1239_
timestamp 1644511149
transform 1 0 5520 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1240_
timestamp 1644511149
transform 1 0 8648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1241_
timestamp 1644511149
transform 1 0 9108 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1242_
timestamp 1644511149
transform 1 0 8832 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1243_
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1244_
timestamp 1644511149
transform 1 0 8004 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1245_
timestamp 1644511149
transform 1 0 7360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1246_
timestamp 1644511149
transform 1 0 6440 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1247_
timestamp 1644511149
transform 1 0 10028 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1248_
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1249_
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1250_
timestamp 1644511149
transform 1 0 6808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1251_
timestamp 1644511149
transform 1 0 10396 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1252_
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1253_
timestamp 1644511149
transform 1 0 9752 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1254_
timestamp 1644511149
transform 1 0 9936 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1255_
timestamp 1644511149
transform 1 0 9108 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1256_
timestamp 1644511149
transform 1 0 5612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1257_
timestamp 1644511149
transform 1 0 10120 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1258_
timestamp 1644511149
transform 1 0 9936 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1259_
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1260_
timestamp 1644511149
transform 1 0 9568 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1261_
timestamp 1644511149
transform 1 0 9936 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1262_
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1263_
timestamp 1644511149
transform 1 0 10304 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1264_
timestamp 1644511149
transform 1 0 9476 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1265_
timestamp 1644511149
transform 1 0 11040 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1266_
timestamp 1644511149
transform 1 0 14444 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1267_
timestamp 1644511149
transform 1 0 10948 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1268_
timestamp 1644511149
transform 1 0 10580 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1269_
timestamp 1644511149
transform 1 0 7544 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1270_
timestamp 1644511149
transform 1 0 11408 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1271_
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1272_
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1273_
timestamp 1644511149
transform 1 0 11960 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1274_
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1275_
timestamp 1644511149
transform 1 0 10580 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1276_
timestamp 1644511149
transform 1 0 12696 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1277_
timestamp 1644511149
transform 1 0 14628 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1278_
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1279_
timestamp 1644511149
transform 1 0 13340 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1280_
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1281_
timestamp 1644511149
transform 1 0 11868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1282_
timestamp 1644511149
transform 1 0 12788 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1283_
timestamp 1644511149
transform 1 0 12696 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1284_
timestamp 1644511149
transform 1 0 5244 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1285_
timestamp 1644511149
transform 1 0 12972 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1286_
timestamp 1644511149
transform 1 0 12880 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1287_
timestamp 1644511149
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1288_
timestamp 1644511149
transform 1 0 12972 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1289_
timestamp 1644511149
transform 1 0 13524 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1290_
timestamp 1644511149
transform 1 0 7820 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1291_
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1292_
timestamp 1644511149
transform 1 0 13432 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1293_
timestamp 1644511149
transform 1 0 6716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1294_
timestamp 1644511149
transform 1 0 15916 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1295_
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1296_
timestamp 1644511149
transform 1 0 21160 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1297_
timestamp 1644511149
transform 1 0 15456 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1298_
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1299_
timestamp 1644511149
transform 1 0 4968 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1300_
timestamp 1644511149
transform 1 0 15456 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1301_
timestamp 1644511149
transform 1 0 15732 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1302_
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1303_
timestamp 1644511149
transform 1 0 15364 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1304_
timestamp 1644511149
transform 1 0 15640 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1305_
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1306_
timestamp 1644511149
transform 1 0 18676 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1307_
timestamp 1644511149
transform 1 0 18032 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1308_
timestamp 1644511149
transform 1 0 13156 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1309_
timestamp 1644511149
transform 1 0 14628 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1310_
timestamp 1644511149
transform 1 0 14444 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1311_
timestamp 1644511149
transform 1 0 15824 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1312_
timestamp 1644511149
transform 1 0 20056 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1313_
timestamp 1644511149
transform 1 0 19320 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1314_
timestamp 1644511149
transform 1 0 14720 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1315_
timestamp 1644511149
transform 1 0 9844 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1316_
timestamp 1644511149
transform 1 0 13524 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1317_
timestamp 1644511149
transform 1 0 10672 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1318_
timestamp 1644511149
transform 1 0 11684 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1319_
timestamp 1644511149
transform 1 0 12880 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1320_
timestamp 1644511149
transform 1 0 17204 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1321_
timestamp 1644511149
transform 1 0 17940 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _1322_
timestamp 1644511149
transform 1 0 16836 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1323_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13248 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1324_
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1325_
timestamp 1644511149
transform 1 0 11960 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1326_
timestamp 1644511149
transform 1 0 12512 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1327_
timestamp 1644511149
transform 1 0 12144 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1328_
timestamp 1644511149
transform 1 0 13156 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1329_
timestamp 1644511149
transform 1 0 12696 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1330_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12052 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1331_
timestamp 1644511149
transform 1 0 14812 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1332_
timestamp 1644511149
transform 1 0 13984 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _1333_
timestamp 1644511149
transform 1 0 12880 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1334_
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1335_
timestamp 1644511149
transform 1 0 10672 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1336_
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _1337_
timestamp 1644511149
transform 1 0 13432 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1338_
timestamp 1644511149
transform 1 0 13064 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1339_
timestamp 1644511149
transform 1 0 8096 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1340_
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1341_
timestamp 1644511149
transform 1 0 12972 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1342_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1343_
timestamp 1644511149
transform 1 0 14168 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1344_
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1345_
timestamp 1644511149
transform 1 0 9108 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1346_
timestamp 1644511149
transform 1 0 8924 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _1347_
timestamp 1644511149
transform 1 0 9936 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1348_
timestamp 1644511149
transform 1 0 10212 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1349_
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1350_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7728 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1351_
timestamp 1644511149
transform 1 0 14076 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1352_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7728 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1353_
timestamp 1644511149
transform 1 0 7544 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1354_
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1355_
timestamp 1644511149
transform 1 0 7176 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1356_
timestamp 1644511149
transform 1 0 6900 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1357_
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1358_
timestamp 1644511149
transform 1 0 8188 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1359_
timestamp 1644511149
transform 1 0 9476 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1360_
timestamp 1644511149
transform 1 0 8740 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1361_
timestamp 1644511149
transform 1 0 8004 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1362_
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1363_
timestamp 1644511149
transform 1 0 7728 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1364_
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1365_
timestamp 1644511149
transform 1 0 9200 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1366_
timestamp 1644511149
transform 1 0 8004 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1367_
timestamp 1644511149
transform 1 0 7728 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1368_
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1369_
timestamp 1644511149
transform 1 0 9568 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _1370_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8004 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1371_
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1372_
timestamp 1644511149
transform 1 0 9936 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1373_
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1374_
timestamp 1644511149
transform 1 0 8464 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1375_
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1376_
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1377_
timestamp 1644511149
transform 1 0 7084 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1378_
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1379_
timestamp 1644511149
transform 1 0 10304 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1380_
timestamp 1644511149
transform 1 0 10764 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _1381_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13248 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_2  _1382_
timestamp 1644511149
transform 1 0 14720 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _1383_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15640 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1384_
timestamp 1644511149
transform 1 0 15548 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1385_
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_2  _1386_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15916 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1387_
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _1388_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1389_
timestamp 1644511149
transform 1 0 19136 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1390_
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1391_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1392_
timestamp 1644511149
transform 1 0 17940 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1393_
timestamp 1644511149
transform 1 0 18308 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1394_
timestamp 1644511149
transform 1 0 20516 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1395_
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1396_
timestamp 1644511149
transform 1 0 20424 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1397_
timestamp 1644511149
transform 1 0 17940 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1398_
timestamp 1644511149
transform 1 0 19044 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1399_
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1400_
timestamp 1644511149
transform 1 0 20148 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1401_
timestamp 1644511149
transform 1 0 17020 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1402_
timestamp 1644511149
transform 1 0 24196 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1403_
timestamp 1644511149
transform 1 0 22724 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1404_
timestamp 1644511149
transform 1 0 23092 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1405_
timestamp 1644511149
transform 1 0 21804 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1406_
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1407_
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1408_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1409_
timestamp 1644511149
transform 1 0 21896 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1410_
timestamp 1644511149
transform 1 0 22172 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1411_
timestamp 1644511149
transform 1 0 20516 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1412_
timestamp 1644511149
transform 1 0 25760 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1413_
timestamp 1644511149
transform 1 0 24840 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1414_
timestamp 1644511149
transform 1 0 24288 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1415_
timestamp 1644511149
transform 1 0 28152 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1416_
timestamp 1644511149
transform 1 0 26128 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1417_
timestamp 1644511149
transform 1 0 25484 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1418_
timestamp 1644511149
transform 1 0 25668 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1419_
timestamp 1644511149
transform 1 0 28060 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1420_
timestamp 1644511149
transform 1 0 25668 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1421_
timestamp 1644511149
transform 1 0 28796 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1422_
timestamp 1644511149
transform 1 0 26128 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1423_
timestamp 1644511149
transform 1 0 28152 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1424_
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1425_
timestamp 1644511149
transform 1 0 27416 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1426_
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1427_
timestamp 1644511149
transform 1 0 28336 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1428_
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1429_
timestamp 1644511149
transform 1 0 24840 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1430_
timestamp 1644511149
transform 1 0 17848 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1431_
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1432_
timestamp 1644511149
transform 1 0 20792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1433_
timestamp 1644511149
transform 1 0 21804 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1434_
timestamp 1644511149
transform 1 0 26128 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1435_
timestamp 1644511149
transform 1 0 19872 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1436_
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1437_
timestamp 1644511149
transform 1 0 21068 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1438_
timestamp 1644511149
transform 1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1439_
timestamp 1644511149
transform 1 0 23920 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1440_
timestamp 1644511149
transform 1 0 23092 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1441_
timestamp 1644511149
transform 1 0 23276 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1442_
timestamp 1644511149
transform 1 0 19872 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1443_
timestamp 1644511149
transform 1 0 28704 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1444_
timestamp 1644511149
transform 1 0 23920 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1445_
timestamp 1644511149
transform 1 0 23920 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1446_
timestamp 1644511149
transform 1 0 4968 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1447_
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1448_
timestamp 1644511149
transform 1 0 22816 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1449_
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1450_
timestamp 1644511149
transform 1 0 22172 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1451_
timestamp 1644511149
transform 1 0 26036 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1452_
timestamp 1644511149
transform 1 0 28060 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1453_
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1454_
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1455_
timestamp 1644511149
transform 1 0 28244 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1456_
timestamp 1644511149
transform 1 0 29808 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1457_
timestamp 1644511149
transform 1 0 25208 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1458_
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1459_
timestamp 1644511149
transform 1 0 29348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1460_
timestamp 1644511149
transform 1 0 26680 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1461_
timestamp 1644511149
transform 1 0 28152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1462_
timestamp 1644511149
transform 1 0 20792 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1463_
timestamp 1644511149
transform 1 0 28796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1464_
timestamp 1644511149
transform 1 0 26036 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1465_
timestamp 1644511149
transform 1 0 28796 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1466_
timestamp 1644511149
transform 1 0 28520 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1467_
timestamp 1644511149
transform 1 0 30176 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1468_
timestamp 1644511149
transform 1 0 28796 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1469_
timestamp 1644511149
transform 1 0 27508 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1470_
timestamp 1644511149
transform 1 0 27600 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1471_
timestamp 1644511149
transform 1 0 28796 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1472_
timestamp 1644511149
transform 1 0 30820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1473_
timestamp 1644511149
transform 1 0 28520 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1474_
timestamp 1644511149
transform 1 0 30452 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1475_
timestamp 1644511149
transform 1 0 30452 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1476_
timestamp 1644511149
transform 1 0 30084 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1477_
timestamp 1644511149
transform 1 0 32200 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1478_
timestamp 1644511149
transform 1 0 31924 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1479_
timestamp 1644511149
transform 1 0 33212 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1480_
timestamp 1644511149
transform 1 0 32292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1481_
timestamp 1644511149
transform 1 0 30360 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1482_
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1483_
timestamp 1644511149
transform 1 0 32936 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1484_
timestamp 1644511149
transform 1 0 31004 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1485_
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1486_
timestamp 1644511149
transform 1 0 35604 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1487_
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1488_
timestamp 1644511149
transform 1 0 34408 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1489_
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1490_
timestamp 1644511149
transform 1 0 35604 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1491_
timestamp 1644511149
transform 1 0 35788 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1492_
timestamp 1644511149
transform 1 0 36248 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1493_
timestamp 1644511149
transform 1 0 32844 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1494_
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1495_
timestamp 1644511149
transform 1 0 21896 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _1496_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1497_
timestamp 1644511149
transform 1 0 26220 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1498_
timestamp 1644511149
transform 1 0 28704 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1499_
timestamp 1644511149
transform 1 0 15548 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1500_
timestamp 1644511149
transform 1 0 9292 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1501_
timestamp 1644511149
transform 1 0 17112 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1502_
timestamp 1644511149
transform 1 0 17112 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1503_
timestamp 1644511149
transform 1 0 16744 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1504_
timestamp 1644511149
transform 1 0 13340 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1505_
timestamp 1644511149
transform 1 0 17664 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1506_
timestamp 1644511149
transform 1 0 17296 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1507_
timestamp 1644511149
transform 1 0 17204 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1508_
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1509_
timestamp 1644511149
transform 1 0 14536 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1510_
timestamp 1644511149
transform 1 0 14260 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1511_
timestamp 1644511149
transform 1 0 12512 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1512_
timestamp 1644511149
transform 1 0 12880 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1513_
timestamp 1644511149
transform 1 0 11868 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1514_
timestamp 1644511149
transform 1 0 12788 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1515_
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1516_
timestamp 1644511149
transform 1 0 12788 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1517_
timestamp 1644511149
transform 1 0 23460 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _1518_
timestamp 1644511149
transform 1 0 15732 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1519_
timestamp 1644511149
transform 1 0 14720 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1520_
timestamp 1644511149
transform 1 0 23460 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1521_
timestamp 1644511149
transform 1 0 23276 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1522_
timestamp 1644511149
transform 1 0 19688 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1523_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14904 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1524_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15088 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1525_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14628 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1526_
timestamp 1644511149
transform 1 0 14444 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1527_
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1528_
timestamp 1644511149
transform 1 0 16468 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1529_
timestamp 1644511149
transform 1 0 15364 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1530_
timestamp 1644511149
transform 1 0 15088 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1531_
timestamp 1644511149
transform 1 0 17020 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1532_
timestamp 1644511149
transform 1 0 15456 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1533_
timestamp 1644511149
transform 1 0 15916 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1534_
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1535_
timestamp 1644511149
transform 1 0 15272 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1536_
timestamp 1644511149
transform 1 0 14352 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1537_
timestamp 1644511149
transform 1 0 14812 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1538_
timestamp 1644511149
transform 1 0 17848 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1539_
timestamp 1644511149
transform 1 0 15732 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1540_
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1541_
timestamp 1644511149
transform 1 0 15732 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1542_
timestamp 1644511149
transform 1 0 14720 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1543_
timestamp 1644511149
transform 1 0 17296 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1544_
timestamp 1644511149
transform 1 0 18492 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1545_
timestamp 1644511149
transform 1 0 19872 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1546_
timestamp 1644511149
transform 1 0 19504 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1547_
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1548_
timestamp 1644511149
transform 1 0 20148 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1549_
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1550_
timestamp 1644511149
transform 1 0 18308 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1551_
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1552_
timestamp 1644511149
transform 1 0 18124 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1553_
timestamp 1644511149
transform 1 0 16744 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1554_
timestamp 1644511149
transform 1 0 16744 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1555_
timestamp 1644511149
transform 1 0 20516 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1556_
timestamp 1644511149
transform 1 0 20148 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1557_
timestamp 1644511149
transform 1 0 22632 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1558_
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1559_
timestamp 1644511149
transform 1 0 18584 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1560_
timestamp 1644511149
transform 1 0 17940 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1561_
timestamp 1644511149
transform 1 0 15732 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1562_
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1563_
timestamp 1644511149
transform 1 0 23276 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1564_
timestamp 1644511149
transform 1 0 21896 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1565_
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1566_
timestamp 1644511149
transform 1 0 19780 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1567_
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1568_
timestamp 1644511149
transform 1 0 18308 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1569_
timestamp 1644511149
transform 1 0 17664 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1570_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20424 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1571_
timestamp 1644511149
transform 1 0 18952 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1572_
timestamp 1644511149
transform 1 0 18124 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1573_
timestamp 1644511149
transform 1 0 17296 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1574_
timestamp 1644511149
transform 1 0 16836 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1575_
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1576_
timestamp 1644511149
transform 1 0 20792 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1577_
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1578_
timestamp 1644511149
transform 1 0 20240 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1579_
timestamp 1644511149
transform 1 0 19136 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1580_
timestamp 1644511149
transform 1 0 17480 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1581_
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1582_
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1583_
timestamp 1644511149
transform 1 0 23000 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1584_
timestamp 1644511149
transform 1 0 21712 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1585_
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1586_
timestamp 1644511149
transform 1 0 21252 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1587_
timestamp 1644511149
transform 1 0 20884 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1588_
timestamp 1644511149
transform 1 0 22908 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1589_
timestamp 1644511149
transform 1 0 20240 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1590_
timestamp 1644511149
transform 1 0 22908 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1591_
timestamp 1644511149
transform 1 0 23368 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1592_
timestamp 1644511149
transform 1 0 22816 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1593_
timestamp 1644511149
transform 1 0 23092 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1594_
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1595_
timestamp 1644511149
transform 1 0 24196 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1596_
timestamp 1644511149
transform 1 0 21528 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1597_
timestamp 1644511149
transform 1 0 21896 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1598_
timestamp 1644511149
transform 1 0 22080 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1599_
timestamp 1644511149
transform 1 0 22448 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1600_
timestamp 1644511149
transform 1 0 23276 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1601_
timestamp 1644511149
transform 1 0 20516 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1602_
timestamp 1644511149
transform 1 0 20516 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1603_
timestamp 1644511149
transform 1 0 20700 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1604_
timestamp 1644511149
transform 1 0 20884 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1605_
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1606_
timestamp 1644511149
transform 1 0 22632 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1607_
timestamp 1644511149
transform 1 0 23000 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1608_
timestamp 1644511149
transform 1 0 24196 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1609_
timestamp 1644511149
transform 1 0 25208 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1610_
timestamp 1644511149
transform 1 0 25208 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1611_
timestamp 1644511149
transform 1 0 23644 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1612_
timestamp 1644511149
transform 1 0 24656 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1613_
timestamp 1644511149
transform 1 0 24564 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1614_
timestamp 1644511149
transform 1 0 22816 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1615_
timestamp 1644511149
transform 1 0 25484 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1616_
timestamp 1644511149
transform 1 0 24288 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1617_
timestamp 1644511149
transform 1 0 25668 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1618_
timestamp 1644511149
transform 1 0 26680 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1619_
timestamp 1644511149
transform 1 0 26864 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1620_
timestamp 1644511149
transform 1 0 21896 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1621_
timestamp 1644511149
transform 1 0 25944 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1622_
timestamp 1644511149
transform 1 0 25852 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1623_
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1624_
timestamp 1644511149
transform 1 0 27784 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1625_
timestamp 1644511149
transform 1 0 23460 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1626_
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1627_
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1628_
timestamp 1644511149
transform 1 0 27968 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1629_
timestamp 1644511149
transform 1 0 27508 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1630_
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1631_
timestamp 1644511149
transform 1 0 25576 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1632_
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1633_
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1634_
timestamp 1644511149
transform 1 0 28244 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1635_
timestamp 1644511149
transform 1 0 23552 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1636_
timestamp 1644511149
transform 1 0 24656 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1637_
timestamp 1644511149
transform 1 0 24932 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1638_
timestamp 1644511149
transform 1 0 25944 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1639_
timestamp 1644511149
transform 1 0 26036 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1640_
timestamp 1644511149
transform 1 0 24104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1641_
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1642_
timestamp 1644511149
transform 1 0 23368 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1643_
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1644_
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1645_
timestamp 1644511149
transform 1 0 26036 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1646_
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _1647_
timestamp 1644511149
transform 1 0 16376 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1648_
timestamp 1644511149
transform 1 0 26128 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1649_
timestamp 1644511149
transform 1 0 23092 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1650_
timestamp 1644511149
transform 1 0 23092 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1651_
timestamp 1644511149
transform 1 0 20608 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1652_
timestamp 1644511149
transform 1 0 24748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1653_
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1654_
timestamp 1644511149
transform 1 0 23644 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a221o_1  _1655_
timestamp 1644511149
transform 1 0 21988 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1656_
timestamp 1644511149
transform 1 0 26036 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1657_
timestamp 1644511149
transform 1 0 23368 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1658_
timestamp 1644511149
transform 1 0 23920 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1659_
timestamp 1644511149
transform 1 0 25392 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1660_
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1661_
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1662_
timestamp 1644511149
transform 1 0 24380 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1663_
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1664_
timestamp 1644511149
transform 1 0 23184 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1665_
timestamp 1644511149
transform 1 0 23368 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1666_
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1667_
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1668_
timestamp 1644511149
transform 1 0 21988 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1669_
timestamp 1644511149
transform 1 0 26772 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1670_
timestamp 1644511149
transform 1 0 28152 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1671_
timestamp 1644511149
transform 1 0 28428 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1672_
timestamp 1644511149
transform 1 0 25484 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1673_
timestamp 1644511149
transform 1 0 27508 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1674_
timestamp 1644511149
transform 1 0 28244 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1675_
timestamp 1644511149
transform 1 0 28980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1676_
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1677_
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1678_
timestamp 1644511149
transform 1 0 28520 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1679_
timestamp 1644511149
transform 1 0 28152 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1680_
timestamp 1644511149
transform 1 0 26956 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1681_
timestamp 1644511149
transform 1 0 27508 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1682_
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1683_
timestamp 1644511149
transform 1 0 29624 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1684_
timestamp 1644511149
transform 1 0 25668 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1685_
timestamp 1644511149
transform 1 0 17388 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1686_
timestamp 1644511149
transform 1 0 18124 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1687_
timestamp 1644511149
transform 1 0 16560 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1688_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1689_
timestamp 1644511149
transform 1 0 7820 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1690_
timestamp 1644511149
transform 1 0 10304 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1691_
timestamp 1644511149
transform 1 0 7820 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1692_
timestamp 1644511149
transform 1 0 10396 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1693_
timestamp 1644511149
transform 1 0 6992 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1694_
timestamp 1644511149
transform 1 0 10396 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1695_
timestamp 1644511149
transform 1 0 7820 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1696_
timestamp 1644511149
transform 1 0 7820 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1697_
timestamp 1644511149
transform 1 0 10396 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1698_
timestamp 1644511149
transform 1 0 8464 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1699_
timestamp 1644511149
transform 1 0 17296 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1700_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14536 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1701_
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1702_
timestamp 1644511149
transform 1 0 17020 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1703_
timestamp 1644511149
transform 1 0 17020 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1704_
timestamp 1644511149
transform 1 0 17296 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1705_
timestamp 1644511149
transform 1 0 18124 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1706_
timestamp 1644511149
transform 1 0 19320 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1707_
timestamp 1644511149
transform 1 0 19872 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1708_
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1709_
timestamp 1644511149
transform 1 0 21804 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1710_
timestamp 1644511149
transform 1 0 22448 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1711_
timestamp 1644511149
transform 1 0 22264 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1712_
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1713_
timestamp 1644511149
transform 1 0 24932 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 1644511149
transform 1 0 25760 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 1644511149
transform 1 0 25208 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1716_
timestamp 1644511149
transform 1 0 24932 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1717_
timestamp 1644511149
transform 1 0 23276 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1718_
timestamp 1644511149
transform 1 0 13156 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1719_
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 1644511149
transform 1 0 10580 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1721_
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1722_
timestamp 1644511149
transform 1 0 8280 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1723_
timestamp 1644511149
transform 1 0 3864 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1724_
timestamp 1644511149
transform 1 0 3956 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1725_
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1726_
timestamp 1644511149
transform 1 0 3864 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1727_
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1728_
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1729_
timestamp 1644511149
transform 1 0 5244 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1730_
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1731_
timestamp 1644511149
transform 1 0 5796 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1732_
timestamp 1644511149
transform 1 0 6624 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1733_
timestamp 1644511149
transform 1 0 8188 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1734_
timestamp 1644511149
transform 1 0 7360 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1735_
timestamp 1644511149
transform 1 0 8740 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1736_
timestamp 1644511149
transform 1 0 9200 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1737_
timestamp 1644511149
transform 1 0 8832 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1738_
timestamp 1644511149
transform 1 0 9200 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1739_
timestamp 1644511149
transform 1 0 10304 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1740_
timestamp 1644511149
transform 1 0 10396 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1741_
timestamp 1644511149
transform 1 0 10304 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1742_
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1743_
timestamp 1644511149
transform 1 0 11868 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1744_
timestamp 1644511149
transform 1 0 11776 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1745_
timestamp 1644511149
transform 1 0 12144 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1746_
timestamp 1644511149
transform 1 0 13616 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1747_
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1748_
timestamp 1644511149
transform 1 0 14812 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1749_
timestamp 1644511149
transform 1 0 14720 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1750_
timestamp 1644511149
transform 1 0 15088 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1751_
timestamp 1644511149
transform 1 0 17848 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1752_
timestamp 1644511149
transform 1 0 12696 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1753_
timestamp 1644511149
transform 1 0 14536 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1754_
timestamp 1644511149
transform 1 0 11684 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1755_
timestamp 1644511149
transform 1 0 12144 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1756_
timestamp 1644511149
transform 1 0 8464 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1757_
timestamp 1644511149
transform 1 0 6624 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1758_
timestamp 1644511149
transform 1 0 7268 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1759_
timestamp 1644511149
transform 1 0 6992 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1760_
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1761_
timestamp 1644511149
transform 1 0 9200 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1762_
timestamp 1644511149
transform 1 0 10672 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1763_
timestamp 1644511149
transform 1 0 19044 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1764_
timestamp 1644511149
transform 1 0 19228 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1765_
timestamp 1644511149
transform 1 0 19780 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1766_
timestamp 1644511149
transform 1 0 20056 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1767_
timestamp 1644511149
transform 1 0 19780 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1768_
timestamp 1644511149
transform 1 0 22448 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1769_
timestamp 1644511149
transform 1 0 22356 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1770_
timestamp 1644511149
transform 1 0 21620 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1771_
timestamp 1644511149
transform 1 0 24472 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1772_
timestamp 1644511149
transform 1 0 23920 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1773_
timestamp 1644511149
transform 1 0 27416 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1774_
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1775_
timestamp 1644511149
transform 1 0 27600 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1776_
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1777_
timestamp 1644511149
transform 1 0 26680 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1778_
timestamp 1644511149
transform 1 0 24564 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1779_
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1780_
timestamp 1644511149
transform 1 0 19780 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1781_
timestamp 1644511149
transform 1 0 19872 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1782_
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1783_
timestamp 1644511149
transform 1 0 19596 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1784_
timestamp 1644511149
transform 1 0 23644 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1785_
timestamp 1644511149
transform 1 0 22080 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1786_
timestamp 1644511149
transform 1 0 21896 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1787_
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1788_
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1789_
timestamp 1644511149
transform 1 0 27324 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1790_
timestamp 1644511149
transform 1 0 24840 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1791_
timestamp 1644511149
transform 1 0 27600 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1792_
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1793_
timestamp 1644511149
transform 1 0 21988 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1794_
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1795_
timestamp 1644511149
transform 1 0 27416 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1796_
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1797_
timestamp 1644511149
transform 1 0 29256 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1798_
timestamp 1644511149
transform 1 0 27140 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1799_
timestamp 1644511149
transform 1 0 29716 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1800_
timestamp 1644511149
transform 1 0 29716 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1801_
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1802_
timestamp 1644511149
transform 1 0 30084 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1803_
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1804_
timestamp 1644511149
transform 1 0 30084 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1805_
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1806_
timestamp 1644511149
transform 1 0 33672 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1807_
timestamp 1644511149
transform 1 0 34408 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1808_
timestamp 1644511149
transform 1 0 33764 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1809_
timestamp 1644511149
transform 1 0 33948 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1810_
timestamp 1644511149
transform 1 0 32292 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1811_
timestamp 1644511149
transform 1 0 15824 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1812_
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1813_
timestamp 1644511149
transform 1 0 14168 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1814_
timestamp 1644511149
transform 1 0 16836 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1815_
timestamp 1644511149
transform 1 0 18216 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1816_
timestamp 1644511149
transform 1 0 17296 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1817_
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1818_
timestamp 1644511149
transform 1 0 10580 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1819_
timestamp 1644511149
transform 1 0 8648 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1820_
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1821_
timestamp 1644511149
transform 1 0 15456 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1822_
timestamp 1644511149
transform 1 0 17848 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1823_
timestamp 1644511149
transform 1 0 14168 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1644511149
transform 1 0 14628 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1644511149
transform 1 0 16468 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1644511149
transform 1 0 14076 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1644511149
transform 1 0 16100 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1828_
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1644511149
transform 1 0 16376 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1644511149
transform 1 0 18308 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1831_
timestamp 1644511149
transform 1 0 16928 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1832_
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1833_
timestamp 1644511149
transform 1 0 20516 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1834_
timestamp 1644511149
transform 1 0 23368 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1835_
timestamp 1644511149
transform 1 0 22356 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1836_
timestamp 1644511149
transform 1 0 21068 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1837_
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1838_
timestamp 1644511149
transform 1 0 26864 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1839_
timestamp 1644511149
transform 1 0 27140 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1840_
timestamp 1644511149
transform 1 0 27140 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1841_
timestamp 1644511149
transform 1 0 26404 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1842_
timestamp 1644511149
transform 1 0 25024 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1843_
timestamp 1644511149
transform 1 0 23644 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1844_
timestamp 1644511149
transform 1 0 20608 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1845_
timestamp 1644511149
transform 1 0 20148 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1846_
timestamp 1644511149
transform 1 0 24472 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1847_
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1848_
timestamp 1644511149
transform 1 0 24656 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1849_
timestamp 1644511149
transform 1 0 23644 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1850_
timestamp 1644511149
transform 1 0 23644 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1851_
timestamp 1644511149
transform 1 0 21528 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1852_
timestamp 1644511149
transform 1 0 27508 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1853_
timestamp 1644511149
transform 1 0 24748 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1854_
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1855_
timestamp 1644511149
transform 1 0 27416 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1856_
timestamp 1644511149
transform 1 0 28796 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1857_
timestamp 1644511149
transform 1 0 27600 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1858_
timestamp 1644511149
transform 1 0 28520 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1859_
timestamp 1644511149
transform 1 0 25668 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1860_
timestamp 1644511149
transform 1 0 17204 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1861_
timestamp 1644511149
transform 1 0 17204 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1862__90 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1863__91
timestamp 1644511149
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CLK pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19596 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_CLK
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_CLK
timestamp 1644511149
transform 1 0 11776 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_CLK
timestamp 1644511149
transform 1 0 12880 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_CLK
timestamp 1644511149
transform 1 0 15364 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_CLK
timestamp 1644511149
transform 1 0 23276 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_CLK
timestamp 1644511149
transform 1 0 26680 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_CLK
timestamp 1644511149
transform 1 0 21252 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_CLK
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_CLK
timestamp 1644511149
transform 1 0 10856 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_CLK
timestamp 1644511149
transform 1 0 10120 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_CLK
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_CLK
timestamp 1644511149
transform 1 0 10672 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_CLK
timestamp 1644511149
transform 1 0 12512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_CLK
timestamp 1644511149
transform 1 0 10672 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_CLK
timestamp 1644511149
transform 1 0 15824 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_CLK
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_CLK
timestamp 1644511149
transform 1 0 23276 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_CLK
timestamp 1644511149
transform 1 0 23276 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_CLK
timestamp 1644511149
transform 1 0 27508 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_CLK
timestamp 1644511149
transform 1 0 27416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_CLK
timestamp 1644511149
transform 1 0 20976 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_CLK
timestamp 1644511149
transform 1 0 20976 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_CLK
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_CLK
timestamp 1644511149
transform 1 0 25300 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 3680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1644511149
transform 1 0 2392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform 1 0 2392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 3220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1644511149
transform 1 0 2392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform 1 0 2576 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1644511149
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1644511149
transform 1 0 4692 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform 1 0 1932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform 1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1644511149
transform 1 0 2944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform 1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform 1 0 2300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1644511149
transform 1 0 1748 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform 1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform 1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform 1 0 2392 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 2208 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 1564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1644511149
transform 1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1644511149
transform 1 0 4324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 2392 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 2944 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 4324 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform 1 0 1748 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 3680 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1644511149
transform 1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1644511149
transform 1 0 3036 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1644511149
transform 1 0 29716 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1644511149
transform 1 0 31464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1644511149
transform 1 0 30360 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1644511149
transform 1 0 30360 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1644511149
transform 1 0 31096 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1644511149
transform 1 0 31004 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform 1 0 31004 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1644511149
transform 1 0 29992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1644511149
transform 1 0 31004 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1644511149
transform 1 0 31648 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1644511149
transform 1 0 30176 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform 1 0 30636 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input52
timestamp 1644511149
transform 1 0 36064 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input53
timestamp 1644511149
transform 1 0 4140 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1644511149
transform 1 0 23552 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1644511149
transform 1 0 26404 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1644511149
transform 1 0 30268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1644511149
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1644511149
transform 1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1644511149
transform 1 0 19964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1644511149
transform 1 0 32844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1644511149
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1644511149
transform 1 0 34592 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1644511149
transform 1 0 35420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1644511149
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1644511149
transform 1 0 37628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1644511149
transform 1 0 37812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1644511149
transform 1 0 37812 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1644511149
transform 1 0 37812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1644511149
transform 1 0 22448 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1644511149
transform 1 0 23644 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1644511149
transform 1 0 22540 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1644511149
transform 1 0 23184 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1644511149
transform 1 0 25116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1644511149
transform 1 0 12052 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1644511149
transform 1 0 20056 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 406 592
<< labels >>
rlabel metal2 s 202 0 258 800 6 CLK
port 0 nsew signal input
rlabel metal2 s 570 0 626 800 6 RST_N
port 1 nsew signal input
rlabel metal2 s 3146 0 3202 800 6 slave_ack_o
port 2 nsew signal tristate
rlabel metal2 s 4250 0 4306 800 6 slave_adr_i[0]
port 3 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 slave_adr_i[10]
port 4 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 slave_adr_i[11]
port 5 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 slave_adr_i[12]
port 6 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 slave_adr_i[13]
port 7 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 slave_adr_i[14]
port 8 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 slave_adr_i[15]
port 9 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 slave_adr_i[16]
port 10 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 slave_adr_i[17]
port 11 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 slave_adr_i[18]
port 12 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 slave_adr_i[19]
port 13 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 slave_adr_i[1]
port 14 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 slave_adr_i[20]
port 15 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 slave_adr_i[21]
port 16 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 slave_adr_i[22]
port 17 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 slave_adr_i[23]
port 18 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 slave_adr_i[24]
port 19 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 slave_adr_i[25]
port 20 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 slave_adr_i[26]
port 21 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 slave_adr_i[27]
port 22 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 slave_adr_i[28]
port 23 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 slave_adr_i[29]
port 24 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 slave_adr_i[2]
port 25 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 slave_adr_i[30]
port 26 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 slave_adr_i[31]
port 27 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 slave_adr_i[3]
port 28 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 slave_adr_i[4]
port 29 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 slave_adr_i[5]
port 30 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 slave_adr_i[6]
port 31 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 slave_adr_i[7]
port 32 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 slave_adr_i[8]
port 33 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 slave_adr_i[9]
port 34 nsew signal input
rlabel metal2 s 938 0 994 800 6 slave_cyc_i
port 35 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 slave_dat_i[0]
port 36 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 slave_dat_i[10]
port 37 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 slave_dat_i[11]
port 38 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 slave_dat_i[12]
port 39 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 slave_dat_i[13]
port 40 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 slave_dat_i[14]
port 41 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 slave_dat_i[15]
port 42 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 slave_dat_i[16]
port 43 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 slave_dat_i[17]
port 44 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 slave_dat_i[18]
port 45 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 slave_dat_i[19]
port 46 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 slave_dat_i[1]
port 47 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 slave_dat_i[20]
port 48 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 slave_dat_i[21]
port 49 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 slave_dat_i[22]
port 50 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 slave_dat_i[23]
port 51 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 slave_dat_i[24]
port 52 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 slave_dat_i[25]
port 53 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 slave_dat_i[26]
port 54 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 slave_dat_i[27]
port 55 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 slave_dat_i[28]
port 56 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 slave_dat_i[29]
port 57 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 slave_dat_i[2]
port 58 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 slave_dat_i[30]
port 59 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 slave_dat_i[31]
port 60 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 slave_dat_i[3]
port 61 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 slave_dat_i[4]
port 62 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 slave_dat_i[5]
port 63 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 slave_dat_i[6]
port 64 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 slave_dat_i[7]
port 65 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 slave_dat_i[8]
port 66 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 slave_dat_i[9]
port 67 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 slave_dat_o[0]
port 68 nsew signal tristate
rlabel metal2 s 24122 0 24178 800 6 slave_dat_o[10]
port 69 nsew signal tristate
rlabel metal2 s 24858 0 24914 800 6 slave_dat_o[11]
port 70 nsew signal tristate
rlabel metal2 s 25594 0 25650 800 6 slave_dat_o[12]
port 71 nsew signal tristate
rlabel metal2 s 26330 0 26386 800 6 slave_dat_o[13]
port 72 nsew signal tristate
rlabel metal2 s 27066 0 27122 800 6 slave_dat_o[14]
port 73 nsew signal tristate
rlabel metal2 s 27802 0 27858 800 6 slave_dat_o[15]
port 74 nsew signal tristate
rlabel metal2 s 28538 0 28594 800 6 slave_dat_o[16]
port 75 nsew signal tristate
rlabel metal2 s 29366 0 29422 800 6 slave_dat_o[17]
port 76 nsew signal tristate
rlabel metal2 s 30102 0 30158 800 6 slave_dat_o[18]
port 77 nsew signal tristate
rlabel metal2 s 30838 0 30894 800 6 slave_dat_o[19]
port 78 nsew signal tristate
rlabel metal2 s 17406 0 17462 800 6 slave_dat_o[1]
port 79 nsew signal tristate
rlabel metal2 s 31574 0 31630 800 6 slave_dat_o[20]
port 80 nsew signal tristate
rlabel metal2 s 32310 0 32366 800 6 slave_dat_o[21]
port 81 nsew signal tristate
rlabel metal2 s 33046 0 33102 800 6 slave_dat_o[22]
port 82 nsew signal tristate
rlabel metal2 s 33782 0 33838 800 6 slave_dat_o[23]
port 83 nsew signal tristate
rlabel metal2 s 34610 0 34666 800 6 slave_dat_o[24]
port 84 nsew signal tristate
rlabel metal2 s 35346 0 35402 800 6 slave_dat_o[25]
port 85 nsew signal tristate
rlabel metal2 s 36082 0 36138 800 6 slave_dat_o[26]
port 86 nsew signal tristate
rlabel metal2 s 36818 0 36874 800 6 slave_dat_o[27]
port 87 nsew signal tristate
rlabel metal2 s 37554 0 37610 800 6 slave_dat_o[28]
port 88 nsew signal tristate
rlabel metal2 s 38290 0 38346 800 6 slave_dat_o[29]
port 89 nsew signal tristate
rlabel metal2 s 18142 0 18198 800 6 slave_dat_o[2]
port 90 nsew signal tristate
rlabel metal2 s 39026 0 39082 800 6 slave_dat_o[30]
port 91 nsew signal tristate
rlabel metal2 s 39762 0 39818 800 6 slave_dat_o[31]
port 92 nsew signal tristate
rlabel metal2 s 18878 0 18934 800 6 slave_dat_o[3]
port 93 nsew signal tristate
rlabel metal2 s 19614 0 19670 800 6 slave_dat_o[4]
port 94 nsew signal tristate
rlabel metal2 s 20350 0 20406 800 6 slave_dat_o[5]
port 95 nsew signal tristate
rlabel metal2 s 21086 0 21142 800 6 slave_dat_o[6]
port 96 nsew signal tristate
rlabel metal2 s 21822 0 21878 800 6 slave_dat_o[7]
port 97 nsew signal tristate
rlabel metal2 s 22558 0 22614 800 6 slave_dat_o[8]
port 98 nsew signal tristate
rlabel metal2 s 23386 0 23442 800 6 slave_dat_o[9]
port 99 nsew signal tristate
rlabel metal2 s 3514 0 3570 800 6 slave_err_o
port 100 nsew signal tristate
rlabel metal2 s 3882 0 3938 800 6 slave_rty_o
port 101 nsew signal tristate
rlabel metal2 s 1674 0 1730 800 6 slave_sel_i[0]
port 102 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 slave_sel_i[1]
port 103 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 slave_sel_i[2]
port 104 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 slave_sel_i[3]
port 105 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 slave_stb_i
port 106 nsew signal input
rlabel metal2 s 35990 49200 36046 50000 6 slave_we_i
port 107 nsew signal input
rlabel metal2 s 3974 49200 4030 50000 6 spiMaster_miso
port 108 nsew signal input
rlabel metal2 s 11978 49200 12034 50000 6 spiMaster_mosi
port 109 nsew signal tristate
rlabel metal2 s 19982 49200 20038 50000 6 spiMaster_mosi_oe
port 110 nsew signal tristate
rlabel metal2 s 27986 49200 28042 50000 6 spiMaster_sclk
port 111 nsew signal tristate
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 112 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 112 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 113 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 40000 50000
<< end >>
