VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mkLanaiCPU
  CLASS BLOCK ;
  FOREIGN mkLanaiCPU ;
  ORIGIN 0.000 0.000 ;
  SIZE 840.545 BY 851.265 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END CLK
  PIN EN_dmem_client_request_get
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 847.265 2.210 851.265 ;
    END
  END EN_dmem_client_request_get
  PIN EN_dmem_client_response_put
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 847.265 5.890 851.265 ;
    END
  END EN_dmem_client_response_put
  PIN EN_imem_client_request_get
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 847.265 538.570 851.265 ;
    END
  END EN_imem_client_request_get
  PIN EN_imem_client_response_put
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 847.265 542.710 851.265 ;
    END
  END EN_imem_client_response_put
  PIN RDY_dmem_client_request_get
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 847.265 10.030 851.265 ;
    END
  END RDY_dmem_client_request_get
  PIN RDY_dmem_client_response_put
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 847.265 13.710 851.265 ;
    END
  END RDY_dmem_client_response_put
  PIN RDY_imem_client_request_get
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 847.265 546.390 851.265 ;
    END
  END RDY_imem_client_request_get
  PIN RDY_imem_client_response_put
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 847.265 550.530 851.265 ;
    END
  END RDY_imem_client_response_put
  PIN RDY_readPC
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END RDY_readPC
  PIN RST_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END RST_N
  PIN dmem_client_request_get[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 847.265 17.850 851.265 ;
    END
  END dmem_client_request_get[0]
  PIN dmem_client_request_get[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 847.265 96.510 851.265 ;
    END
  END dmem_client_request_get[10]
  PIN dmem_client_request_get[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 847.265 104.790 851.265 ;
    END
  END dmem_client_request_get[11]
  PIN dmem_client_request_get[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 847.265 112.610 851.265 ;
    END
  END dmem_client_request_get[12]
  PIN dmem_client_request_get[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 847.265 120.430 851.265 ;
    END
  END dmem_client_request_get[13]
  PIN dmem_client_request_get[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 847.265 128.250 851.265 ;
    END
  END dmem_client_request_get[14]
  PIN dmem_client_request_get[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 847.265 136.070 851.265 ;
    END
  END dmem_client_request_get[15]
  PIN dmem_client_request_get[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 847.265 143.890 851.265 ;
    END
  END dmem_client_request_get[16]
  PIN dmem_client_request_get[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 847.265 151.710 851.265 ;
    END
  END dmem_client_request_get[17]
  PIN dmem_client_request_get[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 847.265 159.990 851.265 ;
    END
  END dmem_client_request_get[18]
  PIN dmem_client_request_get[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 847.265 167.810 851.265 ;
    END
  END dmem_client_request_get[19]
  PIN dmem_client_request_get[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 847.265 25.670 851.265 ;
    END
  END dmem_client_request_get[1]
  PIN dmem_client_request_get[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 847.265 175.630 851.265 ;
    END
  END dmem_client_request_get[20]
  PIN dmem_client_request_get[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 847.265 183.450 851.265 ;
    END
  END dmem_client_request_get[21]
  PIN dmem_client_request_get[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 847.265 191.270 851.265 ;
    END
  END dmem_client_request_get[22]
  PIN dmem_client_request_get[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 847.265 199.090 851.265 ;
    END
  END dmem_client_request_get[23]
  PIN dmem_client_request_get[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 847.265 207.370 851.265 ;
    END
  END dmem_client_request_get[24]
  PIN dmem_client_request_get[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 847.265 215.190 851.265 ;
    END
  END dmem_client_request_get[25]
  PIN dmem_client_request_get[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 847.265 223.010 851.265 ;
    END
  END dmem_client_request_get[26]
  PIN dmem_client_request_get[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 847.265 230.830 851.265 ;
    END
  END dmem_client_request_get[27]
  PIN dmem_client_request_get[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 847.265 238.650 851.265 ;
    END
  END dmem_client_request_get[28]
  PIN dmem_client_request_get[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 847.265 246.470 851.265 ;
    END
  END dmem_client_request_get[29]
  PIN dmem_client_request_get[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 847.265 33.490 851.265 ;
    END
  END dmem_client_request_get[2]
  PIN dmem_client_request_get[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 847.265 254.290 851.265 ;
    END
  END dmem_client_request_get[30]
  PIN dmem_client_request_get[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 847.265 262.570 851.265 ;
    END
  END dmem_client_request_get[31]
  PIN dmem_client_request_get[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 847.265 270.390 851.265 ;
    END
  END dmem_client_request_get[32]
  PIN dmem_client_request_get[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 847.265 274.070 851.265 ;
    END
  END dmem_client_request_get[33]
  PIN dmem_client_request_get[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 847.265 278.210 851.265 ;
    END
  END dmem_client_request_get[34]
  PIN dmem_client_request_get[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 847.265 282.350 851.265 ;
    END
  END dmem_client_request_get[35]
  PIN dmem_client_request_get[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 847.265 286.030 851.265 ;
    END
  END dmem_client_request_get[36]
  PIN dmem_client_request_get[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 847.265 290.170 851.265 ;
    END
  END dmem_client_request_get[37]
  PIN dmem_client_request_get[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 847.265 293.850 851.265 ;
    END
  END dmem_client_request_get[38]
  PIN dmem_client_request_get[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 847.265 297.990 851.265 ;
    END
  END dmem_client_request_get[39]
  PIN dmem_client_request_get[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 847.265 41.310 851.265 ;
    END
  END dmem_client_request_get[3]
  PIN dmem_client_request_get[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 847.265 301.670 851.265 ;
    END
  END dmem_client_request_get[40]
  PIN dmem_client_request_get[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 847.265 305.810 851.265 ;
    END
  END dmem_client_request_get[41]
  PIN dmem_client_request_get[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 847.265 309.950 851.265 ;
    END
  END dmem_client_request_get[42]
  PIN dmem_client_request_get[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 847.265 313.630 851.265 ;
    END
  END dmem_client_request_get[43]
  PIN dmem_client_request_get[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 847.265 317.770 851.265 ;
    END
  END dmem_client_request_get[44]
  PIN dmem_client_request_get[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 847.265 321.450 851.265 ;
    END
  END dmem_client_request_get[45]
  PIN dmem_client_request_get[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 847.265 325.590 851.265 ;
    END
  END dmem_client_request_get[46]
  PIN dmem_client_request_get[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 847.265 329.270 851.265 ;
    END
  END dmem_client_request_get[47]
  PIN dmem_client_request_get[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 847.265 333.410 851.265 ;
    END
  END dmem_client_request_get[48]
  PIN dmem_client_request_get[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 847.265 337.550 851.265 ;
    END
  END dmem_client_request_get[49]
  PIN dmem_client_request_get[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 847.265 49.130 851.265 ;
    END
  END dmem_client_request_get[4]
  PIN dmem_client_request_get[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 847.265 341.230 851.265 ;
    END
  END dmem_client_request_get[50]
  PIN dmem_client_request_get[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 847.265 345.370 851.265 ;
    END
  END dmem_client_request_get[51]
  PIN dmem_client_request_get[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 847.265 349.050 851.265 ;
    END
  END dmem_client_request_get[52]
  PIN dmem_client_request_get[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 847.265 353.190 851.265 ;
    END
  END dmem_client_request_get[53]
  PIN dmem_client_request_get[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.590 847.265 356.870 851.265 ;
    END
  END dmem_client_request_get[54]
  PIN dmem_client_request_get[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 847.265 361.010 851.265 ;
    END
  END dmem_client_request_get[55]
  PIN dmem_client_request_get[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 847.265 365.150 851.265 ;
    END
  END dmem_client_request_get[56]
  PIN dmem_client_request_get[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 847.265 368.830 851.265 ;
    END
  END dmem_client_request_get[57]
  PIN dmem_client_request_get[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 847.265 372.970 851.265 ;
    END
  END dmem_client_request_get[58]
  PIN dmem_client_request_get[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 847.265 376.650 851.265 ;
    END
  END dmem_client_request_get[59]
  PIN dmem_client_request_get[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 847.265 57.410 851.265 ;
    END
  END dmem_client_request_get[5]
  PIN dmem_client_request_get[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 847.265 380.790 851.265 ;
    END
  END dmem_client_request_get[60]
  PIN dmem_client_request_get[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 847.265 384.930 851.265 ;
    END
  END dmem_client_request_get[61]
  PIN dmem_client_request_get[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 847.265 388.610 851.265 ;
    END
  END dmem_client_request_get[62]
  PIN dmem_client_request_get[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 847.265 392.750 851.265 ;
    END
  END dmem_client_request_get[63]
  PIN dmem_client_request_get[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 847.265 396.430 851.265 ;
    END
  END dmem_client_request_get[64]
  PIN dmem_client_request_get[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 847.265 400.570 851.265 ;
    END
  END dmem_client_request_get[65]
  PIN dmem_client_request_get[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 847.265 404.250 851.265 ;
    END
  END dmem_client_request_get[66]
  PIN dmem_client_request_get[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 847.265 408.390 851.265 ;
    END
  END dmem_client_request_get[67]
  PIN dmem_client_request_get[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 847.265 412.530 851.265 ;
    END
  END dmem_client_request_get[68]
  PIN dmem_client_request_get[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 847.265 416.210 851.265 ;
    END
  END dmem_client_request_get[69]
  PIN dmem_client_request_get[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 847.265 65.230 851.265 ;
    END
  END dmem_client_request_get[6]
  PIN dmem_client_request_get[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 847.265 420.350 851.265 ;
    END
  END dmem_client_request_get[70]
  PIN dmem_client_request_get[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 847.265 424.030 851.265 ;
    END
  END dmem_client_request_get[71]
  PIN dmem_client_request_get[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 847.265 428.170 851.265 ;
    END
  END dmem_client_request_get[72]
  PIN dmem_client_request_get[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 847.265 431.850 851.265 ;
    END
  END dmem_client_request_get[73]
  PIN dmem_client_request_get[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 847.265 435.990 851.265 ;
    END
  END dmem_client_request_get[74]
  PIN dmem_client_request_get[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 847.265 440.130 851.265 ;
    END
  END dmem_client_request_get[75]
  PIN dmem_client_request_get[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 847.265 443.810 851.265 ;
    END
  END dmem_client_request_get[76]
  PIN dmem_client_request_get[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 847.265 447.950 851.265 ;
    END
  END dmem_client_request_get[77]
  PIN dmem_client_request_get[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 847.265 451.630 851.265 ;
    END
  END dmem_client_request_get[78]
  PIN dmem_client_request_get[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 847.265 455.770 851.265 ;
    END
  END dmem_client_request_get[79]
  PIN dmem_client_request_get[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 847.265 73.050 851.265 ;
    END
  END dmem_client_request_get[7]
  PIN dmem_client_request_get[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.170 847.265 459.450 851.265 ;
    END
  END dmem_client_request_get[80]
  PIN dmem_client_request_get[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 847.265 463.590 851.265 ;
    END
  END dmem_client_request_get[81]
  PIN dmem_client_request_get[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 847.265 467.730 851.265 ;
    END
  END dmem_client_request_get[82]
  PIN dmem_client_request_get[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 847.265 471.410 851.265 ;
    END
  END dmem_client_request_get[83]
  PIN dmem_client_request_get[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 847.265 475.550 851.265 ;
    END
  END dmem_client_request_get[84]
  PIN dmem_client_request_get[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 847.265 479.230 851.265 ;
    END
  END dmem_client_request_get[85]
  PIN dmem_client_request_get[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 847.265 483.370 851.265 ;
    END
  END dmem_client_request_get[86]
  PIN dmem_client_request_get[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 847.265 487.510 851.265 ;
    END
  END dmem_client_request_get[87]
  PIN dmem_client_request_get[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 847.265 491.190 851.265 ;
    END
  END dmem_client_request_get[88]
  PIN dmem_client_request_get[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 847.265 495.330 851.265 ;
    END
  END dmem_client_request_get[89]
  PIN dmem_client_request_get[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 847.265 80.870 851.265 ;
    END
  END dmem_client_request_get[8]
  PIN dmem_client_request_get[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 847.265 499.010 851.265 ;
    END
  END dmem_client_request_get[90]
  PIN dmem_client_request_get[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 847.265 503.150 851.265 ;
    END
  END dmem_client_request_get[91]
  PIN dmem_client_request_get[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 847.265 506.830 851.265 ;
    END
  END dmem_client_request_get[92]
  PIN dmem_client_request_get[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 847.265 510.970 851.265 ;
    END
  END dmem_client_request_get[93]
  PIN dmem_client_request_get[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 847.265 515.110 851.265 ;
    END
  END dmem_client_request_get[94]
  PIN dmem_client_request_get[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 847.265 518.790 851.265 ;
    END
  END dmem_client_request_get[95]
  PIN dmem_client_request_get[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.650 847.265 522.930 851.265 ;
    END
  END dmem_client_request_get[96]
  PIN dmem_client_request_get[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 847.265 526.610 851.265 ;
    END
  END dmem_client_request_get[97]
  PIN dmem_client_request_get[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 847.265 530.750 851.265 ;
    END
  END dmem_client_request_get[98]
  PIN dmem_client_request_get[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 847.265 534.430 851.265 ;
    END
  END dmem_client_request_get[99]
  PIN dmem_client_request_get[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 847.265 88.690 851.265 ;
    END
  END dmem_client_request_get[9]
  PIN dmem_client_response_put[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 847.265 21.530 851.265 ;
    END
  END dmem_client_response_put[0]
  PIN dmem_client_response_put[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 847.265 100.650 851.265 ;
    END
  END dmem_client_response_put[10]
  PIN dmem_client_response_put[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 847.265 108.470 851.265 ;
    END
  END dmem_client_response_put[11]
  PIN dmem_client_response_put[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 847.265 116.290 851.265 ;
    END
  END dmem_client_response_put[12]
  PIN dmem_client_response_put[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 847.265 124.110 851.265 ;
    END
  END dmem_client_response_put[13]
  PIN dmem_client_response_put[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 847.265 132.390 851.265 ;
    END
  END dmem_client_response_put[14]
  PIN dmem_client_response_put[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 847.265 140.210 851.265 ;
    END
  END dmem_client_response_put[15]
  PIN dmem_client_response_put[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 847.265 148.030 851.265 ;
    END
  END dmem_client_response_put[16]
  PIN dmem_client_response_put[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 847.265 155.850 851.265 ;
    END
  END dmem_client_response_put[17]
  PIN dmem_client_response_put[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 847.265 163.670 851.265 ;
    END
  END dmem_client_response_put[18]
  PIN dmem_client_response_put[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 847.265 171.490 851.265 ;
    END
  END dmem_client_response_put[19]
  PIN dmem_client_response_put[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 847.265 29.810 851.265 ;
    END
  END dmem_client_response_put[1]
  PIN dmem_client_response_put[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 847.265 179.310 851.265 ;
    END
  END dmem_client_response_put[20]
  PIN dmem_client_response_put[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 847.265 187.590 851.265 ;
    END
  END dmem_client_response_put[21]
  PIN dmem_client_response_put[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 847.265 195.410 851.265 ;
    END
  END dmem_client_response_put[22]
  PIN dmem_client_response_put[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 847.265 203.230 851.265 ;
    END
  END dmem_client_response_put[23]
  PIN dmem_client_response_put[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 847.265 211.050 851.265 ;
    END
  END dmem_client_response_put[24]
  PIN dmem_client_response_put[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 847.265 218.870 851.265 ;
    END
  END dmem_client_response_put[25]
  PIN dmem_client_response_put[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 847.265 226.690 851.265 ;
    END
  END dmem_client_response_put[26]
  PIN dmem_client_response_put[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 847.265 234.970 851.265 ;
    END
  END dmem_client_response_put[27]
  PIN dmem_client_response_put[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 847.265 242.790 851.265 ;
    END
  END dmem_client_response_put[28]
  PIN dmem_client_response_put[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 847.265 250.610 851.265 ;
    END
  END dmem_client_response_put[29]
  PIN dmem_client_response_put[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 847.265 37.630 851.265 ;
    END
  END dmem_client_response_put[2]
  PIN dmem_client_response_put[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 847.265 258.430 851.265 ;
    END
  END dmem_client_response_put[30]
  PIN dmem_client_response_put[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 847.265 266.250 851.265 ;
    END
  END dmem_client_response_put[31]
  PIN dmem_client_response_put[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 847.265 45.450 851.265 ;
    END
  END dmem_client_response_put[3]
  PIN dmem_client_response_put[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 847.265 53.270 851.265 ;
    END
  END dmem_client_response_put[4]
  PIN dmem_client_response_put[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 847.265 61.090 851.265 ;
    END
  END dmem_client_response_put[5]
  PIN dmem_client_response_put[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 847.265 68.910 851.265 ;
    END
  END dmem_client_response_put[6]
  PIN dmem_client_response_put[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 847.265 76.730 851.265 ;
    END
  END dmem_client_response_put[7]
  PIN dmem_client_response_put[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 847.265 85.010 851.265 ;
    END
  END dmem_client_response_put[8]
  PIN dmem_client_response_put[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 847.265 92.830 851.265 ;
    END
  END dmem_client_response_put[9]
  PIN imem_client_request_get[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 847.265 554.210 851.265 ;
    END
  END imem_client_request_get[0]
  PIN imem_client_request_get[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 847.265 633.330 851.265 ;
    END
  END imem_client_request_get[10]
  PIN imem_client_request_get[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 847.265 641.150 851.265 ;
    END
  END imem_client_request_get[11]
  PIN imem_client_request_get[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 847.265 648.970 851.265 ;
    END
  END imem_client_request_get[12]
  PIN imem_client_request_get[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 847.265 656.790 851.265 ;
    END
  END imem_client_request_get[13]
  PIN imem_client_request_get[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 847.265 665.070 851.265 ;
    END
  END imem_client_request_get[14]
  PIN imem_client_request_get[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 847.265 672.890 851.265 ;
    END
  END imem_client_request_get[15]
  PIN imem_client_request_get[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 847.265 680.710 851.265 ;
    END
  END imem_client_request_get[16]
  PIN imem_client_request_get[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 847.265 688.530 851.265 ;
    END
  END imem_client_request_get[17]
  PIN imem_client_request_get[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 847.265 696.350 851.265 ;
    END
  END imem_client_request_get[18]
  PIN imem_client_request_get[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 847.265 704.170 851.265 ;
    END
  END imem_client_request_get[19]
  PIN imem_client_request_get[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 847.265 562.490 851.265 ;
    END
  END imem_client_request_get[1]
  PIN imem_client_request_get[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 847.265 711.990 851.265 ;
    END
  END imem_client_request_get[20]
  PIN imem_client_request_get[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.990 847.265 720.270 851.265 ;
    END
  END imem_client_request_get[21]
  PIN imem_client_request_get[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 847.265 728.090 851.265 ;
    END
  END imem_client_request_get[22]
  PIN imem_client_request_get[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 847.265 735.910 851.265 ;
    END
  END imem_client_request_get[23]
  PIN imem_client_request_get[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.450 847.265 743.730 851.265 ;
    END
  END imem_client_request_get[24]
  PIN imem_client_request_get[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.270 847.265 751.550 851.265 ;
    END
  END imem_client_request_get[25]
  PIN imem_client_request_get[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 847.265 759.370 851.265 ;
    END
  END imem_client_request_get[26]
  PIN imem_client_request_get[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 847.265 767.650 851.265 ;
    END
  END imem_client_request_get[27]
  PIN imem_client_request_get[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 847.265 775.470 851.265 ;
    END
  END imem_client_request_get[28]
  PIN imem_client_request_get[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.010 847.265 783.290 851.265 ;
    END
  END imem_client_request_get[29]
  PIN imem_client_request_get[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 847.265 570.310 851.265 ;
    END
  END imem_client_request_get[2]
  PIN imem_client_request_get[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.830 847.265 791.110 851.265 ;
    END
  END imem_client_request_get[30]
  PIN imem_client_request_get[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 847.265 798.930 851.265 ;
    END
  END imem_client_request_get[31]
  PIN imem_client_request_get[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 847.265 578.130 851.265 ;
    END
  END imem_client_request_get[3]
  PIN imem_client_request_get[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 847.265 585.950 851.265 ;
    END
  END imem_client_request_get[4]
  PIN imem_client_request_get[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 847.265 593.770 851.265 ;
    END
  END imem_client_request_get[5]
  PIN imem_client_request_get[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 847.265 601.590 851.265 ;
    END
  END imem_client_request_get[6]
  PIN imem_client_request_get[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 847.265 609.410 851.265 ;
    END
  END imem_client_request_get[7]
  PIN imem_client_request_get[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 847.265 617.690 851.265 ;
    END
  END imem_client_request_get[8]
  PIN imem_client_request_get[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.230 847.265 625.510 851.265 ;
    END
  END imem_client_request_get[9]
  PIN imem_client_response_put[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 847.265 558.350 851.265 ;
    END
  END imem_client_response_put[0]
  PIN imem_client_response_put[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.730 847.265 637.010 851.265 ;
    END
  END imem_client_response_put[10]
  PIN imem_client_response_put[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 847.265 645.290 851.265 ;
    END
  END imem_client_response_put[11]
  PIN imem_client_response_put[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 847.265 653.110 851.265 ;
    END
  END imem_client_response_put[12]
  PIN imem_client_response_put[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 847.265 660.930 851.265 ;
    END
  END imem_client_response_put[13]
  PIN imem_client_response_put[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.470 847.265 668.750 851.265 ;
    END
  END imem_client_response_put[14]
  PIN imem_client_response_put[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 847.265 676.570 851.265 ;
    END
  END imem_client_response_put[15]
  PIN imem_client_response_put[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 847.265 684.390 851.265 ;
    END
  END imem_client_response_put[16]
  PIN imem_client_response_put[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 847.265 692.670 851.265 ;
    END
  END imem_client_response_put[17]
  PIN imem_client_response_put[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 847.265 700.490 851.265 ;
    END
  END imem_client_response_put[18]
  PIN imem_client_response_put[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 847.265 708.310 851.265 ;
    END
  END imem_client_response_put[19]
  PIN imem_client_response_put[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 847.265 566.170 851.265 ;
    END
  END imem_client_response_put[1]
  PIN imem_client_response_put[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.850 847.265 716.130 851.265 ;
    END
  END imem_client_response_put[20]
  PIN imem_client_response_put[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.670 847.265 723.950 851.265 ;
    END
  END imem_client_response_put[21]
  PIN imem_client_response_put[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 847.265 731.770 851.265 ;
    END
  END imem_client_response_put[22]
  PIN imem_client_response_put[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 847.265 739.590 851.265 ;
    END
  END imem_client_response_put[23]
  PIN imem_client_response_put[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.590 847.265 747.870 851.265 ;
    END
  END imem_client_response_put[24]
  PIN imem_client_response_put[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.410 847.265 755.690 851.265 ;
    END
  END imem_client_response_put[25]
  PIN imem_client_response_put[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 847.265 763.510 851.265 ;
    END
  END imem_client_response_put[26]
  PIN imem_client_response_put[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.050 847.265 771.330 851.265 ;
    END
  END imem_client_response_put[27]
  PIN imem_client_response_put[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.870 847.265 779.150 851.265 ;
    END
  END imem_client_response_put[28]
  PIN imem_client_response_put[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 847.265 786.970 851.265 ;
    END
  END imem_client_response_put[29]
  PIN imem_client_response_put[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 847.265 573.990 851.265 ;
    END
  END imem_client_response_put[2]
  PIN imem_client_response_put[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.970 847.265 795.250 851.265 ;
    END
  END imem_client_response_put[30]
  PIN imem_client_response_put[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.790 847.265 803.070 851.265 ;
    END
  END imem_client_response_put[31]
  PIN imem_client_response_put[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 847.265 581.810 851.265 ;
    END
  END imem_client_response_put[3]
  PIN imem_client_response_put[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 847.265 590.090 851.265 ;
    END
  END imem_client_response_put[4]
  PIN imem_client_response_put[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 847.265 597.910 851.265 ;
    END
  END imem_client_response_put[5]
  PIN imem_client_response_put[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 847.265 605.730 851.265 ;
    END
  END imem_client_response_put[6]
  PIN imem_client_response_put[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 847.265 613.550 851.265 ;
    END
  END imem_client_response_put[7]
  PIN imem_client_response_put[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 847.265 621.370 851.265 ;
    END
  END imem_client_response_put[8]
  PIN imem_client_response_put[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 847.265 629.190 851.265 ;
    END
  END imem_client_response_put[9]
  PIN readPC[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END readPC[0]
  PIN readPC[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 824.200 840.545 824.800 ;
    END
  END readPC[10]
  PIN readPC[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 0.000 420.350 4.000 ;
    END
  END readPC[11]
  PIN readPC[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 847.265 814.570 851.265 ;
    END
  END readPC[12]
  PIN readPC[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END readPC[13]
  PIN readPC[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 831.680 840.545 832.280 ;
    END
  END readPC[14]
  PIN readPC[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END readPC[15]
  PIN readPC[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 0.000 513.730 4.000 ;
    END
  END readPC[16]
  PIN readPC[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.880 4.000 553.480 ;
    END
  END readPC[17]
  PIN readPC[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 839.160 840.545 839.760 ;
    END
  END readPC[18]
  PIN readPC[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.430 847.265 818.710 851.265 ;
    END
  END readPC[19]
  PIN readPC[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.200 4.000 127.800 ;
    END
  END readPC[1]
  PIN readPC[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.570 847.265 822.850 851.265 ;
    END
  END readPC[20]
  PIN readPC[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.250 847.265 826.530 851.265 ;
    END
  END readPC[21]
  PIN readPC[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.880 4.000 638.480 ;
    END
  END readPC[22]
  PIN readPC[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 0.000 607.110 4.000 ;
    END
  END readPC[23]
  PIN readPC[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.880 4.000 723.480 ;
    END
  END readPC[24]
  PIN readPC[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 4.000 ;
    END
  END readPC[25]
  PIN readPC[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.390 847.265 830.670 851.265 ;
    END
  END readPC[26]
  PIN readPC[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 847.265 834.350 851.265 ;
    END
  END readPC[27]
  PIN readPC[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END readPC[28]
  PIN readPC[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.210 847.265 838.490 851.265 ;
    END
  END readPC[29]
  PIN readPC[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END readPC[2]
  PIN readPC[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 846.640 840.545 847.240 ;
    END
  END readPC[30]
  PIN readPC[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.880 4.000 808.480 ;
    END
  END readPC[31]
  PIN readPC[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.470 847.265 806.750 851.265 ;
    END
  END readPC[3]
  PIN readPC[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.610 847.265 810.890 851.265 ;
    END
  END readPC[4]
  PIN readPC[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 801.760 840.545 802.360 ;
    END
  END readPC[5]
  PIN readPC[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 809.240 840.545 809.840 ;
    END
  END readPC[6]
  PIN readPC[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END readPC[7]
  PIN readPC[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END readPC[8]
  PIN readPC[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 816.720 840.545 817.320 ;
    END
  END readPC[9]
  PIN sysmem_client_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 3.440 840.545 4.040 ;
    END
  END sysmem_client_ack_i
  PIN sysmem_client_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 48.320 840.545 48.920 ;
    END
  END sysmem_client_adr_o[0]
  PIN sysmem_client_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 304.680 840.545 305.280 ;
    END
  END sysmem_client_adr_o[10]
  PIN sysmem_client_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 327.120 840.545 327.720 ;
    END
  END sysmem_client_adr_o[11]
  PIN sysmem_client_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 349.560 840.545 350.160 ;
    END
  END sysmem_client_adr_o[12]
  PIN sysmem_client_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 372.000 840.545 372.600 ;
    END
  END sysmem_client_adr_o[13]
  PIN sysmem_client_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 395.120 840.545 395.720 ;
    END
  END sysmem_client_adr_o[14]
  PIN sysmem_client_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 417.560 840.545 418.160 ;
    END
  END sysmem_client_adr_o[15]
  PIN sysmem_client_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 440.000 840.545 440.600 ;
    END
  END sysmem_client_adr_o[16]
  PIN sysmem_client_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 462.440 840.545 463.040 ;
    END
  END sysmem_client_adr_o[17]
  PIN sysmem_client_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 485.560 840.545 486.160 ;
    END
  END sysmem_client_adr_o[18]
  PIN sysmem_client_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 508.000 840.545 508.600 ;
    END
  END sysmem_client_adr_o[19]
  PIN sysmem_client_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 78.240 840.545 78.840 ;
    END
  END sysmem_client_adr_o[1]
  PIN sysmem_client_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 530.440 840.545 531.040 ;
    END
  END sysmem_client_adr_o[20]
  PIN sysmem_client_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 552.880 840.545 553.480 ;
    END
  END sysmem_client_adr_o[21]
  PIN sysmem_client_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 576.000 840.545 576.600 ;
    END
  END sysmem_client_adr_o[22]
  PIN sysmem_client_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 598.440 840.545 599.040 ;
    END
  END sysmem_client_adr_o[23]
  PIN sysmem_client_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 620.880 840.545 621.480 ;
    END
  END sysmem_client_adr_o[24]
  PIN sysmem_client_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 643.320 840.545 643.920 ;
    END
  END sysmem_client_adr_o[25]
  PIN sysmem_client_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 666.440 840.545 667.040 ;
    END
  END sysmem_client_adr_o[26]
  PIN sysmem_client_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 688.880 840.545 689.480 ;
    END
  END sysmem_client_adr_o[27]
  PIN sysmem_client_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 711.320 840.545 711.920 ;
    END
  END sysmem_client_adr_o[28]
  PIN sysmem_client_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 733.760 840.545 734.360 ;
    END
  END sysmem_client_adr_o[29]
  PIN sysmem_client_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 108.840 840.545 109.440 ;
    END
  END sysmem_client_adr_o[2]
  PIN sysmem_client_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 756.200 840.545 756.800 ;
    END
  END sysmem_client_adr_o[30]
  PIN sysmem_client_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 779.320 840.545 779.920 ;
    END
  END sysmem_client_adr_o[31]
  PIN sysmem_client_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 138.760 840.545 139.360 ;
    END
  END sysmem_client_adr_o[3]
  PIN sysmem_client_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 168.680 840.545 169.280 ;
    END
  END sysmem_client_adr_o[4]
  PIN sysmem_client_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 191.120 840.545 191.720 ;
    END
  END sysmem_client_adr_o[5]
  PIN sysmem_client_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 214.240 840.545 214.840 ;
    END
  END sysmem_client_adr_o[6]
  PIN sysmem_client_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 236.680 840.545 237.280 ;
    END
  END sysmem_client_adr_o[7]
  PIN sysmem_client_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 259.120 840.545 259.720 ;
    END
  END sysmem_client_adr_o[8]
  PIN sysmem_client_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 281.560 840.545 282.160 ;
    END
  END sysmem_client_adr_o[9]
  PIN sysmem_client_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 10.920 840.545 11.520 ;
    END
  END sysmem_client_cyc_o
  PIN sysmem_client_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 55.800 840.545 56.400 ;
    END
  END sysmem_client_dat_i[0]
  PIN sysmem_client_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 312.160 840.545 312.760 ;
    END
  END sysmem_client_dat_i[10]
  PIN sysmem_client_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 334.600 840.545 335.200 ;
    END
  END sysmem_client_dat_i[11]
  PIN sysmem_client_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 357.040 840.545 357.640 ;
    END
  END sysmem_client_dat_i[12]
  PIN sysmem_client_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 379.480 840.545 380.080 ;
    END
  END sysmem_client_dat_i[13]
  PIN sysmem_client_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 402.600 840.545 403.200 ;
    END
  END sysmem_client_dat_i[14]
  PIN sysmem_client_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 425.040 840.545 425.640 ;
    END
  END sysmem_client_dat_i[15]
  PIN sysmem_client_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 447.480 840.545 448.080 ;
    END
  END sysmem_client_dat_i[16]
  PIN sysmem_client_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 469.920 840.545 470.520 ;
    END
  END sysmem_client_dat_i[17]
  PIN sysmem_client_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 493.040 840.545 493.640 ;
    END
  END sysmem_client_dat_i[18]
  PIN sysmem_client_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 515.480 840.545 516.080 ;
    END
  END sysmem_client_dat_i[19]
  PIN sysmem_client_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 85.720 840.545 86.320 ;
    END
  END sysmem_client_dat_i[1]
  PIN sysmem_client_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 537.920 840.545 538.520 ;
    END
  END sysmem_client_dat_i[20]
  PIN sysmem_client_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 560.360 840.545 560.960 ;
    END
  END sysmem_client_dat_i[21]
  PIN sysmem_client_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 583.480 840.545 584.080 ;
    END
  END sysmem_client_dat_i[22]
  PIN sysmem_client_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 605.920 840.545 606.520 ;
    END
  END sysmem_client_dat_i[23]
  PIN sysmem_client_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 628.360 840.545 628.960 ;
    END
  END sysmem_client_dat_i[24]
  PIN sysmem_client_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 650.800 840.545 651.400 ;
    END
  END sysmem_client_dat_i[25]
  PIN sysmem_client_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 673.920 840.545 674.520 ;
    END
  END sysmem_client_dat_i[26]
  PIN sysmem_client_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 696.360 840.545 696.960 ;
    END
  END sysmem_client_dat_i[27]
  PIN sysmem_client_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 718.800 840.545 719.400 ;
    END
  END sysmem_client_dat_i[28]
  PIN sysmem_client_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 741.240 840.545 741.840 ;
    END
  END sysmem_client_dat_i[29]
  PIN sysmem_client_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 116.320 840.545 116.920 ;
    END
  END sysmem_client_dat_i[2]
  PIN sysmem_client_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 764.360 840.545 764.960 ;
    END
  END sysmem_client_dat_i[30]
  PIN sysmem_client_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 786.800 840.545 787.400 ;
    END
  END sysmem_client_dat_i[31]
  PIN sysmem_client_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 146.240 840.545 146.840 ;
    END
  END sysmem_client_dat_i[3]
  PIN sysmem_client_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 176.160 840.545 176.760 ;
    END
  END sysmem_client_dat_i[4]
  PIN sysmem_client_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 199.280 840.545 199.880 ;
    END
  END sysmem_client_dat_i[5]
  PIN sysmem_client_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 221.720 840.545 222.320 ;
    END
  END sysmem_client_dat_i[6]
  PIN sysmem_client_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 244.160 840.545 244.760 ;
    END
  END sysmem_client_dat_i[7]
  PIN sysmem_client_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 266.600 840.545 267.200 ;
    END
  END sysmem_client_dat_i[8]
  PIN sysmem_client_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 289.720 840.545 290.320 ;
    END
  END sysmem_client_dat_i[9]
  PIN sysmem_client_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 63.280 840.545 63.880 ;
    END
  END sysmem_client_dat_o[0]
  PIN sysmem_client_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 319.640 840.545 320.240 ;
    END
  END sysmem_client_dat_o[10]
  PIN sysmem_client_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 342.080 840.545 342.680 ;
    END
  END sysmem_client_dat_o[11]
  PIN sysmem_client_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 364.520 840.545 365.120 ;
    END
  END sysmem_client_dat_o[12]
  PIN sysmem_client_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 387.640 840.545 388.240 ;
    END
  END sysmem_client_dat_o[13]
  PIN sysmem_client_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 410.080 840.545 410.680 ;
    END
  END sysmem_client_dat_o[14]
  PIN sysmem_client_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 432.520 840.545 433.120 ;
    END
  END sysmem_client_dat_o[15]
  PIN sysmem_client_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 454.960 840.545 455.560 ;
    END
  END sysmem_client_dat_o[16]
  PIN sysmem_client_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 478.080 840.545 478.680 ;
    END
  END sysmem_client_dat_o[17]
  PIN sysmem_client_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 500.520 840.545 501.120 ;
    END
  END sysmem_client_dat_o[18]
  PIN sysmem_client_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 522.960 840.545 523.560 ;
    END
  END sysmem_client_dat_o[19]
  PIN sysmem_client_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 93.200 840.545 93.800 ;
    END
  END sysmem_client_dat_o[1]
  PIN sysmem_client_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 545.400 840.545 546.000 ;
    END
  END sysmem_client_dat_o[20]
  PIN sysmem_client_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 567.840 840.545 568.440 ;
    END
  END sysmem_client_dat_o[21]
  PIN sysmem_client_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 590.960 840.545 591.560 ;
    END
  END sysmem_client_dat_o[22]
  PIN sysmem_client_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 613.400 840.545 614.000 ;
    END
  END sysmem_client_dat_o[23]
  PIN sysmem_client_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 635.840 840.545 636.440 ;
    END
  END sysmem_client_dat_o[24]
  PIN sysmem_client_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 658.280 840.545 658.880 ;
    END
  END sysmem_client_dat_o[25]
  PIN sysmem_client_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 681.400 840.545 682.000 ;
    END
  END sysmem_client_dat_o[26]
  PIN sysmem_client_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 703.840 840.545 704.440 ;
    END
  END sysmem_client_dat_o[27]
  PIN sysmem_client_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 726.280 840.545 726.880 ;
    END
  END sysmem_client_dat_o[28]
  PIN sysmem_client_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 748.720 840.545 749.320 ;
    END
  END sysmem_client_dat_o[29]
  PIN sysmem_client_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 123.800 840.545 124.400 ;
    END
  END sysmem_client_dat_o[2]
  PIN sysmem_client_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 771.840 840.545 772.440 ;
    END
  END sysmem_client_dat_o[30]
  PIN sysmem_client_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 794.280 840.545 794.880 ;
    END
  END sysmem_client_dat_o[31]
  PIN sysmem_client_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 153.720 840.545 154.320 ;
    END
  END sysmem_client_dat_o[3]
  PIN sysmem_client_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 183.640 840.545 184.240 ;
    END
  END sysmem_client_dat_o[4]
  PIN sysmem_client_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 206.760 840.545 207.360 ;
    END
  END sysmem_client_dat_o[5]
  PIN sysmem_client_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 229.200 840.545 229.800 ;
    END
  END sysmem_client_dat_o[6]
  PIN sysmem_client_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 251.640 840.545 252.240 ;
    END
  END sysmem_client_dat_o[7]
  PIN sysmem_client_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 274.080 840.545 274.680 ;
    END
  END sysmem_client_dat_o[8]
  PIN sysmem_client_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 297.200 840.545 297.800 ;
    END
  END sysmem_client_dat_o[9]
  PIN sysmem_client_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 18.400 840.545 19.000 ;
    END
  END sysmem_client_err_i
  PIN sysmem_client_rty_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 25.880 840.545 26.480 ;
    END
  END sysmem_client_rty_i
  PIN sysmem_client_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 70.760 840.545 71.360 ;
    END
  END sysmem_client_sel_o[0]
  PIN sysmem_client_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 101.360 840.545 101.960 ;
    END
  END sysmem_client_sel_o[1]
  PIN sysmem_client_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 131.280 840.545 131.880 ;
    END
  END sysmem_client_sel_o[2]
  PIN sysmem_client_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 161.200 840.545 161.800 ;
    END
  END sysmem_client_sel_o[3]
  PIN sysmem_client_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 33.360 840.545 33.960 ;
    END
  END sysmem_client_stb_o
  PIN sysmem_client_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 836.545 40.840 840.545 41.440 ;
    END
  END sysmem_client_we_o
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 838.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 838.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 838.000 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 834.900 837.845 ;
      LAYER met1 ;
        RECT 0.070 10.640 840.350 841.800 ;
      LAYER met2 ;
        RECT 0.100 846.985 1.650 847.690 ;
        RECT 2.490 846.985 5.330 847.690 ;
        RECT 6.170 846.985 9.470 847.690 ;
        RECT 10.310 846.985 13.150 847.690 ;
        RECT 13.990 846.985 17.290 847.690 ;
        RECT 18.130 846.985 20.970 847.690 ;
        RECT 21.810 846.985 25.110 847.690 ;
        RECT 25.950 846.985 29.250 847.690 ;
        RECT 30.090 846.985 32.930 847.690 ;
        RECT 33.770 846.985 37.070 847.690 ;
        RECT 37.910 846.985 40.750 847.690 ;
        RECT 41.590 846.985 44.890 847.690 ;
        RECT 45.730 846.985 48.570 847.690 ;
        RECT 49.410 846.985 52.710 847.690 ;
        RECT 53.550 846.985 56.850 847.690 ;
        RECT 57.690 846.985 60.530 847.690 ;
        RECT 61.370 846.985 64.670 847.690 ;
        RECT 65.510 846.985 68.350 847.690 ;
        RECT 69.190 846.985 72.490 847.690 ;
        RECT 73.330 846.985 76.170 847.690 ;
        RECT 77.010 846.985 80.310 847.690 ;
        RECT 81.150 846.985 84.450 847.690 ;
        RECT 85.290 846.985 88.130 847.690 ;
        RECT 88.970 846.985 92.270 847.690 ;
        RECT 93.110 846.985 95.950 847.690 ;
        RECT 96.790 846.985 100.090 847.690 ;
        RECT 100.930 846.985 104.230 847.690 ;
        RECT 105.070 846.985 107.910 847.690 ;
        RECT 108.750 846.985 112.050 847.690 ;
        RECT 112.890 846.985 115.730 847.690 ;
        RECT 116.570 846.985 119.870 847.690 ;
        RECT 120.710 846.985 123.550 847.690 ;
        RECT 124.390 846.985 127.690 847.690 ;
        RECT 128.530 846.985 131.830 847.690 ;
        RECT 132.670 846.985 135.510 847.690 ;
        RECT 136.350 846.985 139.650 847.690 ;
        RECT 140.490 846.985 143.330 847.690 ;
        RECT 144.170 846.985 147.470 847.690 ;
        RECT 148.310 846.985 151.150 847.690 ;
        RECT 151.990 846.985 155.290 847.690 ;
        RECT 156.130 846.985 159.430 847.690 ;
        RECT 160.270 846.985 163.110 847.690 ;
        RECT 163.950 846.985 167.250 847.690 ;
        RECT 168.090 846.985 170.930 847.690 ;
        RECT 171.770 846.985 175.070 847.690 ;
        RECT 175.910 846.985 178.750 847.690 ;
        RECT 179.590 846.985 182.890 847.690 ;
        RECT 183.730 846.985 187.030 847.690 ;
        RECT 187.870 846.985 190.710 847.690 ;
        RECT 191.550 846.985 194.850 847.690 ;
        RECT 195.690 846.985 198.530 847.690 ;
        RECT 199.370 846.985 202.670 847.690 ;
        RECT 203.510 846.985 206.810 847.690 ;
        RECT 207.650 846.985 210.490 847.690 ;
        RECT 211.330 846.985 214.630 847.690 ;
        RECT 215.470 846.985 218.310 847.690 ;
        RECT 219.150 846.985 222.450 847.690 ;
        RECT 223.290 846.985 226.130 847.690 ;
        RECT 226.970 846.985 230.270 847.690 ;
        RECT 231.110 846.985 234.410 847.690 ;
        RECT 235.250 846.985 238.090 847.690 ;
        RECT 238.930 846.985 242.230 847.690 ;
        RECT 243.070 846.985 245.910 847.690 ;
        RECT 246.750 846.985 250.050 847.690 ;
        RECT 250.890 846.985 253.730 847.690 ;
        RECT 254.570 846.985 257.870 847.690 ;
        RECT 258.710 846.985 262.010 847.690 ;
        RECT 262.850 846.985 265.690 847.690 ;
        RECT 266.530 846.985 269.830 847.690 ;
        RECT 270.670 846.985 273.510 847.690 ;
        RECT 274.350 846.985 277.650 847.690 ;
        RECT 278.490 846.985 281.790 847.690 ;
        RECT 282.630 846.985 285.470 847.690 ;
        RECT 286.310 846.985 289.610 847.690 ;
        RECT 290.450 846.985 293.290 847.690 ;
        RECT 294.130 846.985 297.430 847.690 ;
        RECT 298.270 846.985 301.110 847.690 ;
        RECT 301.950 846.985 305.250 847.690 ;
        RECT 306.090 846.985 309.390 847.690 ;
        RECT 310.230 846.985 313.070 847.690 ;
        RECT 313.910 846.985 317.210 847.690 ;
        RECT 318.050 846.985 320.890 847.690 ;
        RECT 321.730 846.985 325.030 847.690 ;
        RECT 325.870 846.985 328.710 847.690 ;
        RECT 329.550 846.985 332.850 847.690 ;
        RECT 333.690 846.985 336.990 847.690 ;
        RECT 337.830 846.985 340.670 847.690 ;
        RECT 341.510 846.985 344.810 847.690 ;
        RECT 345.650 846.985 348.490 847.690 ;
        RECT 349.330 846.985 352.630 847.690 ;
        RECT 353.470 846.985 356.310 847.690 ;
        RECT 357.150 846.985 360.450 847.690 ;
        RECT 361.290 846.985 364.590 847.690 ;
        RECT 365.430 846.985 368.270 847.690 ;
        RECT 369.110 846.985 372.410 847.690 ;
        RECT 373.250 846.985 376.090 847.690 ;
        RECT 376.930 846.985 380.230 847.690 ;
        RECT 381.070 846.985 384.370 847.690 ;
        RECT 385.210 846.985 388.050 847.690 ;
        RECT 388.890 846.985 392.190 847.690 ;
        RECT 393.030 846.985 395.870 847.690 ;
        RECT 396.710 846.985 400.010 847.690 ;
        RECT 400.850 846.985 403.690 847.690 ;
        RECT 404.530 846.985 407.830 847.690 ;
        RECT 408.670 846.985 411.970 847.690 ;
        RECT 412.810 846.985 415.650 847.690 ;
        RECT 416.490 846.985 419.790 847.690 ;
        RECT 420.630 846.985 423.470 847.690 ;
        RECT 424.310 846.985 427.610 847.690 ;
        RECT 428.450 846.985 431.290 847.690 ;
        RECT 432.130 846.985 435.430 847.690 ;
        RECT 436.270 846.985 439.570 847.690 ;
        RECT 440.410 846.985 443.250 847.690 ;
        RECT 444.090 846.985 447.390 847.690 ;
        RECT 448.230 846.985 451.070 847.690 ;
        RECT 451.910 846.985 455.210 847.690 ;
        RECT 456.050 846.985 458.890 847.690 ;
        RECT 459.730 846.985 463.030 847.690 ;
        RECT 463.870 846.985 467.170 847.690 ;
        RECT 468.010 846.985 470.850 847.690 ;
        RECT 471.690 846.985 474.990 847.690 ;
        RECT 475.830 846.985 478.670 847.690 ;
        RECT 479.510 846.985 482.810 847.690 ;
        RECT 483.650 846.985 486.950 847.690 ;
        RECT 487.790 846.985 490.630 847.690 ;
        RECT 491.470 846.985 494.770 847.690 ;
        RECT 495.610 846.985 498.450 847.690 ;
        RECT 499.290 846.985 502.590 847.690 ;
        RECT 503.430 846.985 506.270 847.690 ;
        RECT 507.110 846.985 510.410 847.690 ;
        RECT 511.250 846.985 514.550 847.690 ;
        RECT 515.390 846.985 518.230 847.690 ;
        RECT 519.070 846.985 522.370 847.690 ;
        RECT 523.210 846.985 526.050 847.690 ;
        RECT 526.890 846.985 530.190 847.690 ;
        RECT 531.030 846.985 533.870 847.690 ;
        RECT 534.710 846.985 538.010 847.690 ;
        RECT 538.850 846.985 542.150 847.690 ;
        RECT 542.990 846.985 545.830 847.690 ;
        RECT 546.670 846.985 549.970 847.690 ;
        RECT 550.810 846.985 553.650 847.690 ;
        RECT 554.490 846.985 557.790 847.690 ;
        RECT 558.630 846.985 561.930 847.690 ;
        RECT 562.770 846.985 565.610 847.690 ;
        RECT 566.450 846.985 569.750 847.690 ;
        RECT 570.590 846.985 573.430 847.690 ;
        RECT 574.270 846.985 577.570 847.690 ;
        RECT 578.410 846.985 581.250 847.690 ;
        RECT 582.090 846.985 585.390 847.690 ;
        RECT 586.230 846.985 589.530 847.690 ;
        RECT 590.370 846.985 593.210 847.690 ;
        RECT 594.050 846.985 597.350 847.690 ;
        RECT 598.190 846.985 601.030 847.690 ;
        RECT 601.870 846.985 605.170 847.690 ;
        RECT 606.010 846.985 608.850 847.690 ;
        RECT 609.690 846.985 612.990 847.690 ;
        RECT 613.830 846.985 617.130 847.690 ;
        RECT 617.970 846.985 620.810 847.690 ;
        RECT 621.650 846.985 624.950 847.690 ;
        RECT 625.790 846.985 628.630 847.690 ;
        RECT 629.470 846.985 632.770 847.690 ;
        RECT 633.610 846.985 636.450 847.690 ;
        RECT 637.290 846.985 640.590 847.690 ;
        RECT 641.430 846.985 644.730 847.690 ;
        RECT 645.570 846.985 648.410 847.690 ;
        RECT 649.250 846.985 652.550 847.690 ;
        RECT 653.390 846.985 656.230 847.690 ;
        RECT 657.070 846.985 660.370 847.690 ;
        RECT 661.210 846.985 664.510 847.690 ;
        RECT 665.350 846.985 668.190 847.690 ;
        RECT 669.030 846.985 672.330 847.690 ;
        RECT 673.170 846.985 676.010 847.690 ;
        RECT 676.850 846.985 680.150 847.690 ;
        RECT 680.990 846.985 683.830 847.690 ;
        RECT 684.670 846.985 687.970 847.690 ;
        RECT 688.810 846.985 692.110 847.690 ;
        RECT 692.950 846.985 695.790 847.690 ;
        RECT 696.630 846.985 699.930 847.690 ;
        RECT 700.770 846.985 703.610 847.690 ;
        RECT 704.450 846.985 707.750 847.690 ;
        RECT 708.590 846.985 711.430 847.690 ;
        RECT 712.270 846.985 715.570 847.690 ;
        RECT 716.410 846.985 719.710 847.690 ;
        RECT 720.550 846.985 723.390 847.690 ;
        RECT 724.230 846.985 727.530 847.690 ;
        RECT 728.370 846.985 731.210 847.690 ;
        RECT 732.050 846.985 735.350 847.690 ;
        RECT 736.190 846.985 739.030 847.690 ;
        RECT 739.870 846.985 743.170 847.690 ;
        RECT 744.010 846.985 747.310 847.690 ;
        RECT 748.150 846.985 750.990 847.690 ;
        RECT 751.830 846.985 755.130 847.690 ;
        RECT 755.970 846.985 758.810 847.690 ;
        RECT 759.650 846.985 762.950 847.690 ;
        RECT 763.790 846.985 767.090 847.690 ;
        RECT 767.930 846.985 770.770 847.690 ;
        RECT 771.610 846.985 774.910 847.690 ;
        RECT 775.750 846.985 778.590 847.690 ;
        RECT 779.430 846.985 782.730 847.690 ;
        RECT 783.570 846.985 786.410 847.690 ;
        RECT 787.250 846.985 790.550 847.690 ;
        RECT 791.390 846.985 794.690 847.690 ;
        RECT 795.530 846.985 798.370 847.690 ;
        RECT 799.210 846.985 802.510 847.690 ;
        RECT 803.350 846.985 806.190 847.690 ;
        RECT 807.030 846.985 810.330 847.690 ;
        RECT 811.170 846.985 814.010 847.690 ;
        RECT 814.850 846.985 818.150 847.690 ;
        RECT 818.990 846.985 822.290 847.690 ;
        RECT 823.130 846.985 825.970 847.690 ;
        RECT 826.810 846.985 830.110 847.690 ;
        RECT 830.950 846.985 833.790 847.690 ;
        RECT 834.630 846.985 837.930 847.690 ;
        RECT 838.770 846.985 840.320 847.690 ;
        RECT 0.100 4.280 840.320 846.985 ;
        RECT 0.100 3.555 46.270 4.280 ;
        RECT 47.110 3.555 139.650 4.280 ;
        RECT 140.490 3.555 233.030 4.280 ;
        RECT 233.870 3.555 326.410 4.280 ;
        RECT 327.250 3.555 419.790 4.280 ;
        RECT 420.630 3.555 513.170 4.280 ;
        RECT 514.010 3.555 606.550 4.280 ;
        RECT 607.390 3.555 699.930 4.280 ;
        RECT 700.770 3.555 793.310 4.280 ;
        RECT 794.150 3.555 840.320 4.280 ;
      LAYER met3 ;
        RECT 4.000 846.240 836.145 847.105 ;
        RECT 4.000 840.160 836.890 846.240 ;
        RECT 4.000 838.760 836.145 840.160 ;
        RECT 4.000 832.680 836.890 838.760 ;
        RECT 4.000 831.280 836.145 832.680 ;
        RECT 4.000 825.200 836.890 831.280 ;
        RECT 4.000 823.800 836.145 825.200 ;
        RECT 4.000 817.720 836.890 823.800 ;
        RECT 4.000 816.320 836.145 817.720 ;
        RECT 4.000 810.240 836.890 816.320 ;
        RECT 4.000 808.880 836.145 810.240 ;
        RECT 4.400 808.840 836.145 808.880 ;
        RECT 4.400 807.480 836.890 808.840 ;
        RECT 4.000 802.760 836.890 807.480 ;
        RECT 4.000 801.360 836.145 802.760 ;
        RECT 4.000 795.280 836.890 801.360 ;
        RECT 4.000 793.880 836.145 795.280 ;
        RECT 4.000 787.800 836.890 793.880 ;
        RECT 4.000 786.400 836.145 787.800 ;
        RECT 4.000 780.320 836.890 786.400 ;
        RECT 4.000 778.920 836.145 780.320 ;
        RECT 4.000 772.840 836.890 778.920 ;
        RECT 4.000 771.440 836.145 772.840 ;
        RECT 4.000 765.360 836.890 771.440 ;
        RECT 4.000 763.960 836.145 765.360 ;
        RECT 4.000 757.200 836.890 763.960 ;
        RECT 4.000 755.800 836.145 757.200 ;
        RECT 4.000 749.720 836.890 755.800 ;
        RECT 4.000 748.320 836.145 749.720 ;
        RECT 4.000 742.240 836.890 748.320 ;
        RECT 4.000 740.840 836.145 742.240 ;
        RECT 4.000 734.760 836.890 740.840 ;
        RECT 4.000 733.360 836.145 734.760 ;
        RECT 4.000 727.280 836.890 733.360 ;
        RECT 4.000 725.880 836.145 727.280 ;
        RECT 4.000 723.880 836.890 725.880 ;
        RECT 4.400 722.480 836.890 723.880 ;
        RECT 4.000 719.800 836.890 722.480 ;
        RECT 4.000 718.400 836.145 719.800 ;
        RECT 4.000 712.320 836.890 718.400 ;
        RECT 4.000 710.920 836.145 712.320 ;
        RECT 4.000 704.840 836.890 710.920 ;
        RECT 4.000 703.440 836.145 704.840 ;
        RECT 4.000 697.360 836.890 703.440 ;
        RECT 4.000 695.960 836.145 697.360 ;
        RECT 4.000 689.880 836.890 695.960 ;
        RECT 4.000 688.480 836.145 689.880 ;
        RECT 4.000 682.400 836.890 688.480 ;
        RECT 4.000 681.000 836.145 682.400 ;
        RECT 4.000 674.920 836.890 681.000 ;
        RECT 4.000 673.520 836.145 674.920 ;
        RECT 4.000 667.440 836.890 673.520 ;
        RECT 4.000 666.040 836.145 667.440 ;
        RECT 4.000 659.280 836.890 666.040 ;
        RECT 4.000 657.880 836.145 659.280 ;
        RECT 4.000 651.800 836.890 657.880 ;
        RECT 4.000 650.400 836.145 651.800 ;
        RECT 4.000 644.320 836.890 650.400 ;
        RECT 4.000 642.920 836.145 644.320 ;
        RECT 4.000 638.880 836.890 642.920 ;
        RECT 4.400 637.480 836.890 638.880 ;
        RECT 4.000 636.840 836.890 637.480 ;
        RECT 4.000 635.440 836.145 636.840 ;
        RECT 4.000 629.360 836.890 635.440 ;
        RECT 4.000 627.960 836.145 629.360 ;
        RECT 4.000 621.880 836.890 627.960 ;
        RECT 4.000 620.480 836.145 621.880 ;
        RECT 4.000 614.400 836.890 620.480 ;
        RECT 4.000 613.000 836.145 614.400 ;
        RECT 4.000 606.920 836.890 613.000 ;
        RECT 4.000 605.520 836.145 606.920 ;
        RECT 4.000 599.440 836.890 605.520 ;
        RECT 4.000 598.040 836.145 599.440 ;
        RECT 4.000 591.960 836.890 598.040 ;
        RECT 4.000 590.560 836.145 591.960 ;
        RECT 4.000 584.480 836.890 590.560 ;
        RECT 4.000 583.080 836.145 584.480 ;
        RECT 4.000 577.000 836.890 583.080 ;
        RECT 4.000 575.600 836.145 577.000 ;
        RECT 4.000 568.840 836.890 575.600 ;
        RECT 4.000 567.440 836.145 568.840 ;
        RECT 4.000 561.360 836.890 567.440 ;
        RECT 4.000 559.960 836.145 561.360 ;
        RECT 4.000 553.880 836.890 559.960 ;
        RECT 4.400 552.480 836.145 553.880 ;
        RECT 4.000 546.400 836.890 552.480 ;
        RECT 4.000 545.000 836.145 546.400 ;
        RECT 4.000 538.920 836.890 545.000 ;
        RECT 4.000 537.520 836.145 538.920 ;
        RECT 4.000 531.440 836.890 537.520 ;
        RECT 4.000 530.040 836.145 531.440 ;
        RECT 4.000 523.960 836.890 530.040 ;
        RECT 4.000 522.560 836.145 523.960 ;
        RECT 4.000 516.480 836.890 522.560 ;
        RECT 4.000 515.080 836.145 516.480 ;
        RECT 4.000 509.000 836.890 515.080 ;
        RECT 4.000 507.600 836.145 509.000 ;
        RECT 4.000 501.520 836.890 507.600 ;
        RECT 4.000 500.120 836.145 501.520 ;
        RECT 4.000 494.040 836.890 500.120 ;
        RECT 4.000 492.640 836.145 494.040 ;
        RECT 4.000 486.560 836.890 492.640 ;
        RECT 4.000 485.160 836.145 486.560 ;
        RECT 4.000 479.080 836.890 485.160 ;
        RECT 4.000 477.680 836.145 479.080 ;
        RECT 4.000 470.920 836.890 477.680 ;
        RECT 4.000 469.520 836.145 470.920 ;
        RECT 4.000 468.880 836.890 469.520 ;
        RECT 4.400 467.480 836.890 468.880 ;
        RECT 4.000 463.440 836.890 467.480 ;
        RECT 4.000 462.040 836.145 463.440 ;
        RECT 4.000 455.960 836.890 462.040 ;
        RECT 4.000 454.560 836.145 455.960 ;
        RECT 4.000 448.480 836.890 454.560 ;
        RECT 4.000 447.080 836.145 448.480 ;
        RECT 4.000 441.000 836.890 447.080 ;
        RECT 4.000 439.600 836.145 441.000 ;
        RECT 4.000 433.520 836.890 439.600 ;
        RECT 4.000 432.120 836.145 433.520 ;
        RECT 4.000 426.040 836.890 432.120 ;
        RECT 4.000 424.640 836.145 426.040 ;
        RECT 4.000 418.560 836.890 424.640 ;
        RECT 4.000 417.160 836.145 418.560 ;
        RECT 4.000 411.080 836.890 417.160 ;
        RECT 4.000 409.680 836.145 411.080 ;
        RECT 4.000 403.600 836.890 409.680 ;
        RECT 4.000 402.200 836.145 403.600 ;
        RECT 4.000 396.120 836.890 402.200 ;
        RECT 4.000 394.720 836.145 396.120 ;
        RECT 4.000 388.640 836.890 394.720 ;
        RECT 4.000 387.240 836.145 388.640 ;
        RECT 4.000 383.200 836.890 387.240 ;
        RECT 4.400 381.800 836.890 383.200 ;
        RECT 4.000 380.480 836.890 381.800 ;
        RECT 4.000 379.080 836.145 380.480 ;
        RECT 4.000 373.000 836.890 379.080 ;
        RECT 4.000 371.600 836.145 373.000 ;
        RECT 4.000 365.520 836.890 371.600 ;
        RECT 4.000 364.120 836.145 365.520 ;
        RECT 4.000 358.040 836.890 364.120 ;
        RECT 4.000 356.640 836.145 358.040 ;
        RECT 4.000 350.560 836.890 356.640 ;
        RECT 4.000 349.160 836.145 350.560 ;
        RECT 4.000 343.080 836.890 349.160 ;
        RECT 4.000 341.680 836.145 343.080 ;
        RECT 4.000 335.600 836.890 341.680 ;
        RECT 4.000 334.200 836.145 335.600 ;
        RECT 4.000 328.120 836.890 334.200 ;
        RECT 4.000 326.720 836.145 328.120 ;
        RECT 4.000 320.640 836.890 326.720 ;
        RECT 4.000 319.240 836.145 320.640 ;
        RECT 4.000 313.160 836.890 319.240 ;
        RECT 4.000 311.760 836.145 313.160 ;
        RECT 4.000 305.680 836.890 311.760 ;
        RECT 4.000 304.280 836.145 305.680 ;
        RECT 4.000 298.200 836.890 304.280 ;
        RECT 4.400 296.800 836.145 298.200 ;
        RECT 4.000 290.720 836.890 296.800 ;
        RECT 4.000 289.320 836.145 290.720 ;
        RECT 4.000 282.560 836.890 289.320 ;
        RECT 4.000 281.160 836.145 282.560 ;
        RECT 4.000 275.080 836.890 281.160 ;
        RECT 4.000 273.680 836.145 275.080 ;
        RECT 4.000 267.600 836.890 273.680 ;
        RECT 4.000 266.200 836.145 267.600 ;
        RECT 4.000 260.120 836.890 266.200 ;
        RECT 4.000 258.720 836.145 260.120 ;
        RECT 4.000 252.640 836.890 258.720 ;
        RECT 4.000 251.240 836.145 252.640 ;
        RECT 4.000 245.160 836.890 251.240 ;
        RECT 4.000 243.760 836.145 245.160 ;
        RECT 4.000 237.680 836.890 243.760 ;
        RECT 4.000 236.280 836.145 237.680 ;
        RECT 4.000 230.200 836.890 236.280 ;
        RECT 4.000 228.800 836.145 230.200 ;
        RECT 4.000 222.720 836.890 228.800 ;
        RECT 4.000 221.320 836.145 222.720 ;
        RECT 4.000 215.240 836.890 221.320 ;
        RECT 4.000 213.840 836.145 215.240 ;
        RECT 4.000 213.200 836.890 213.840 ;
        RECT 4.400 211.800 836.890 213.200 ;
        RECT 4.000 207.760 836.890 211.800 ;
        RECT 4.000 206.360 836.145 207.760 ;
        RECT 4.000 200.280 836.890 206.360 ;
        RECT 4.000 198.880 836.145 200.280 ;
        RECT 4.000 192.120 836.890 198.880 ;
        RECT 4.000 190.720 836.145 192.120 ;
        RECT 4.000 184.640 836.890 190.720 ;
        RECT 4.000 183.240 836.145 184.640 ;
        RECT 4.000 177.160 836.890 183.240 ;
        RECT 4.000 175.760 836.145 177.160 ;
        RECT 4.000 169.680 836.890 175.760 ;
        RECT 4.000 168.280 836.145 169.680 ;
        RECT 4.000 162.200 836.890 168.280 ;
        RECT 4.000 160.800 836.145 162.200 ;
        RECT 4.000 154.720 836.890 160.800 ;
        RECT 4.000 153.320 836.145 154.720 ;
        RECT 4.000 147.240 836.890 153.320 ;
        RECT 4.000 145.840 836.145 147.240 ;
        RECT 4.000 139.760 836.890 145.840 ;
        RECT 4.000 138.360 836.145 139.760 ;
        RECT 4.000 132.280 836.890 138.360 ;
        RECT 4.000 130.880 836.145 132.280 ;
        RECT 4.000 128.200 836.890 130.880 ;
        RECT 4.400 126.800 836.890 128.200 ;
        RECT 4.000 124.800 836.890 126.800 ;
        RECT 4.000 123.400 836.145 124.800 ;
        RECT 4.000 117.320 836.890 123.400 ;
        RECT 4.000 115.920 836.145 117.320 ;
        RECT 4.000 109.840 836.890 115.920 ;
        RECT 4.000 108.440 836.145 109.840 ;
        RECT 4.000 102.360 836.890 108.440 ;
        RECT 4.000 100.960 836.145 102.360 ;
        RECT 4.000 94.200 836.890 100.960 ;
        RECT 4.000 92.800 836.145 94.200 ;
        RECT 4.000 86.720 836.890 92.800 ;
        RECT 4.000 85.320 836.145 86.720 ;
        RECT 4.000 79.240 836.890 85.320 ;
        RECT 4.000 77.840 836.145 79.240 ;
        RECT 4.000 71.760 836.890 77.840 ;
        RECT 4.000 70.360 836.145 71.760 ;
        RECT 4.000 64.280 836.890 70.360 ;
        RECT 4.000 62.880 836.145 64.280 ;
        RECT 4.000 56.800 836.890 62.880 ;
        RECT 4.000 55.400 836.145 56.800 ;
        RECT 4.000 49.320 836.890 55.400 ;
        RECT 4.000 47.920 836.145 49.320 ;
        RECT 4.000 43.200 836.890 47.920 ;
        RECT 4.400 41.840 836.890 43.200 ;
        RECT 4.400 41.800 836.145 41.840 ;
        RECT 4.000 40.440 836.145 41.800 ;
        RECT 4.000 34.360 836.890 40.440 ;
        RECT 4.000 32.960 836.145 34.360 ;
        RECT 4.000 26.880 836.890 32.960 ;
        RECT 4.000 25.480 836.145 26.880 ;
        RECT 4.000 19.400 836.890 25.480 ;
        RECT 4.000 18.000 836.145 19.400 ;
        RECT 4.000 11.920 836.890 18.000 ;
        RECT 4.000 10.520 836.145 11.920 ;
        RECT 4.000 4.440 836.890 10.520 ;
        RECT 4.000 3.575 836.145 4.440 ;
      LAYER met4 ;
        RECT 23.295 16.495 97.440 828.745 ;
        RECT 99.840 16.495 174.240 828.745 ;
        RECT 176.640 16.495 251.040 828.745 ;
        RECT 253.440 16.495 327.840 828.745 ;
        RECT 330.240 16.495 404.640 828.745 ;
        RECT 407.040 16.495 481.440 828.745 ;
        RECT 483.840 16.495 558.240 828.745 ;
        RECT 560.640 16.495 635.040 828.745 ;
        RECT 637.440 16.495 711.840 828.745 ;
        RECT 714.240 16.495 788.640 828.745 ;
        RECT 791.040 16.495 827.705 828.745 ;
  END
END mkLanaiCPU
END LIBRARY

