magic
tech sky130A
magscale 1 2
timestamp 1647708161
<< obsli1 >>
rect 1104 2159 166796 167569
<< obsm1 >>
rect 14 2128 167610 168224
<< metal2 >>
rect 386 169318 442 170118
rect 1122 169318 1178 170118
rect 1950 169318 2006 170118
rect 2778 169318 2834 170118
rect 3514 169318 3570 170118
rect 4342 169318 4398 170118
rect 5170 169318 5226 170118
rect 5906 169318 5962 170118
rect 6734 169318 6790 170118
rect 7562 169318 7618 170118
rect 8298 169318 8354 170118
rect 9126 169318 9182 170118
rect 9954 169318 10010 170118
rect 10782 169318 10838 170118
rect 11518 169318 11574 170118
rect 12346 169318 12402 170118
rect 13174 169318 13230 170118
rect 13910 169318 13966 170118
rect 14738 169318 14794 170118
rect 15566 169318 15622 170118
rect 16302 169318 16358 170118
rect 17130 169318 17186 170118
rect 17958 169318 18014 170118
rect 18694 169318 18750 170118
rect 19522 169318 19578 170118
rect 20350 169318 20406 170118
rect 21178 169318 21234 170118
rect 21914 169318 21970 170118
rect 22742 169318 22798 170118
rect 23570 169318 23626 170118
rect 24306 169318 24362 170118
rect 25134 169318 25190 170118
rect 25962 169318 26018 170118
rect 26698 169318 26754 170118
rect 27526 169318 27582 170118
rect 28354 169318 28410 170118
rect 29182 169318 29238 170118
rect 29918 169318 29974 170118
rect 30746 169318 30802 170118
rect 31574 169318 31630 170118
rect 32310 169318 32366 170118
rect 33138 169318 33194 170118
rect 33966 169318 34022 170118
rect 34702 169318 34758 170118
rect 35530 169318 35586 170118
rect 36358 169318 36414 170118
rect 37094 169318 37150 170118
rect 37922 169318 37978 170118
rect 38750 169318 38806 170118
rect 39578 169318 39634 170118
rect 40314 169318 40370 170118
rect 41142 169318 41198 170118
rect 41970 169318 42026 170118
rect 42706 169318 42762 170118
rect 43534 169318 43590 170118
rect 44362 169318 44418 170118
rect 45098 169318 45154 170118
rect 45926 169318 45982 170118
rect 46754 169318 46810 170118
rect 47582 169318 47638 170118
rect 48318 169318 48374 170118
rect 49146 169318 49202 170118
rect 49974 169318 50030 170118
rect 50710 169318 50766 170118
rect 51538 169318 51594 170118
rect 52366 169318 52422 170118
rect 53102 169318 53158 170118
rect 53930 169318 53986 170118
rect 54758 169318 54814 170118
rect 55494 169318 55550 170118
rect 56322 169318 56378 170118
rect 57150 169318 57206 170118
rect 57978 169318 58034 170118
rect 58714 169318 58770 170118
rect 59542 169318 59598 170118
rect 60370 169318 60426 170118
rect 61106 169318 61162 170118
rect 61934 169318 61990 170118
rect 62762 169318 62818 170118
rect 63498 169318 63554 170118
rect 64326 169318 64382 170118
rect 65154 169318 65210 170118
rect 65982 169318 66038 170118
rect 66718 169318 66774 170118
rect 67546 169318 67602 170118
rect 68374 169318 68430 170118
rect 69110 169318 69166 170118
rect 69938 169318 69994 170118
rect 70766 169318 70822 170118
rect 71502 169318 71558 170118
rect 72330 169318 72386 170118
rect 73158 169318 73214 170118
rect 73894 169318 73950 170118
rect 74722 169318 74778 170118
rect 75550 169318 75606 170118
rect 76378 169318 76434 170118
rect 77114 169318 77170 170118
rect 77942 169318 77998 170118
rect 78770 169318 78826 170118
rect 79506 169318 79562 170118
rect 80334 169318 80390 170118
rect 81162 169318 81218 170118
rect 81898 169318 81954 170118
rect 82726 169318 82782 170118
rect 83554 169318 83610 170118
rect 84382 169318 84438 170118
rect 85118 169318 85174 170118
rect 85946 169318 86002 170118
rect 86774 169318 86830 170118
rect 87510 169318 87566 170118
rect 88338 169318 88394 170118
rect 89166 169318 89222 170118
rect 89902 169318 89958 170118
rect 90730 169318 90786 170118
rect 91558 169318 91614 170118
rect 92294 169318 92350 170118
rect 93122 169318 93178 170118
rect 93950 169318 94006 170118
rect 94778 169318 94834 170118
rect 95514 169318 95570 170118
rect 96342 169318 96398 170118
rect 97170 169318 97226 170118
rect 97906 169318 97962 170118
rect 98734 169318 98790 170118
rect 99562 169318 99618 170118
rect 100298 169318 100354 170118
rect 101126 169318 101182 170118
rect 101954 169318 102010 170118
rect 102690 169318 102746 170118
rect 103518 169318 103574 170118
rect 104346 169318 104402 170118
rect 105174 169318 105230 170118
rect 105910 169318 105966 170118
rect 106738 169318 106794 170118
rect 107566 169318 107622 170118
rect 108302 169318 108358 170118
rect 109130 169318 109186 170118
rect 109958 169318 110014 170118
rect 110694 169318 110750 170118
rect 111522 169318 111578 170118
rect 112350 169318 112406 170118
rect 113178 169318 113234 170118
rect 113914 169318 113970 170118
rect 114742 169318 114798 170118
rect 115570 169318 115626 170118
rect 116306 169318 116362 170118
rect 117134 169318 117190 170118
rect 117962 169318 118018 170118
rect 118698 169318 118754 170118
rect 119526 169318 119582 170118
rect 120354 169318 120410 170118
rect 121090 169318 121146 170118
rect 121918 169318 121974 170118
rect 122746 169318 122802 170118
rect 123574 169318 123630 170118
rect 124310 169318 124366 170118
rect 125138 169318 125194 170118
rect 125966 169318 126022 170118
rect 126702 169318 126758 170118
rect 127530 169318 127586 170118
rect 128358 169318 128414 170118
rect 129094 169318 129150 170118
rect 129922 169318 129978 170118
rect 130750 169318 130806 170118
rect 131578 169318 131634 170118
rect 132314 169318 132370 170118
rect 133142 169318 133198 170118
rect 133970 169318 134026 170118
rect 134706 169318 134762 170118
rect 135534 169318 135590 170118
rect 136362 169318 136418 170118
rect 137098 169318 137154 170118
rect 137926 169318 137982 170118
rect 138754 169318 138810 170118
rect 139490 169318 139546 170118
rect 140318 169318 140374 170118
rect 141146 169318 141202 170118
rect 141974 169318 142030 170118
rect 142710 169318 142766 170118
rect 143538 169318 143594 170118
rect 144366 169318 144422 170118
rect 145102 169318 145158 170118
rect 145930 169318 145986 170118
rect 146758 169318 146814 170118
rect 147494 169318 147550 170118
rect 148322 169318 148378 170118
rect 149150 169318 149206 170118
rect 149978 169318 150034 170118
rect 150714 169318 150770 170118
rect 151542 169318 151598 170118
rect 152370 169318 152426 170118
rect 153106 169318 153162 170118
rect 153934 169318 153990 170118
rect 154762 169318 154818 170118
rect 155498 169318 155554 170118
rect 156326 169318 156382 170118
rect 157154 169318 157210 170118
rect 157890 169318 157946 170118
rect 158718 169318 158774 170118
rect 159546 169318 159602 170118
rect 160374 169318 160430 170118
rect 161110 169318 161166 170118
rect 161938 169318 161994 170118
rect 162766 169318 162822 170118
rect 163502 169318 163558 170118
rect 164330 169318 164386 170118
rect 165158 169318 165214 170118
rect 165894 169318 165950 170118
rect 166722 169318 166778 170118
rect 167550 169318 167606 170118
rect 16762 0 16818 800
rect 50342 0 50398 800
rect 83922 0 83978 800
rect 117502 0 117558 800
rect 151082 0 151138 800
<< obsm2 >>
rect 20 169262 330 169402
rect 498 169262 1066 169402
rect 1234 169262 1894 169402
rect 2062 169262 2722 169402
rect 2890 169262 3458 169402
rect 3626 169262 4286 169402
rect 4454 169262 5114 169402
rect 5282 169262 5850 169402
rect 6018 169262 6678 169402
rect 6846 169262 7506 169402
rect 7674 169262 8242 169402
rect 8410 169262 9070 169402
rect 9238 169262 9898 169402
rect 10066 169262 10726 169402
rect 10894 169262 11462 169402
rect 11630 169262 12290 169402
rect 12458 169262 13118 169402
rect 13286 169262 13854 169402
rect 14022 169262 14682 169402
rect 14850 169262 15510 169402
rect 15678 169262 16246 169402
rect 16414 169262 17074 169402
rect 17242 169262 17902 169402
rect 18070 169262 18638 169402
rect 18806 169262 19466 169402
rect 19634 169262 20294 169402
rect 20462 169262 21122 169402
rect 21290 169262 21858 169402
rect 22026 169262 22686 169402
rect 22854 169262 23514 169402
rect 23682 169262 24250 169402
rect 24418 169262 25078 169402
rect 25246 169262 25906 169402
rect 26074 169262 26642 169402
rect 26810 169262 27470 169402
rect 27638 169262 28298 169402
rect 28466 169262 29126 169402
rect 29294 169262 29862 169402
rect 30030 169262 30690 169402
rect 30858 169262 31518 169402
rect 31686 169262 32254 169402
rect 32422 169262 33082 169402
rect 33250 169262 33910 169402
rect 34078 169262 34646 169402
rect 34814 169262 35474 169402
rect 35642 169262 36302 169402
rect 36470 169262 37038 169402
rect 37206 169262 37866 169402
rect 38034 169262 38694 169402
rect 38862 169262 39522 169402
rect 39690 169262 40258 169402
rect 40426 169262 41086 169402
rect 41254 169262 41914 169402
rect 42082 169262 42650 169402
rect 42818 169262 43478 169402
rect 43646 169262 44306 169402
rect 44474 169262 45042 169402
rect 45210 169262 45870 169402
rect 46038 169262 46698 169402
rect 46866 169262 47526 169402
rect 47694 169262 48262 169402
rect 48430 169262 49090 169402
rect 49258 169262 49918 169402
rect 50086 169262 50654 169402
rect 50822 169262 51482 169402
rect 51650 169262 52310 169402
rect 52478 169262 53046 169402
rect 53214 169262 53874 169402
rect 54042 169262 54702 169402
rect 54870 169262 55438 169402
rect 55606 169262 56266 169402
rect 56434 169262 57094 169402
rect 57262 169262 57922 169402
rect 58090 169262 58658 169402
rect 58826 169262 59486 169402
rect 59654 169262 60314 169402
rect 60482 169262 61050 169402
rect 61218 169262 61878 169402
rect 62046 169262 62706 169402
rect 62874 169262 63442 169402
rect 63610 169262 64270 169402
rect 64438 169262 65098 169402
rect 65266 169262 65926 169402
rect 66094 169262 66662 169402
rect 66830 169262 67490 169402
rect 67658 169262 68318 169402
rect 68486 169262 69054 169402
rect 69222 169262 69882 169402
rect 70050 169262 70710 169402
rect 70878 169262 71446 169402
rect 71614 169262 72274 169402
rect 72442 169262 73102 169402
rect 73270 169262 73838 169402
rect 74006 169262 74666 169402
rect 74834 169262 75494 169402
rect 75662 169262 76322 169402
rect 76490 169262 77058 169402
rect 77226 169262 77886 169402
rect 78054 169262 78714 169402
rect 78882 169262 79450 169402
rect 79618 169262 80278 169402
rect 80446 169262 81106 169402
rect 81274 169262 81842 169402
rect 82010 169262 82670 169402
rect 82838 169262 83498 169402
rect 83666 169262 84326 169402
rect 84494 169262 85062 169402
rect 85230 169262 85890 169402
rect 86058 169262 86718 169402
rect 86886 169262 87454 169402
rect 87622 169262 88282 169402
rect 88450 169262 89110 169402
rect 89278 169262 89846 169402
rect 90014 169262 90674 169402
rect 90842 169262 91502 169402
rect 91670 169262 92238 169402
rect 92406 169262 93066 169402
rect 93234 169262 93894 169402
rect 94062 169262 94722 169402
rect 94890 169262 95458 169402
rect 95626 169262 96286 169402
rect 96454 169262 97114 169402
rect 97282 169262 97850 169402
rect 98018 169262 98678 169402
rect 98846 169262 99506 169402
rect 99674 169262 100242 169402
rect 100410 169262 101070 169402
rect 101238 169262 101898 169402
rect 102066 169262 102634 169402
rect 102802 169262 103462 169402
rect 103630 169262 104290 169402
rect 104458 169262 105118 169402
rect 105286 169262 105854 169402
rect 106022 169262 106682 169402
rect 106850 169262 107510 169402
rect 107678 169262 108246 169402
rect 108414 169262 109074 169402
rect 109242 169262 109902 169402
rect 110070 169262 110638 169402
rect 110806 169262 111466 169402
rect 111634 169262 112294 169402
rect 112462 169262 113122 169402
rect 113290 169262 113858 169402
rect 114026 169262 114686 169402
rect 114854 169262 115514 169402
rect 115682 169262 116250 169402
rect 116418 169262 117078 169402
rect 117246 169262 117906 169402
rect 118074 169262 118642 169402
rect 118810 169262 119470 169402
rect 119638 169262 120298 169402
rect 120466 169262 121034 169402
rect 121202 169262 121862 169402
rect 122030 169262 122690 169402
rect 122858 169262 123518 169402
rect 123686 169262 124254 169402
rect 124422 169262 125082 169402
rect 125250 169262 125910 169402
rect 126078 169262 126646 169402
rect 126814 169262 127474 169402
rect 127642 169262 128302 169402
rect 128470 169262 129038 169402
rect 129206 169262 129866 169402
rect 130034 169262 130694 169402
rect 130862 169262 131522 169402
rect 131690 169262 132258 169402
rect 132426 169262 133086 169402
rect 133254 169262 133914 169402
rect 134082 169262 134650 169402
rect 134818 169262 135478 169402
rect 135646 169262 136306 169402
rect 136474 169262 137042 169402
rect 137210 169262 137870 169402
rect 138038 169262 138698 169402
rect 138866 169262 139434 169402
rect 139602 169262 140262 169402
rect 140430 169262 141090 169402
rect 141258 169262 141918 169402
rect 142086 169262 142654 169402
rect 142822 169262 143482 169402
rect 143650 169262 144310 169402
rect 144478 169262 145046 169402
rect 145214 169262 145874 169402
rect 146042 169262 146702 169402
rect 146870 169262 147438 169402
rect 147606 169262 148266 169402
rect 148434 169262 149094 169402
rect 149262 169262 149922 169402
rect 150090 169262 150658 169402
rect 150826 169262 151486 169402
rect 151654 169262 152314 169402
rect 152482 169262 153050 169402
rect 153218 169262 153878 169402
rect 154046 169262 154706 169402
rect 154874 169262 155442 169402
rect 155610 169262 156270 169402
rect 156438 169262 157098 169402
rect 157266 169262 157834 169402
rect 158002 169262 158662 169402
rect 158830 169262 159490 169402
rect 159658 169262 160318 169402
rect 160486 169262 161054 169402
rect 161222 169262 161882 169402
rect 162050 169262 162710 169402
rect 162878 169262 163446 169402
rect 163614 169262 164274 169402
rect 164442 169262 165102 169402
rect 165270 169262 165838 169402
rect 166006 169262 166666 169402
rect 166834 169262 167494 169402
rect 20 856 167604 169262
rect 20 711 16706 856
rect 16874 711 50286 856
rect 50454 711 83866 856
rect 84034 711 117446 856
rect 117614 711 151026 856
rect 151194 711 167604 856
<< metal3 >>
rect 167174 169328 167974 169448
rect 167174 167832 167974 167952
rect 167174 166336 167974 166456
rect 167174 164976 167974 165096
rect 0 163480 800 163600
rect 167174 163480 167974 163600
rect 167174 161984 167974 162104
rect 167174 160624 167974 160744
rect 167174 159128 167974 159248
rect 167174 157632 167974 157752
rect 167174 156272 167974 156392
rect 167174 154776 167974 154896
rect 167174 153280 167974 153400
rect 167174 151920 167974 152040
rect 0 150424 800 150544
rect 167174 150424 167974 150544
rect 167174 148928 167974 149048
rect 167174 147432 167974 147552
rect 167174 146072 167974 146192
rect 167174 144576 167974 144696
rect 167174 143080 167974 143200
rect 167174 141720 167974 141840
rect 167174 140224 167974 140344
rect 167174 138728 167974 138848
rect 0 137368 800 137488
rect 167174 137368 167974 137488
rect 167174 135872 167974 135992
rect 167174 134376 167974 134496
rect 167174 133016 167974 133136
rect 167174 131520 167974 131640
rect 167174 130024 167974 130144
rect 167174 128528 167974 128648
rect 167174 127168 167974 127288
rect 167174 125672 167974 125792
rect 0 124312 800 124432
rect 167174 124176 167974 124296
rect 167174 122816 167974 122936
rect 167174 121320 167974 121440
rect 167174 119824 167974 119944
rect 167174 118464 167974 118584
rect 167174 116968 167974 117088
rect 167174 115472 167974 115592
rect 167174 114112 167974 114232
rect 167174 112616 167974 112736
rect 0 111120 800 111240
rect 167174 111120 167974 111240
rect 167174 109624 167974 109744
rect 167174 108264 167974 108384
rect 167174 106768 167974 106888
rect 167174 105272 167974 105392
rect 167174 103912 167974 104032
rect 167174 102416 167974 102536
rect 167174 100920 167974 101040
rect 167174 99560 167974 99680
rect 0 98064 800 98184
rect 167174 98064 167974 98184
rect 167174 96568 167974 96688
rect 167174 95208 167974 95328
rect 167174 93712 167974 93832
rect 167174 92216 167974 92336
rect 167174 90720 167974 90840
rect 167174 89360 167974 89480
rect 167174 87864 167974 87984
rect 167174 86368 167974 86488
rect 0 85008 800 85128
rect 167174 85008 167974 85128
rect 167174 83512 167974 83632
rect 167174 82016 167974 82136
rect 167174 80656 167974 80776
rect 167174 79160 167974 79280
rect 167174 77664 167974 77784
rect 167174 76304 167974 76424
rect 167174 74808 167974 74928
rect 167174 73312 167974 73432
rect 0 71952 800 72072
rect 167174 71816 167974 71936
rect 167174 70456 167974 70576
rect 167174 68960 167974 69080
rect 167174 67464 167974 67584
rect 167174 66104 167974 66224
rect 167174 64608 167974 64728
rect 167174 63112 167974 63232
rect 167174 61752 167974 61872
rect 167174 60256 167974 60376
rect 0 58760 800 58880
rect 167174 58760 167974 58880
rect 167174 57400 167974 57520
rect 167174 55904 167974 56024
rect 167174 54408 167974 54528
rect 167174 52912 167974 53032
rect 167174 51552 167974 51672
rect 167174 50056 167974 50176
rect 167174 48560 167974 48680
rect 167174 47200 167974 47320
rect 0 45704 800 45824
rect 167174 45704 167974 45824
rect 167174 44208 167974 44328
rect 167174 42848 167974 42968
rect 167174 41352 167974 41472
rect 167174 39856 167974 39976
rect 167174 38496 167974 38616
rect 167174 37000 167974 37120
rect 167174 35504 167974 35624
rect 167174 34008 167974 34128
rect 0 32648 800 32768
rect 167174 32648 167974 32768
rect 167174 31152 167974 31272
rect 167174 29656 167974 29776
rect 167174 28296 167974 28416
rect 167174 26800 167974 26920
rect 167174 25304 167974 25424
rect 167174 23944 167974 24064
rect 167174 22448 167974 22568
rect 167174 20952 167974 21072
rect 0 19592 800 19712
rect 167174 19592 167974 19712
rect 167174 18096 167974 18216
rect 167174 16600 167974 16720
rect 167174 15104 167974 15224
rect 167174 13744 167974 13864
rect 167174 12248 167974 12368
rect 167174 10752 167974 10872
rect 167174 9392 167974 9512
rect 167174 7896 167974 8016
rect 0 6536 800 6656
rect 167174 6400 167974 6520
rect 167174 5040 167974 5160
rect 167174 3544 167974 3664
rect 167174 2048 167974 2168
rect 167174 688 167974 808
<< obsm3 >>
rect 800 169248 167094 169418
rect 800 168032 167174 169248
rect 800 167752 167094 168032
rect 800 166536 167174 167752
rect 800 166256 167094 166536
rect 800 165176 167174 166256
rect 800 164896 167094 165176
rect 800 163680 167174 164896
rect 880 163400 167094 163680
rect 800 162184 167174 163400
rect 800 161904 167094 162184
rect 800 160824 167174 161904
rect 800 160544 167094 160824
rect 800 159328 167174 160544
rect 800 159048 167094 159328
rect 800 157832 167174 159048
rect 800 157552 167094 157832
rect 800 156472 167174 157552
rect 800 156192 167094 156472
rect 800 154976 167174 156192
rect 800 154696 167094 154976
rect 800 153480 167174 154696
rect 800 153200 167094 153480
rect 800 152120 167174 153200
rect 800 151840 167094 152120
rect 800 150624 167174 151840
rect 880 150344 167094 150624
rect 800 149128 167174 150344
rect 800 148848 167094 149128
rect 800 147632 167174 148848
rect 800 147352 167094 147632
rect 800 146272 167174 147352
rect 800 145992 167094 146272
rect 800 144776 167174 145992
rect 800 144496 167094 144776
rect 800 143280 167174 144496
rect 800 143000 167094 143280
rect 800 141920 167174 143000
rect 800 141640 167094 141920
rect 800 140424 167174 141640
rect 800 140144 167094 140424
rect 800 138928 167174 140144
rect 800 138648 167094 138928
rect 800 137568 167174 138648
rect 880 137288 167094 137568
rect 800 136072 167174 137288
rect 800 135792 167094 136072
rect 800 134576 167174 135792
rect 800 134296 167094 134576
rect 800 133216 167174 134296
rect 800 132936 167094 133216
rect 800 131720 167174 132936
rect 800 131440 167094 131720
rect 800 130224 167174 131440
rect 800 129944 167094 130224
rect 800 128728 167174 129944
rect 800 128448 167094 128728
rect 800 127368 167174 128448
rect 800 127088 167094 127368
rect 800 125872 167174 127088
rect 800 125592 167094 125872
rect 800 124512 167174 125592
rect 880 124376 167174 124512
rect 880 124232 167094 124376
rect 800 124096 167094 124232
rect 800 123016 167174 124096
rect 800 122736 167094 123016
rect 800 121520 167174 122736
rect 800 121240 167094 121520
rect 800 120024 167174 121240
rect 800 119744 167094 120024
rect 800 118664 167174 119744
rect 800 118384 167094 118664
rect 800 117168 167174 118384
rect 800 116888 167094 117168
rect 800 115672 167174 116888
rect 800 115392 167094 115672
rect 800 114312 167174 115392
rect 800 114032 167094 114312
rect 800 112816 167174 114032
rect 800 112536 167094 112816
rect 800 111320 167174 112536
rect 880 111040 167094 111320
rect 800 109824 167174 111040
rect 800 109544 167094 109824
rect 800 108464 167174 109544
rect 800 108184 167094 108464
rect 800 106968 167174 108184
rect 800 106688 167094 106968
rect 800 105472 167174 106688
rect 800 105192 167094 105472
rect 800 104112 167174 105192
rect 800 103832 167094 104112
rect 800 102616 167174 103832
rect 800 102336 167094 102616
rect 800 101120 167174 102336
rect 800 100840 167094 101120
rect 800 99760 167174 100840
rect 800 99480 167094 99760
rect 800 98264 167174 99480
rect 880 97984 167094 98264
rect 800 96768 167174 97984
rect 800 96488 167094 96768
rect 800 95408 167174 96488
rect 800 95128 167094 95408
rect 800 93912 167174 95128
rect 800 93632 167094 93912
rect 800 92416 167174 93632
rect 800 92136 167094 92416
rect 800 90920 167174 92136
rect 800 90640 167094 90920
rect 800 89560 167174 90640
rect 800 89280 167094 89560
rect 800 88064 167174 89280
rect 800 87784 167094 88064
rect 800 86568 167174 87784
rect 800 86288 167094 86568
rect 800 85208 167174 86288
rect 880 84928 167094 85208
rect 800 83712 167174 84928
rect 800 83432 167094 83712
rect 800 82216 167174 83432
rect 800 81936 167094 82216
rect 800 80856 167174 81936
rect 800 80576 167094 80856
rect 800 79360 167174 80576
rect 800 79080 167094 79360
rect 800 77864 167174 79080
rect 800 77584 167094 77864
rect 800 76504 167174 77584
rect 800 76224 167094 76504
rect 800 75008 167174 76224
rect 800 74728 167094 75008
rect 800 73512 167174 74728
rect 800 73232 167094 73512
rect 800 72152 167174 73232
rect 880 72016 167174 72152
rect 880 71872 167094 72016
rect 800 71736 167094 71872
rect 800 70656 167174 71736
rect 800 70376 167094 70656
rect 800 69160 167174 70376
rect 800 68880 167094 69160
rect 800 67664 167174 68880
rect 800 67384 167094 67664
rect 800 66304 167174 67384
rect 800 66024 167094 66304
rect 800 64808 167174 66024
rect 800 64528 167094 64808
rect 800 63312 167174 64528
rect 800 63032 167094 63312
rect 800 61952 167174 63032
rect 800 61672 167094 61952
rect 800 60456 167174 61672
rect 800 60176 167094 60456
rect 800 58960 167174 60176
rect 880 58680 167094 58960
rect 800 57600 167174 58680
rect 800 57320 167094 57600
rect 800 56104 167174 57320
rect 800 55824 167094 56104
rect 800 54608 167174 55824
rect 800 54328 167094 54608
rect 800 53112 167174 54328
rect 800 52832 167094 53112
rect 800 51752 167174 52832
rect 800 51472 167094 51752
rect 800 50256 167174 51472
rect 800 49976 167094 50256
rect 800 48760 167174 49976
rect 800 48480 167094 48760
rect 800 47400 167174 48480
rect 800 47120 167094 47400
rect 800 45904 167174 47120
rect 880 45624 167094 45904
rect 800 44408 167174 45624
rect 800 44128 167094 44408
rect 800 43048 167174 44128
rect 800 42768 167094 43048
rect 800 41552 167174 42768
rect 800 41272 167094 41552
rect 800 40056 167174 41272
rect 800 39776 167094 40056
rect 800 38696 167174 39776
rect 800 38416 167094 38696
rect 800 37200 167174 38416
rect 800 36920 167094 37200
rect 800 35704 167174 36920
rect 800 35424 167094 35704
rect 800 34208 167174 35424
rect 800 33928 167094 34208
rect 800 32848 167174 33928
rect 880 32568 167094 32848
rect 800 31352 167174 32568
rect 800 31072 167094 31352
rect 800 29856 167174 31072
rect 800 29576 167094 29856
rect 800 28496 167174 29576
rect 800 28216 167094 28496
rect 800 27000 167174 28216
rect 800 26720 167094 27000
rect 800 25504 167174 26720
rect 800 25224 167094 25504
rect 800 24144 167174 25224
rect 800 23864 167094 24144
rect 800 22648 167174 23864
rect 800 22368 167094 22648
rect 800 21152 167174 22368
rect 800 20872 167094 21152
rect 800 19792 167174 20872
rect 880 19512 167094 19792
rect 800 18296 167174 19512
rect 800 18016 167094 18296
rect 800 16800 167174 18016
rect 800 16520 167094 16800
rect 800 15304 167174 16520
rect 800 15024 167094 15304
rect 800 13944 167174 15024
rect 800 13664 167094 13944
rect 800 12448 167174 13664
rect 800 12168 167094 12448
rect 800 10952 167174 12168
rect 800 10672 167094 10952
rect 800 9592 167174 10672
rect 800 9312 167094 9592
rect 800 8096 167174 9312
rect 800 7816 167094 8096
rect 800 6736 167174 7816
rect 880 6600 167174 6736
rect 880 6456 167094 6600
rect 800 6320 167094 6456
rect 800 5240 167174 6320
rect 800 4960 167094 5240
rect 800 3744 167174 4960
rect 800 3464 167094 3744
rect 800 2248 167174 3464
rect 800 1968 167094 2248
rect 800 888 167174 1968
rect 800 715 167094 888
<< metal4 >>
rect 4208 2128 4528 167600
rect 19568 2128 19888 167600
rect 34928 2128 35248 167600
rect 50288 2128 50608 167600
rect 65648 2128 65968 167600
rect 81008 2128 81328 167600
rect 96368 2128 96688 167600
rect 111728 2128 112048 167600
rect 127088 2128 127408 167600
rect 142448 2128 142768 167600
rect 157808 2128 158128 167600
<< obsm4 >>
rect 19379 3707 19488 164525
rect 19968 3707 34848 164525
rect 35328 3707 50208 164525
rect 50688 3707 65568 164525
rect 66048 3707 80928 164525
rect 81408 3707 96288 164525
rect 96768 3707 111648 164525
rect 112128 3707 127008 164525
rect 127488 3707 142368 164525
rect 142848 3707 157728 164525
rect 158208 3707 165725 164525
<< labels >>
rlabel metal3 s 167174 154776 167974 154896 6 CLK
port 1 nsew signal input
rlabel metal2 s 386 169318 442 170118 6 EN_dmem_client_request_get
port 2 nsew signal input
rlabel metal2 s 1122 169318 1178 170118 6 EN_dmem_client_response_put
port 3 nsew signal input
rlabel metal2 s 109130 169318 109186 170118 6 EN_imem_client_request_get
port 4 nsew signal input
rlabel metal2 s 109958 169318 110014 170118 6 EN_imem_client_response_put
port 5 nsew signal input
rlabel metal2 s 1950 169318 2006 170118 6 RDY_dmem_client_request_get
port 6 nsew signal output
rlabel metal2 s 2778 169318 2834 170118 6 RDY_dmem_client_response_put
port 7 nsew signal output
rlabel metal2 s 110694 169318 110750 170118 6 RDY_imem_client_request_get
port 8 nsew signal output
rlabel metal2 s 111522 169318 111578 170118 6 RDY_imem_client_response_put
port 9 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 RDY_readPC
port 10 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 RST_N
port 11 nsew signal input
rlabel metal2 s 3514 169318 3570 170118 6 dmem_client_request_get[0]
port 12 nsew signal output
rlabel metal2 s 19522 169318 19578 170118 6 dmem_client_request_get[10]
port 13 nsew signal output
rlabel metal2 s 21178 169318 21234 170118 6 dmem_client_request_get[11]
port 14 nsew signal output
rlabel metal2 s 22742 169318 22798 170118 6 dmem_client_request_get[12]
port 15 nsew signal output
rlabel metal2 s 24306 169318 24362 170118 6 dmem_client_request_get[13]
port 16 nsew signal output
rlabel metal2 s 25962 169318 26018 170118 6 dmem_client_request_get[14]
port 17 nsew signal output
rlabel metal2 s 27526 169318 27582 170118 6 dmem_client_request_get[15]
port 18 nsew signal output
rlabel metal2 s 29182 169318 29238 170118 6 dmem_client_request_get[16]
port 19 nsew signal output
rlabel metal2 s 30746 169318 30802 170118 6 dmem_client_request_get[17]
port 20 nsew signal output
rlabel metal2 s 32310 169318 32366 170118 6 dmem_client_request_get[18]
port 21 nsew signal output
rlabel metal2 s 33966 169318 34022 170118 6 dmem_client_request_get[19]
port 22 nsew signal output
rlabel metal2 s 5170 169318 5226 170118 6 dmem_client_request_get[1]
port 23 nsew signal output
rlabel metal2 s 35530 169318 35586 170118 6 dmem_client_request_get[20]
port 24 nsew signal output
rlabel metal2 s 37094 169318 37150 170118 6 dmem_client_request_get[21]
port 25 nsew signal output
rlabel metal2 s 38750 169318 38806 170118 6 dmem_client_request_get[22]
port 26 nsew signal output
rlabel metal2 s 40314 169318 40370 170118 6 dmem_client_request_get[23]
port 27 nsew signal output
rlabel metal2 s 41970 169318 42026 170118 6 dmem_client_request_get[24]
port 28 nsew signal output
rlabel metal2 s 43534 169318 43590 170118 6 dmem_client_request_get[25]
port 29 nsew signal output
rlabel metal2 s 45098 169318 45154 170118 6 dmem_client_request_get[26]
port 30 nsew signal output
rlabel metal2 s 46754 169318 46810 170118 6 dmem_client_request_get[27]
port 31 nsew signal output
rlabel metal2 s 48318 169318 48374 170118 6 dmem_client_request_get[28]
port 32 nsew signal output
rlabel metal2 s 49974 169318 50030 170118 6 dmem_client_request_get[29]
port 33 nsew signal output
rlabel metal2 s 6734 169318 6790 170118 6 dmem_client_request_get[2]
port 34 nsew signal output
rlabel metal2 s 51538 169318 51594 170118 6 dmem_client_request_get[30]
port 35 nsew signal output
rlabel metal2 s 53102 169318 53158 170118 6 dmem_client_request_get[31]
port 36 nsew signal output
rlabel metal2 s 54758 169318 54814 170118 6 dmem_client_request_get[32]
port 37 nsew signal output
rlabel metal2 s 55494 169318 55550 170118 6 dmem_client_request_get[33]
port 38 nsew signal output
rlabel metal2 s 56322 169318 56378 170118 6 dmem_client_request_get[34]
port 39 nsew signal output
rlabel metal2 s 57150 169318 57206 170118 6 dmem_client_request_get[35]
port 40 nsew signal output
rlabel metal2 s 57978 169318 58034 170118 6 dmem_client_request_get[36]
port 41 nsew signal output
rlabel metal2 s 58714 169318 58770 170118 6 dmem_client_request_get[37]
port 42 nsew signal output
rlabel metal2 s 59542 169318 59598 170118 6 dmem_client_request_get[38]
port 43 nsew signal output
rlabel metal2 s 60370 169318 60426 170118 6 dmem_client_request_get[39]
port 44 nsew signal output
rlabel metal2 s 8298 169318 8354 170118 6 dmem_client_request_get[3]
port 45 nsew signal output
rlabel metal2 s 61106 169318 61162 170118 6 dmem_client_request_get[40]
port 46 nsew signal output
rlabel metal2 s 61934 169318 61990 170118 6 dmem_client_request_get[41]
port 47 nsew signal output
rlabel metal2 s 62762 169318 62818 170118 6 dmem_client_request_get[42]
port 48 nsew signal output
rlabel metal2 s 63498 169318 63554 170118 6 dmem_client_request_get[43]
port 49 nsew signal output
rlabel metal2 s 64326 169318 64382 170118 6 dmem_client_request_get[44]
port 50 nsew signal output
rlabel metal2 s 65154 169318 65210 170118 6 dmem_client_request_get[45]
port 51 nsew signal output
rlabel metal2 s 65982 169318 66038 170118 6 dmem_client_request_get[46]
port 52 nsew signal output
rlabel metal2 s 66718 169318 66774 170118 6 dmem_client_request_get[47]
port 53 nsew signal output
rlabel metal2 s 67546 169318 67602 170118 6 dmem_client_request_get[48]
port 54 nsew signal output
rlabel metal2 s 68374 169318 68430 170118 6 dmem_client_request_get[49]
port 55 nsew signal output
rlabel metal2 s 9954 169318 10010 170118 6 dmem_client_request_get[4]
port 56 nsew signal output
rlabel metal2 s 69110 169318 69166 170118 6 dmem_client_request_get[50]
port 57 nsew signal output
rlabel metal2 s 69938 169318 69994 170118 6 dmem_client_request_get[51]
port 58 nsew signal output
rlabel metal2 s 70766 169318 70822 170118 6 dmem_client_request_get[52]
port 59 nsew signal output
rlabel metal2 s 71502 169318 71558 170118 6 dmem_client_request_get[53]
port 60 nsew signal output
rlabel metal2 s 72330 169318 72386 170118 6 dmem_client_request_get[54]
port 61 nsew signal output
rlabel metal2 s 73158 169318 73214 170118 6 dmem_client_request_get[55]
port 62 nsew signal output
rlabel metal2 s 73894 169318 73950 170118 6 dmem_client_request_get[56]
port 63 nsew signal output
rlabel metal2 s 74722 169318 74778 170118 6 dmem_client_request_get[57]
port 64 nsew signal output
rlabel metal2 s 75550 169318 75606 170118 6 dmem_client_request_get[58]
port 65 nsew signal output
rlabel metal2 s 76378 169318 76434 170118 6 dmem_client_request_get[59]
port 66 nsew signal output
rlabel metal2 s 11518 169318 11574 170118 6 dmem_client_request_get[5]
port 67 nsew signal output
rlabel metal2 s 77114 169318 77170 170118 6 dmem_client_request_get[60]
port 68 nsew signal output
rlabel metal2 s 77942 169318 77998 170118 6 dmem_client_request_get[61]
port 69 nsew signal output
rlabel metal2 s 78770 169318 78826 170118 6 dmem_client_request_get[62]
port 70 nsew signal output
rlabel metal2 s 79506 169318 79562 170118 6 dmem_client_request_get[63]
port 71 nsew signal output
rlabel metal2 s 80334 169318 80390 170118 6 dmem_client_request_get[64]
port 72 nsew signal output
rlabel metal2 s 81162 169318 81218 170118 6 dmem_client_request_get[65]
port 73 nsew signal output
rlabel metal2 s 81898 169318 81954 170118 6 dmem_client_request_get[66]
port 74 nsew signal output
rlabel metal2 s 82726 169318 82782 170118 6 dmem_client_request_get[67]
port 75 nsew signal output
rlabel metal2 s 83554 169318 83610 170118 6 dmem_client_request_get[68]
port 76 nsew signal output
rlabel metal2 s 84382 169318 84438 170118 6 dmem_client_request_get[69]
port 77 nsew signal output
rlabel metal2 s 13174 169318 13230 170118 6 dmem_client_request_get[6]
port 78 nsew signal output
rlabel metal2 s 85118 169318 85174 170118 6 dmem_client_request_get[70]
port 79 nsew signal output
rlabel metal2 s 85946 169318 86002 170118 6 dmem_client_request_get[71]
port 80 nsew signal output
rlabel metal2 s 86774 169318 86830 170118 6 dmem_client_request_get[72]
port 81 nsew signal output
rlabel metal2 s 87510 169318 87566 170118 6 dmem_client_request_get[73]
port 82 nsew signal output
rlabel metal2 s 88338 169318 88394 170118 6 dmem_client_request_get[74]
port 83 nsew signal output
rlabel metal2 s 89166 169318 89222 170118 6 dmem_client_request_get[75]
port 84 nsew signal output
rlabel metal2 s 89902 169318 89958 170118 6 dmem_client_request_get[76]
port 85 nsew signal output
rlabel metal2 s 90730 169318 90786 170118 6 dmem_client_request_get[77]
port 86 nsew signal output
rlabel metal2 s 91558 169318 91614 170118 6 dmem_client_request_get[78]
port 87 nsew signal output
rlabel metal2 s 92294 169318 92350 170118 6 dmem_client_request_get[79]
port 88 nsew signal output
rlabel metal2 s 14738 169318 14794 170118 6 dmem_client_request_get[7]
port 89 nsew signal output
rlabel metal2 s 93122 169318 93178 170118 6 dmem_client_request_get[80]
port 90 nsew signal output
rlabel metal2 s 93950 169318 94006 170118 6 dmem_client_request_get[81]
port 91 nsew signal output
rlabel metal2 s 94778 169318 94834 170118 6 dmem_client_request_get[82]
port 92 nsew signal output
rlabel metal2 s 95514 169318 95570 170118 6 dmem_client_request_get[83]
port 93 nsew signal output
rlabel metal2 s 96342 169318 96398 170118 6 dmem_client_request_get[84]
port 94 nsew signal output
rlabel metal2 s 97170 169318 97226 170118 6 dmem_client_request_get[85]
port 95 nsew signal output
rlabel metal2 s 97906 169318 97962 170118 6 dmem_client_request_get[86]
port 96 nsew signal output
rlabel metal2 s 98734 169318 98790 170118 6 dmem_client_request_get[87]
port 97 nsew signal output
rlabel metal2 s 99562 169318 99618 170118 6 dmem_client_request_get[88]
port 98 nsew signal output
rlabel metal2 s 100298 169318 100354 170118 6 dmem_client_request_get[89]
port 99 nsew signal output
rlabel metal2 s 16302 169318 16358 170118 6 dmem_client_request_get[8]
port 100 nsew signal output
rlabel metal2 s 101126 169318 101182 170118 6 dmem_client_request_get[90]
port 101 nsew signal output
rlabel metal2 s 101954 169318 102010 170118 6 dmem_client_request_get[91]
port 102 nsew signal output
rlabel metal2 s 102690 169318 102746 170118 6 dmem_client_request_get[92]
port 103 nsew signal output
rlabel metal2 s 103518 169318 103574 170118 6 dmem_client_request_get[93]
port 104 nsew signal output
rlabel metal2 s 104346 169318 104402 170118 6 dmem_client_request_get[94]
port 105 nsew signal output
rlabel metal2 s 105174 169318 105230 170118 6 dmem_client_request_get[95]
port 106 nsew signal output
rlabel metal2 s 105910 169318 105966 170118 6 dmem_client_request_get[96]
port 107 nsew signal output
rlabel metal2 s 106738 169318 106794 170118 6 dmem_client_request_get[97]
port 108 nsew signal output
rlabel metal2 s 107566 169318 107622 170118 6 dmem_client_request_get[98]
port 109 nsew signal output
rlabel metal2 s 108302 169318 108358 170118 6 dmem_client_request_get[99]
port 110 nsew signal output
rlabel metal2 s 17958 169318 18014 170118 6 dmem_client_request_get[9]
port 111 nsew signal output
rlabel metal2 s 4342 169318 4398 170118 6 dmem_client_response_put[0]
port 112 nsew signal input
rlabel metal2 s 20350 169318 20406 170118 6 dmem_client_response_put[10]
port 113 nsew signal input
rlabel metal2 s 21914 169318 21970 170118 6 dmem_client_response_put[11]
port 114 nsew signal input
rlabel metal2 s 23570 169318 23626 170118 6 dmem_client_response_put[12]
port 115 nsew signal input
rlabel metal2 s 25134 169318 25190 170118 6 dmem_client_response_put[13]
port 116 nsew signal input
rlabel metal2 s 26698 169318 26754 170118 6 dmem_client_response_put[14]
port 117 nsew signal input
rlabel metal2 s 28354 169318 28410 170118 6 dmem_client_response_put[15]
port 118 nsew signal input
rlabel metal2 s 29918 169318 29974 170118 6 dmem_client_response_put[16]
port 119 nsew signal input
rlabel metal2 s 31574 169318 31630 170118 6 dmem_client_response_put[17]
port 120 nsew signal input
rlabel metal2 s 33138 169318 33194 170118 6 dmem_client_response_put[18]
port 121 nsew signal input
rlabel metal2 s 34702 169318 34758 170118 6 dmem_client_response_put[19]
port 122 nsew signal input
rlabel metal2 s 5906 169318 5962 170118 6 dmem_client_response_put[1]
port 123 nsew signal input
rlabel metal2 s 36358 169318 36414 170118 6 dmem_client_response_put[20]
port 124 nsew signal input
rlabel metal2 s 37922 169318 37978 170118 6 dmem_client_response_put[21]
port 125 nsew signal input
rlabel metal2 s 39578 169318 39634 170118 6 dmem_client_response_put[22]
port 126 nsew signal input
rlabel metal2 s 41142 169318 41198 170118 6 dmem_client_response_put[23]
port 127 nsew signal input
rlabel metal2 s 42706 169318 42762 170118 6 dmem_client_response_put[24]
port 128 nsew signal input
rlabel metal2 s 44362 169318 44418 170118 6 dmem_client_response_put[25]
port 129 nsew signal input
rlabel metal2 s 45926 169318 45982 170118 6 dmem_client_response_put[26]
port 130 nsew signal input
rlabel metal2 s 47582 169318 47638 170118 6 dmem_client_response_put[27]
port 131 nsew signal input
rlabel metal2 s 49146 169318 49202 170118 6 dmem_client_response_put[28]
port 132 nsew signal input
rlabel metal2 s 50710 169318 50766 170118 6 dmem_client_response_put[29]
port 133 nsew signal input
rlabel metal2 s 7562 169318 7618 170118 6 dmem_client_response_put[2]
port 134 nsew signal input
rlabel metal2 s 52366 169318 52422 170118 6 dmem_client_response_put[30]
port 135 nsew signal input
rlabel metal2 s 53930 169318 53986 170118 6 dmem_client_response_put[31]
port 136 nsew signal input
rlabel metal2 s 9126 169318 9182 170118 6 dmem_client_response_put[3]
port 137 nsew signal input
rlabel metal2 s 10782 169318 10838 170118 6 dmem_client_response_put[4]
port 138 nsew signal input
rlabel metal2 s 12346 169318 12402 170118 6 dmem_client_response_put[5]
port 139 nsew signal input
rlabel metal2 s 13910 169318 13966 170118 6 dmem_client_response_put[6]
port 140 nsew signal input
rlabel metal2 s 15566 169318 15622 170118 6 dmem_client_response_put[7]
port 141 nsew signal input
rlabel metal2 s 17130 169318 17186 170118 6 dmem_client_response_put[8]
port 142 nsew signal input
rlabel metal2 s 18694 169318 18750 170118 6 dmem_client_response_put[9]
port 143 nsew signal input
rlabel metal2 s 112350 169318 112406 170118 6 imem_client_request_get[0]
port 144 nsew signal output
rlabel metal2 s 128358 169318 128414 170118 6 imem_client_request_get[10]
port 145 nsew signal output
rlabel metal2 s 129922 169318 129978 170118 6 imem_client_request_get[11]
port 146 nsew signal output
rlabel metal2 s 131578 169318 131634 170118 6 imem_client_request_get[12]
port 147 nsew signal output
rlabel metal2 s 133142 169318 133198 170118 6 imem_client_request_get[13]
port 148 nsew signal output
rlabel metal2 s 134706 169318 134762 170118 6 imem_client_request_get[14]
port 149 nsew signal output
rlabel metal2 s 136362 169318 136418 170118 6 imem_client_request_get[15]
port 150 nsew signal output
rlabel metal2 s 137926 169318 137982 170118 6 imem_client_request_get[16]
port 151 nsew signal output
rlabel metal2 s 139490 169318 139546 170118 6 imem_client_request_get[17]
port 152 nsew signal output
rlabel metal2 s 141146 169318 141202 170118 6 imem_client_request_get[18]
port 153 nsew signal output
rlabel metal2 s 142710 169318 142766 170118 6 imem_client_request_get[19]
port 154 nsew signal output
rlabel metal2 s 113914 169318 113970 170118 6 imem_client_request_get[1]
port 155 nsew signal output
rlabel metal2 s 144366 169318 144422 170118 6 imem_client_request_get[20]
port 156 nsew signal output
rlabel metal2 s 145930 169318 145986 170118 6 imem_client_request_get[21]
port 157 nsew signal output
rlabel metal2 s 147494 169318 147550 170118 6 imem_client_request_get[22]
port 158 nsew signal output
rlabel metal2 s 149150 169318 149206 170118 6 imem_client_request_get[23]
port 159 nsew signal output
rlabel metal2 s 150714 169318 150770 170118 6 imem_client_request_get[24]
port 160 nsew signal output
rlabel metal2 s 152370 169318 152426 170118 6 imem_client_request_get[25]
port 161 nsew signal output
rlabel metal2 s 153934 169318 153990 170118 6 imem_client_request_get[26]
port 162 nsew signal output
rlabel metal2 s 155498 169318 155554 170118 6 imem_client_request_get[27]
port 163 nsew signal output
rlabel metal2 s 157154 169318 157210 170118 6 imem_client_request_get[28]
port 164 nsew signal output
rlabel metal2 s 158718 169318 158774 170118 6 imem_client_request_get[29]
port 165 nsew signal output
rlabel metal2 s 115570 169318 115626 170118 6 imem_client_request_get[2]
port 166 nsew signal output
rlabel metal2 s 160374 169318 160430 170118 6 imem_client_request_get[30]
port 167 nsew signal output
rlabel metal2 s 161938 169318 161994 170118 6 imem_client_request_get[31]
port 168 nsew signal output
rlabel metal2 s 117134 169318 117190 170118 6 imem_client_request_get[3]
port 169 nsew signal output
rlabel metal2 s 118698 169318 118754 170118 6 imem_client_request_get[4]
port 170 nsew signal output
rlabel metal2 s 120354 169318 120410 170118 6 imem_client_request_get[5]
port 171 nsew signal output
rlabel metal2 s 121918 169318 121974 170118 6 imem_client_request_get[6]
port 172 nsew signal output
rlabel metal2 s 123574 169318 123630 170118 6 imem_client_request_get[7]
port 173 nsew signal output
rlabel metal2 s 125138 169318 125194 170118 6 imem_client_request_get[8]
port 174 nsew signal output
rlabel metal2 s 126702 169318 126758 170118 6 imem_client_request_get[9]
port 175 nsew signal output
rlabel metal2 s 113178 169318 113234 170118 6 imem_client_response_put[0]
port 176 nsew signal input
rlabel metal2 s 129094 169318 129150 170118 6 imem_client_response_put[10]
port 177 nsew signal input
rlabel metal2 s 130750 169318 130806 170118 6 imem_client_response_put[11]
port 178 nsew signal input
rlabel metal2 s 132314 169318 132370 170118 6 imem_client_response_put[12]
port 179 nsew signal input
rlabel metal2 s 133970 169318 134026 170118 6 imem_client_response_put[13]
port 180 nsew signal input
rlabel metal2 s 135534 169318 135590 170118 6 imem_client_response_put[14]
port 181 nsew signal input
rlabel metal2 s 137098 169318 137154 170118 6 imem_client_response_put[15]
port 182 nsew signal input
rlabel metal2 s 138754 169318 138810 170118 6 imem_client_response_put[16]
port 183 nsew signal input
rlabel metal2 s 140318 169318 140374 170118 6 imem_client_response_put[17]
port 184 nsew signal input
rlabel metal2 s 141974 169318 142030 170118 6 imem_client_response_put[18]
port 185 nsew signal input
rlabel metal2 s 143538 169318 143594 170118 6 imem_client_response_put[19]
port 186 nsew signal input
rlabel metal2 s 114742 169318 114798 170118 6 imem_client_response_put[1]
port 187 nsew signal input
rlabel metal2 s 145102 169318 145158 170118 6 imem_client_response_put[20]
port 188 nsew signal input
rlabel metal2 s 146758 169318 146814 170118 6 imem_client_response_put[21]
port 189 nsew signal input
rlabel metal2 s 148322 169318 148378 170118 6 imem_client_response_put[22]
port 190 nsew signal input
rlabel metal2 s 149978 169318 150034 170118 6 imem_client_response_put[23]
port 191 nsew signal input
rlabel metal2 s 151542 169318 151598 170118 6 imem_client_response_put[24]
port 192 nsew signal input
rlabel metal2 s 153106 169318 153162 170118 6 imem_client_response_put[25]
port 193 nsew signal input
rlabel metal2 s 154762 169318 154818 170118 6 imem_client_response_put[26]
port 194 nsew signal input
rlabel metal2 s 156326 169318 156382 170118 6 imem_client_response_put[27]
port 195 nsew signal input
rlabel metal2 s 157890 169318 157946 170118 6 imem_client_response_put[28]
port 196 nsew signal input
rlabel metal2 s 159546 169318 159602 170118 6 imem_client_response_put[29]
port 197 nsew signal input
rlabel metal2 s 116306 169318 116362 170118 6 imem_client_response_put[2]
port 198 nsew signal input
rlabel metal2 s 161110 169318 161166 170118 6 imem_client_response_put[30]
port 199 nsew signal input
rlabel metal2 s 162766 169318 162822 170118 6 imem_client_response_put[31]
port 200 nsew signal input
rlabel metal2 s 117962 169318 118018 170118 6 imem_client_response_put[3]
port 201 nsew signal input
rlabel metal2 s 119526 169318 119582 170118 6 imem_client_response_put[4]
port 202 nsew signal input
rlabel metal2 s 121090 169318 121146 170118 6 imem_client_response_put[5]
port 203 nsew signal input
rlabel metal2 s 122746 169318 122802 170118 6 imem_client_response_put[6]
port 204 nsew signal input
rlabel metal2 s 124310 169318 124366 170118 6 imem_client_response_put[7]
port 205 nsew signal input
rlabel metal2 s 125966 169318 126022 170118 6 imem_client_response_put[8]
port 206 nsew signal input
rlabel metal2 s 127530 169318 127586 170118 6 imem_client_response_put[9]
port 207 nsew signal input
rlabel metal3 s 167174 156272 167974 156392 6 readPC[0]
port 208 nsew signal output
rlabel metal3 s 0 45704 800 45824 6 readPC[10]
port 209 nsew signal output
rlabel metal2 s 165158 169318 165214 170118 6 readPC[11]
port 210 nsew signal output
rlabel metal3 s 167174 161984 167974 162104 6 readPC[12]
port 211 nsew signal output
rlabel metal2 s 165894 169318 165950 170118 6 readPC[13]
port 212 nsew signal output
rlabel metal3 s 0 58760 800 58880 6 readPC[14]
port 213 nsew signal output
rlabel metal2 s 166722 169318 166778 170118 6 readPC[15]
port 214 nsew signal output
rlabel metal3 s 167174 163480 167974 163600 6 readPC[16]
port 215 nsew signal output
rlabel metal3 s 167174 164976 167974 165096 6 readPC[17]
port 216 nsew signal output
rlabel metal3 s 0 71952 800 72072 6 readPC[18]
port 217 nsew signal output
rlabel metal3 s 0 85008 800 85128 6 readPC[19]
port 218 nsew signal output
rlabel metal3 s 167174 157632 167974 157752 6 readPC[1]
port 219 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 readPC[20]
port 220 nsew signal output
rlabel metal3 s 0 98064 800 98184 6 readPC[21]
port 221 nsew signal output
rlabel metal3 s 167174 166336 167974 166456 6 readPC[22]
port 222 nsew signal output
rlabel metal2 s 151082 0 151138 800 6 readPC[23]
port 223 nsew signal output
rlabel metal3 s 167174 167832 167974 167952 6 readPC[24]
port 224 nsew signal output
rlabel metal3 s 0 111120 800 111240 6 readPC[25]
port 225 nsew signal output
rlabel metal3 s 0 124312 800 124432 6 readPC[26]
port 226 nsew signal output
rlabel metal3 s 0 137368 800 137488 6 readPC[27]
port 227 nsew signal output
rlabel metal3 s 167174 169328 167974 169448 6 readPC[28]
port 228 nsew signal output
rlabel metal2 s 167550 169318 167606 170118 6 readPC[29]
port 229 nsew signal output
rlabel metal3 s 167174 159128 167974 159248 6 readPC[2]
port 230 nsew signal output
rlabel metal3 s 0 150424 800 150544 6 readPC[30]
port 231 nsew signal output
rlabel metal3 s 0 163480 800 163600 6 readPC[31]
port 232 nsew signal output
rlabel metal3 s 167174 160624 167974 160744 6 readPC[3]
port 233 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 readPC[4]
port 234 nsew signal output
rlabel metal2 s 83922 0 83978 800 6 readPC[5]
port 235 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 readPC[6]
port 236 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 readPC[7]
port 237 nsew signal output
rlabel metal2 s 163502 169318 163558 170118 6 readPC[8]
port 238 nsew signal output
rlabel metal2 s 164330 169318 164386 170118 6 readPC[9]
port 239 nsew signal output
rlabel metal3 s 167174 688 167974 808 6 sysmem_client_ack_i
port 240 nsew signal input
rlabel metal3 s 167174 9392 167974 9512 6 sysmem_client_adr_o[0]
port 241 nsew signal output
rlabel metal3 s 167174 58760 167974 58880 6 sysmem_client_adr_o[10]
port 242 nsew signal output
rlabel metal3 s 167174 63112 167974 63232 6 sysmem_client_adr_o[11]
port 243 nsew signal output
rlabel metal3 s 167174 67464 167974 67584 6 sysmem_client_adr_o[12]
port 244 nsew signal output
rlabel metal3 s 167174 71816 167974 71936 6 sysmem_client_adr_o[13]
port 245 nsew signal output
rlabel metal3 s 167174 76304 167974 76424 6 sysmem_client_adr_o[14]
port 246 nsew signal output
rlabel metal3 s 167174 80656 167974 80776 6 sysmem_client_adr_o[15]
port 247 nsew signal output
rlabel metal3 s 167174 85008 167974 85128 6 sysmem_client_adr_o[16]
port 248 nsew signal output
rlabel metal3 s 167174 89360 167974 89480 6 sysmem_client_adr_o[17]
port 249 nsew signal output
rlabel metal3 s 167174 93712 167974 93832 6 sysmem_client_adr_o[18]
port 250 nsew signal output
rlabel metal3 s 167174 98064 167974 98184 6 sysmem_client_adr_o[19]
port 251 nsew signal output
rlabel metal3 s 167174 15104 167974 15224 6 sysmem_client_adr_o[1]
port 252 nsew signal output
rlabel metal3 s 167174 102416 167974 102536 6 sysmem_client_adr_o[20]
port 253 nsew signal output
rlabel metal3 s 167174 106768 167974 106888 6 sysmem_client_adr_o[21]
port 254 nsew signal output
rlabel metal3 s 167174 111120 167974 111240 6 sysmem_client_adr_o[22]
port 255 nsew signal output
rlabel metal3 s 167174 115472 167974 115592 6 sysmem_client_adr_o[23]
port 256 nsew signal output
rlabel metal3 s 167174 119824 167974 119944 6 sysmem_client_adr_o[24]
port 257 nsew signal output
rlabel metal3 s 167174 124176 167974 124296 6 sysmem_client_adr_o[25]
port 258 nsew signal output
rlabel metal3 s 167174 128528 167974 128648 6 sysmem_client_adr_o[26]
port 259 nsew signal output
rlabel metal3 s 167174 133016 167974 133136 6 sysmem_client_adr_o[27]
port 260 nsew signal output
rlabel metal3 s 167174 137368 167974 137488 6 sysmem_client_adr_o[28]
port 261 nsew signal output
rlabel metal3 s 167174 141720 167974 141840 6 sysmem_client_adr_o[29]
port 262 nsew signal output
rlabel metal3 s 167174 20952 167974 21072 6 sysmem_client_adr_o[2]
port 263 nsew signal output
rlabel metal3 s 167174 146072 167974 146192 6 sysmem_client_adr_o[30]
port 264 nsew signal output
rlabel metal3 s 167174 150424 167974 150544 6 sysmem_client_adr_o[31]
port 265 nsew signal output
rlabel metal3 s 167174 26800 167974 26920 6 sysmem_client_adr_o[3]
port 266 nsew signal output
rlabel metal3 s 167174 32648 167974 32768 6 sysmem_client_adr_o[4]
port 267 nsew signal output
rlabel metal3 s 167174 37000 167974 37120 6 sysmem_client_adr_o[5]
port 268 nsew signal output
rlabel metal3 s 167174 41352 167974 41472 6 sysmem_client_adr_o[6]
port 269 nsew signal output
rlabel metal3 s 167174 45704 167974 45824 6 sysmem_client_adr_o[7]
port 270 nsew signal output
rlabel metal3 s 167174 50056 167974 50176 6 sysmem_client_adr_o[8]
port 271 nsew signal output
rlabel metal3 s 167174 54408 167974 54528 6 sysmem_client_adr_o[9]
port 272 nsew signal output
rlabel metal3 s 167174 2048 167974 2168 6 sysmem_client_cyc_o
port 273 nsew signal output
rlabel metal3 s 167174 10752 167974 10872 6 sysmem_client_dat_i[0]
port 274 nsew signal input
rlabel metal3 s 167174 60256 167974 60376 6 sysmem_client_dat_i[10]
port 275 nsew signal input
rlabel metal3 s 167174 64608 167974 64728 6 sysmem_client_dat_i[11]
port 276 nsew signal input
rlabel metal3 s 167174 68960 167974 69080 6 sysmem_client_dat_i[12]
port 277 nsew signal input
rlabel metal3 s 167174 73312 167974 73432 6 sysmem_client_dat_i[13]
port 278 nsew signal input
rlabel metal3 s 167174 77664 167974 77784 6 sysmem_client_dat_i[14]
port 279 nsew signal input
rlabel metal3 s 167174 82016 167974 82136 6 sysmem_client_dat_i[15]
port 280 nsew signal input
rlabel metal3 s 167174 86368 167974 86488 6 sysmem_client_dat_i[16]
port 281 nsew signal input
rlabel metal3 s 167174 90720 167974 90840 6 sysmem_client_dat_i[17]
port 282 nsew signal input
rlabel metal3 s 167174 95208 167974 95328 6 sysmem_client_dat_i[18]
port 283 nsew signal input
rlabel metal3 s 167174 99560 167974 99680 6 sysmem_client_dat_i[19]
port 284 nsew signal input
rlabel metal3 s 167174 16600 167974 16720 6 sysmem_client_dat_i[1]
port 285 nsew signal input
rlabel metal3 s 167174 103912 167974 104032 6 sysmem_client_dat_i[20]
port 286 nsew signal input
rlabel metal3 s 167174 108264 167974 108384 6 sysmem_client_dat_i[21]
port 287 nsew signal input
rlabel metal3 s 167174 112616 167974 112736 6 sysmem_client_dat_i[22]
port 288 nsew signal input
rlabel metal3 s 167174 116968 167974 117088 6 sysmem_client_dat_i[23]
port 289 nsew signal input
rlabel metal3 s 167174 121320 167974 121440 6 sysmem_client_dat_i[24]
port 290 nsew signal input
rlabel metal3 s 167174 125672 167974 125792 6 sysmem_client_dat_i[25]
port 291 nsew signal input
rlabel metal3 s 167174 130024 167974 130144 6 sysmem_client_dat_i[26]
port 292 nsew signal input
rlabel metal3 s 167174 134376 167974 134496 6 sysmem_client_dat_i[27]
port 293 nsew signal input
rlabel metal3 s 167174 138728 167974 138848 6 sysmem_client_dat_i[28]
port 294 nsew signal input
rlabel metal3 s 167174 143080 167974 143200 6 sysmem_client_dat_i[29]
port 295 nsew signal input
rlabel metal3 s 167174 22448 167974 22568 6 sysmem_client_dat_i[2]
port 296 nsew signal input
rlabel metal3 s 167174 147432 167974 147552 6 sysmem_client_dat_i[30]
port 297 nsew signal input
rlabel metal3 s 167174 151920 167974 152040 6 sysmem_client_dat_i[31]
port 298 nsew signal input
rlabel metal3 s 167174 28296 167974 28416 6 sysmem_client_dat_i[3]
port 299 nsew signal input
rlabel metal3 s 167174 34008 167974 34128 6 sysmem_client_dat_i[4]
port 300 nsew signal input
rlabel metal3 s 167174 38496 167974 38616 6 sysmem_client_dat_i[5]
port 301 nsew signal input
rlabel metal3 s 167174 42848 167974 42968 6 sysmem_client_dat_i[6]
port 302 nsew signal input
rlabel metal3 s 167174 47200 167974 47320 6 sysmem_client_dat_i[7]
port 303 nsew signal input
rlabel metal3 s 167174 51552 167974 51672 6 sysmem_client_dat_i[8]
port 304 nsew signal input
rlabel metal3 s 167174 55904 167974 56024 6 sysmem_client_dat_i[9]
port 305 nsew signal input
rlabel metal3 s 167174 12248 167974 12368 6 sysmem_client_dat_o[0]
port 306 nsew signal output
rlabel metal3 s 167174 61752 167974 61872 6 sysmem_client_dat_o[10]
port 307 nsew signal output
rlabel metal3 s 167174 66104 167974 66224 6 sysmem_client_dat_o[11]
port 308 nsew signal output
rlabel metal3 s 167174 70456 167974 70576 6 sysmem_client_dat_o[12]
port 309 nsew signal output
rlabel metal3 s 167174 74808 167974 74928 6 sysmem_client_dat_o[13]
port 310 nsew signal output
rlabel metal3 s 167174 79160 167974 79280 6 sysmem_client_dat_o[14]
port 311 nsew signal output
rlabel metal3 s 167174 83512 167974 83632 6 sysmem_client_dat_o[15]
port 312 nsew signal output
rlabel metal3 s 167174 87864 167974 87984 6 sysmem_client_dat_o[16]
port 313 nsew signal output
rlabel metal3 s 167174 92216 167974 92336 6 sysmem_client_dat_o[17]
port 314 nsew signal output
rlabel metal3 s 167174 96568 167974 96688 6 sysmem_client_dat_o[18]
port 315 nsew signal output
rlabel metal3 s 167174 100920 167974 101040 6 sysmem_client_dat_o[19]
port 316 nsew signal output
rlabel metal3 s 167174 18096 167974 18216 6 sysmem_client_dat_o[1]
port 317 nsew signal output
rlabel metal3 s 167174 105272 167974 105392 6 sysmem_client_dat_o[20]
port 318 nsew signal output
rlabel metal3 s 167174 109624 167974 109744 6 sysmem_client_dat_o[21]
port 319 nsew signal output
rlabel metal3 s 167174 114112 167974 114232 6 sysmem_client_dat_o[22]
port 320 nsew signal output
rlabel metal3 s 167174 118464 167974 118584 6 sysmem_client_dat_o[23]
port 321 nsew signal output
rlabel metal3 s 167174 122816 167974 122936 6 sysmem_client_dat_o[24]
port 322 nsew signal output
rlabel metal3 s 167174 127168 167974 127288 6 sysmem_client_dat_o[25]
port 323 nsew signal output
rlabel metal3 s 167174 131520 167974 131640 6 sysmem_client_dat_o[26]
port 324 nsew signal output
rlabel metal3 s 167174 135872 167974 135992 6 sysmem_client_dat_o[27]
port 325 nsew signal output
rlabel metal3 s 167174 140224 167974 140344 6 sysmem_client_dat_o[28]
port 326 nsew signal output
rlabel metal3 s 167174 144576 167974 144696 6 sysmem_client_dat_o[29]
port 327 nsew signal output
rlabel metal3 s 167174 23944 167974 24064 6 sysmem_client_dat_o[2]
port 328 nsew signal output
rlabel metal3 s 167174 148928 167974 149048 6 sysmem_client_dat_o[30]
port 329 nsew signal output
rlabel metal3 s 167174 153280 167974 153400 6 sysmem_client_dat_o[31]
port 330 nsew signal output
rlabel metal3 s 167174 29656 167974 29776 6 sysmem_client_dat_o[3]
port 331 nsew signal output
rlabel metal3 s 167174 35504 167974 35624 6 sysmem_client_dat_o[4]
port 332 nsew signal output
rlabel metal3 s 167174 39856 167974 39976 6 sysmem_client_dat_o[5]
port 333 nsew signal output
rlabel metal3 s 167174 44208 167974 44328 6 sysmem_client_dat_o[6]
port 334 nsew signal output
rlabel metal3 s 167174 48560 167974 48680 6 sysmem_client_dat_o[7]
port 335 nsew signal output
rlabel metal3 s 167174 52912 167974 53032 6 sysmem_client_dat_o[8]
port 336 nsew signal output
rlabel metal3 s 167174 57400 167974 57520 6 sysmem_client_dat_o[9]
port 337 nsew signal output
rlabel metal3 s 167174 3544 167974 3664 6 sysmem_client_err_i
port 338 nsew signal input
rlabel metal3 s 167174 5040 167974 5160 6 sysmem_client_rty_i
port 339 nsew signal input
rlabel metal3 s 167174 13744 167974 13864 6 sysmem_client_sel_o[0]
port 340 nsew signal output
rlabel metal3 s 167174 19592 167974 19712 6 sysmem_client_sel_o[1]
port 341 nsew signal output
rlabel metal3 s 167174 25304 167974 25424 6 sysmem_client_sel_o[2]
port 342 nsew signal output
rlabel metal3 s 167174 31152 167974 31272 6 sysmem_client_sel_o[3]
port 343 nsew signal output
rlabel metal3 s 167174 6400 167974 6520 6 sysmem_client_stb_o
port 344 nsew signal output
rlabel metal3 s 167174 7896 167974 8016 6 sysmem_client_we_o
port 345 nsew signal output
rlabel metal4 s 4208 2128 4528 167600 6 vccd1
port 346 nsew power input
rlabel metal4 s 34928 2128 35248 167600 6 vccd1
port 346 nsew power input
rlabel metal4 s 65648 2128 65968 167600 6 vccd1
port 346 nsew power input
rlabel metal4 s 96368 2128 96688 167600 6 vccd1
port 346 nsew power input
rlabel metal4 s 127088 2128 127408 167600 6 vccd1
port 346 nsew power input
rlabel metal4 s 157808 2128 158128 167600 6 vccd1
port 346 nsew power input
rlabel metal4 s 19568 2128 19888 167600 6 vssd1
port 347 nsew ground input
rlabel metal4 s 50288 2128 50608 167600 6 vssd1
port 347 nsew ground input
rlabel metal4 s 81008 2128 81328 167600 6 vssd1
port 347 nsew ground input
rlabel metal4 s 111728 2128 112048 167600 6 vssd1
port 347 nsew ground input
rlabel metal4 s 142448 2128 142768 167600 6 vssd1
port 347 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 167974 170118
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 72069912
string GDS_FILE /home/q3k/sky130/qf105/openlane/mkLanaiCPU/runs/mkLanaiCPU/results/finishing/mkLanaiCPU.magic.gds
string GDS_START 1472604
<< end >>

