magic
tech sky130A
magscale 1 2
timestamp 1647788008
<< obsli1 >>
rect 1104 2159 158884 57681
<< obsm1 >>
rect 198 1300 159238 59220
<< metal2 >>
rect 202 59200 258 60000
rect 662 59200 718 60000
rect 1122 59200 1178 60000
rect 1674 59200 1730 60000
rect 2134 59200 2190 60000
rect 2686 59200 2742 60000
rect 3146 59200 3202 60000
rect 3698 59200 3754 60000
rect 4158 59200 4214 60000
rect 4710 59200 4766 60000
rect 5170 59200 5226 60000
rect 5722 59200 5778 60000
rect 6182 59200 6238 60000
rect 6734 59200 6790 60000
rect 7194 59200 7250 60000
rect 7746 59200 7802 60000
rect 8206 59200 8262 60000
rect 8666 59200 8722 60000
rect 9218 59200 9274 60000
rect 9678 59200 9734 60000
rect 10230 59200 10286 60000
rect 10690 59200 10746 60000
rect 11242 59200 11298 60000
rect 11702 59200 11758 60000
rect 12254 59200 12310 60000
rect 12714 59200 12770 60000
rect 13266 59200 13322 60000
rect 13726 59200 13782 60000
rect 14278 59200 14334 60000
rect 14738 59200 14794 60000
rect 15290 59200 15346 60000
rect 15750 59200 15806 60000
rect 16210 59200 16266 60000
rect 16762 59200 16818 60000
rect 17222 59200 17278 60000
rect 17774 59200 17830 60000
rect 18234 59200 18290 60000
rect 18786 59200 18842 60000
rect 19246 59200 19302 60000
rect 19798 59200 19854 60000
rect 20258 59200 20314 60000
rect 20810 59200 20866 60000
rect 21270 59200 21326 60000
rect 21822 59200 21878 60000
rect 22282 59200 22338 60000
rect 22834 59200 22890 60000
rect 23294 59200 23350 60000
rect 23846 59200 23902 60000
rect 24306 59200 24362 60000
rect 24766 59200 24822 60000
rect 25318 59200 25374 60000
rect 25778 59200 25834 60000
rect 26330 59200 26386 60000
rect 26790 59200 26846 60000
rect 27342 59200 27398 60000
rect 27802 59200 27858 60000
rect 28354 59200 28410 60000
rect 28814 59200 28870 60000
rect 29366 59200 29422 60000
rect 29826 59200 29882 60000
rect 30378 59200 30434 60000
rect 30838 59200 30894 60000
rect 31390 59200 31446 60000
rect 31850 59200 31906 60000
rect 32310 59200 32366 60000
rect 32862 59200 32918 60000
rect 33322 59200 33378 60000
rect 33874 59200 33930 60000
rect 34334 59200 34390 60000
rect 34886 59200 34942 60000
rect 35346 59200 35402 60000
rect 35898 59200 35954 60000
rect 36358 59200 36414 60000
rect 36910 59200 36966 60000
rect 37370 59200 37426 60000
rect 37922 59200 37978 60000
rect 38382 59200 38438 60000
rect 38934 59200 38990 60000
rect 39394 59200 39450 60000
rect 39946 59200 40002 60000
rect 40406 59200 40462 60000
rect 40866 59200 40922 60000
rect 41418 59200 41474 60000
rect 41878 59200 41934 60000
rect 42430 59200 42486 60000
rect 42890 59200 42946 60000
rect 43442 59200 43498 60000
rect 43902 59200 43958 60000
rect 44454 59200 44510 60000
rect 44914 59200 44970 60000
rect 45466 59200 45522 60000
rect 45926 59200 45982 60000
rect 46478 59200 46534 60000
rect 46938 59200 46994 60000
rect 47490 59200 47546 60000
rect 47950 59200 48006 60000
rect 48410 59200 48466 60000
rect 48962 59200 49018 60000
rect 49422 59200 49478 60000
rect 49974 59200 50030 60000
rect 50434 59200 50490 60000
rect 50986 59200 51042 60000
rect 51446 59200 51502 60000
rect 51998 59200 52054 60000
rect 52458 59200 52514 60000
rect 53010 59200 53066 60000
rect 53470 59200 53526 60000
rect 54022 59200 54078 60000
rect 54482 59200 54538 60000
rect 55034 59200 55090 60000
rect 55494 59200 55550 60000
rect 56046 59200 56102 60000
rect 56506 59200 56562 60000
rect 56966 59200 57022 60000
rect 57518 59200 57574 60000
rect 57978 59200 58034 60000
rect 58530 59200 58586 60000
rect 58990 59200 59046 60000
rect 59542 59200 59598 60000
rect 60002 59200 60058 60000
rect 60554 59200 60610 60000
rect 61014 59200 61070 60000
rect 61566 59200 61622 60000
rect 62026 59200 62082 60000
rect 62578 59200 62634 60000
rect 63038 59200 63094 60000
rect 63590 59200 63646 60000
rect 64050 59200 64106 60000
rect 64510 59200 64566 60000
rect 65062 59200 65118 60000
rect 65522 59200 65578 60000
rect 66074 59200 66130 60000
rect 66534 59200 66590 60000
rect 67086 59200 67142 60000
rect 67546 59200 67602 60000
rect 68098 59200 68154 60000
rect 68558 59200 68614 60000
rect 69110 59200 69166 60000
rect 69570 59200 69626 60000
rect 70122 59200 70178 60000
rect 70582 59200 70638 60000
rect 71134 59200 71190 60000
rect 71594 59200 71650 60000
rect 72146 59200 72202 60000
rect 72606 59200 72662 60000
rect 73066 59200 73122 60000
rect 73618 59200 73674 60000
rect 74078 59200 74134 60000
rect 74630 59200 74686 60000
rect 75090 59200 75146 60000
rect 75642 59200 75698 60000
rect 76102 59200 76158 60000
rect 76654 59200 76710 60000
rect 77114 59200 77170 60000
rect 77666 59200 77722 60000
rect 78126 59200 78182 60000
rect 78678 59200 78734 60000
rect 79138 59200 79194 60000
rect 79690 59200 79746 60000
rect 80150 59200 80206 60000
rect 80610 59200 80666 60000
rect 81162 59200 81218 60000
rect 81622 59200 81678 60000
rect 82174 59200 82230 60000
rect 82634 59200 82690 60000
rect 83186 59200 83242 60000
rect 83646 59200 83702 60000
rect 84198 59200 84254 60000
rect 84658 59200 84714 60000
rect 85210 59200 85266 60000
rect 85670 59200 85726 60000
rect 86222 59200 86278 60000
rect 86682 59200 86738 60000
rect 87234 59200 87290 60000
rect 87694 59200 87750 60000
rect 88154 59200 88210 60000
rect 88706 59200 88762 60000
rect 89166 59200 89222 60000
rect 89718 59200 89774 60000
rect 90178 59200 90234 60000
rect 90730 59200 90786 60000
rect 91190 59200 91246 60000
rect 91742 59200 91798 60000
rect 92202 59200 92258 60000
rect 92754 59200 92810 60000
rect 93214 59200 93270 60000
rect 93766 59200 93822 60000
rect 94226 59200 94282 60000
rect 94778 59200 94834 60000
rect 95238 59200 95294 60000
rect 95790 59200 95846 60000
rect 96250 59200 96306 60000
rect 96710 59200 96766 60000
rect 97262 59200 97318 60000
rect 97722 59200 97778 60000
rect 98274 59200 98330 60000
rect 98734 59200 98790 60000
rect 99286 59200 99342 60000
rect 99746 59200 99802 60000
rect 100298 59200 100354 60000
rect 100758 59200 100814 60000
rect 101310 59200 101366 60000
rect 101770 59200 101826 60000
rect 102322 59200 102378 60000
rect 102782 59200 102838 60000
rect 103334 59200 103390 60000
rect 103794 59200 103850 60000
rect 104254 59200 104310 60000
rect 104806 59200 104862 60000
rect 105266 59200 105322 60000
rect 105818 59200 105874 60000
rect 106278 59200 106334 60000
rect 106830 59200 106886 60000
rect 107290 59200 107346 60000
rect 107842 59200 107898 60000
rect 108302 59200 108358 60000
rect 108854 59200 108910 60000
rect 109314 59200 109370 60000
rect 109866 59200 109922 60000
rect 110326 59200 110382 60000
rect 110878 59200 110934 60000
rect 111338 59200 111394 60000
rect 111890 59200 111946 60000
rect 112350 59200 112406 60000
rect 112810 59200 112866 60000
rect 113362 59200 113418 60000
rect 113822 59200 113878 60000
rect 114374 59200 114430 60000
rect 114834 59200 114890 60000
rect 115386 59200 115442 60000
rect 115846 59200 115902 60000
rect 116398 59200 116454 60000
rect 116858 59200 116914 60000
rect 117410 59200 117466 60000
rect 117870 59200 117926 60000
rect 118422 59200 118478 60000
rect 118882 59200 118938 60000
rect 119434 59200 119490 60000
rect 119894 59200 119950 60000
rect 120354 59200 120410 60000
rect 120906 59200 120962 60000
rect 121366 59200 121422 60000
rect 121918 59200 121974 60000
rect 122378 59200 122434 60000
rect 122930 59200 122986 60000
rect 123390 59200 123446 60000
rect 123942 59200 123998 60000
rect 124402 59200 124458 60000
rect 124954 59200 125010 60000
rect 125414 59200 125470 60000
rect 125966 59200 126022 60000
rect 126426 59200 126482 60000
rect 126978 59200 127034 60000
rect 127438 59200 127494 60000
rect 127990 59200 128046 60000
rect 128450 59200 128506 60000
rect 128910 59200 128966 60000
rect 129462 59200 129518 60000
rect 129922 59200 129978 60000
rect 130474 59200 130530 60000
rect 130934 59200 130990 60000
rect 131486 59200 131542 60000
rect 131946 59200 132002 60000
rect 132498 59200 132554 60000
rect 132958 59200 133014 60000
rect 133510 59200 133566 60000
rect 133970 59200 134026 60000
rect 134522 59200 134578 60000
rect 134982 59200 135038 60000
rect 135534 59200 135590 60000
rect 135994 59200 136050 60000
rect 136454 59200 136510 60000
rect 137006 59200 137062 60000
rect 137466 59200 137522 60000
rect 138018 59200 138074 60000
rect 138478 59200 138534 60000
rect 139030 59200 139086 60000
rect 139490 59200 139546 60000
rect 140042 59200 140098 60000
rect 140502 59200 140558 60000
rect 141054 59200 141110 60000
rect 141514 59200 141570 60000
rect 142066 59200 142122 60000
rect 142526 59200 142582 60000
rect 143078 59200 143134 60000
rect 143538 59200 143594 60000
rect 144090 59200 144146 60000
rect 144550 59200 144606 60000
rect 145010 59200 145066 60000
rect 145562 59200 145618 60000
rect 146022 59200 146078 60000
rect 146574 59200 146630 60000
rect 147034 59200 147090 60000
rect 147586 59200 147642 60000
rect 148046 59200 148102 60000
rect 148598 59200 148654 60000
rect 149058 59200 149114 60000
rect 149610 59200 149666 60000
rect 150070 59200 150126 60000
rect 150622 59200 150678 60000
rect 151082 59200 151138 60000
rect 151634 59200 151690 60000
rect 152094 59200 152150 60000
rect 152554 59200 152610 60000
rect 153106 59200 153162 60000
rect 153566 59200 153622 60000
rect 154118 59200 154174 60000
rect 154578 59200 154634 60000
rect 155130 59200 155186 60000
rect 155590 59200 155646 60000
rect 156142 59200 156198 60000
rect 156602 59200 156658 60000
rect 157154 59200 157210 60000
rect 157614 59200 157670 60000
rect 158166 59200 158222 60000
rect 158626 59200 158682 60000
rect 159178 59200 159234 60000
rect 159638 59200 159694 60000
<< obsm2 >>
rect 314 59144 606 59945
rect 774 59144 1066 59945
rect 1234 59144 1618 59945
rect 1786 59144 2078 59945
rect 2246 59144 2630 59945
rect 2798 59144 3090 59945
rect 3258 59144 3642 59945
rect 3810 59144 4102 59945
rect 4270 59144 4654 59945
rect 4822 59144 5114 59945
rect 5282 59144 5666 59945
rect 5834 59144 6126 59945
rect 6294 59144 6678 59945
rect 6846 59144 7138 59945
rect 7306 59144 7690 59945
rect 7858 59144 8150 59945
rect 8318 59144 8610 59945
rect 8778 59144 9162 59945
rect 9330 59144 9622 59945
rect 9790 59144 10174 59945
rect 10342 59144 10634 59945
rect 10802 59144 11186 59945
rect 11354 59144 11646 59945
rect 11814 59144 12198 59945
rect 12366 59144 12658 59945
rect 12826 59144 13210 59945
rect 13378 59144 13670 59945
rect 13838 59144 14222 59945
rect 14390 59144 14682 59945
rect 14850 59144 15234 59945
rect 15402 59144 15694 59945
rect 15862 59144 16154 59945
rect 16322 59144 16706 59945
rect 16874 59144 17166 59945
rect 17334 59144 17718 59945
rect 17886 59144 18178 59945
rect 18346 59144 18730 59945
rect 18898 59144 19190 59945
rect 19358 59144 19742 59945
rect 19910 59144 20202 59945
rect 20370 59144 20754 59945
rect 20922 59144 21214 59945
rect 21382 59144 21766 59945
rect 21934 59144 22226 59945
rect 22394 59144 22778 59945
rect 22946 59144 23238 59945
rect 23406 59144 23790 59945
rect 23958 59144 24250 59945
rect 24418 59144 24710 59945
rect 24878 59144 25262 59945
rect 25430 59144 25722 59945
rect 25890 59144 26274 59945
rect 26442 59144 26734 59945
rect 26902 59144 27286 59945
rect 27454 59144 27746 59945
rect 27914 59144 28298 59945
rect 28466 59144 28758 59945
rect 28926 59144 29310 59945
rect 29478 59144 29770 59945
rect 29938 59144 30322 59945
rect 30490 59144 30782 59945
rect 30950 59144 31334 59945
rect 31502 59144 31794 59945
rect 31962 59144 32254 59945
rect 32422 59144 32806 59945
rect 32974 59144 33266 59945
rect 33434 59144 33818 59945
rect 33986 59144 34278 59945
rect 34446 59144 34830 59945
rect 34998 59144 35290 59945
rect 35458 59144 35842 59945
rect 36010 59144 36302 59945
rect 36470 59144 36854 59945
rect 37022 59144 37314 59945
rect 37482 59144 37866 59945
rect 38034 59144 38326 59945
rect 38494 59144 38878 59945
rect 39046 59144 39338 59945
rect 39506 59144 39890 59945
rect 40058 59144 40350 59945
rect 40518 59144 40810 59945
rect 40978 59144 41362 59945
rect 41530 59144 41822 59945
rect 41990 59144 42374 59945
rect 42542 59144 42834 59945
rect 43002 59144 43386 59945
rect 43554 59144 43846 59945
rect 44014 59144 44398 59945
rect 44566 59144 44858 59945
rect 45026 59144 45410 59945
rect 45578 59144 45870 59945
rect 46038 59144 46422 59945
rect 46590 59144 46882 59945
rect 47050 59144 47434 59945
rect 47602 59144 47894 59945
rect 48062 59144 48354 59945
rect 48522 59144 48906 59945
rect 49074 59144 49366 59945
rect 49534 59144 49918 59945
rect 50086 59144 50378 59945
rect 50546 59144 50930 59945
rect 51098 59144 51390 59945
rect 51558 59144 51942 59945
rect 52110 59144 52402 59945
rect 52570 59144 52954 59945
rect 53122 59144 53414 59945
rect 53582 59144 53966 59945
rect 54134 59144 54426 59945
rect 54594 59144 54978 59945
rect 55146 59144 55438 59945
rect 55606 59144 55990 59945
rect 56158 59144 56450 59945
rect 56618 59144 56910 59945
rect 57078 59144 57462 59945
rect 57630 59144 57922 59945
rect 58090 59144 58474 59945
rect 58642 59144 58934 59945
rect 59102 59144 59486 59945
rect 59654 59144 59946 59945
rect 60114 59144 60498 59945
rect 60666 59144 60958 59945
rect 61126 59144 61510 59945
rect 61678 59144 61970 59945
rect 62138 59144 62522 59945
rect 62690 59144 62982 59945
rect 63150 59144 63534 59945
rect 63702 59144 63994 59945
rect 64162 59144 64454 59945
rect 64622 59144 65006 59945
rect 65174 59144 65466 59945
rect 65634 59144 66018 59945
rect 66186 59144 66478 59945
rect 66646 59144 67030 59945
rect 67198 59144 67490 59945
rect 67658 59144 68042 59945
rect 68210 59144 68502 59945
rect 68670 59144 69054 59945
rect 69222 59144 69514 59945
rect 69682 59144 70066 59945
rect 70234 59144 70526 59945
rect 70694 59144 71078 59945
rect 71246 59144 71538 59945
rect 71706 59144 72090 59945
rect 72258 59144 72550 59945
rect 72718 59144 73010 59945
rect 73178 59144 73562 59945
rect 73730 59144 74022 59945
rect 74190 59144 74574 59945
rect 74742 59144 75034 59945
rect 75202 59144 75586 59945
rect 75754 59144 76046 59945
rect 76214 59144 76598 59945
rect 76766 59144 77058 59945
rect 77226 59144 77610 59945
rect 77778 59144 78070 59945
rect 78238 59144 78622 59945
rect 78790 59144 79082 59945
rect 79250 59144 79634 59945
rect 79802 59144 80094 59945
rect 80262 59144 80554 59945
rect 80722 59144 81106 59945
rect 81274 59144 81566 59945
rect 81734 59144 82118 59945
rect 82286 59144 82578 59945
rect 82746 59144 83130 59945
rect 83298 59144 83590 59945
rect 83758 59144 84142 59945
rect 84310 59144 84602 59945
rect 84770 59144 85154 59945
rect 85322 59144 85614 59945
rect 85782 59144 86166 59945
rect 86334 59144 86626 59945
rect 86794 59144 87178 59945
rect 87346 59144 87638 59945
rect 87806 59144 88098 59945
rect 88266 59144 88650 59945
rect 88818 59144 89110 59945
rect 89278 59144 89662 59945
rect 89830 59144 90122 59945
rect 90290 59144 90674 59945
rect 90842 59144 91134 59945
rect 91302 59144 91686 59945
rect 91854 59144 92146 59945
rect 92314 59144 92698 59945
rect 92866 59144 93158 59945
rect 93326 59144 93710 59945
rect 93878 59144 94170 59945
rect 94338 59144 94722 59945
rect 94890 59144 95182 59945
rect 95350 59144 95734 59945
rect 95902 59144 96194 59945
rect 96362 59144 96654 59945
rect 96822 59144 97206 59945
rect 97374 59144 97666 59945
rect 97834 59144 98218 59945
rect 98386 59144 98678 59945
rect 98846 59144 99230 59945
rect 99398 59144 99690 59945
rect 99858 59144 100242 59945
rect 100410 59144 100702 59945
rect 100870 59144 101254 59945
rect 101422 59144 101714 59945
rect 101882 59144 102266 59945
rect 102434 59144 102726 59945
rect 102894 59144 103278 59945
rect 103446 59144 103738 59945
rect 103906 59144 104198 59945
rect 104366 59144 104750 59945
rect 104918 59144 105210 59945
rect 105378 59144 105762 59945
rect 105930 59144 106222 59945
rect 106390 59144 106774 59945
rect 106942 59144 107234 59945
rect 107402 59144 107786 59945
rect 107954 59144 108246 59945
rect 108414 59144 108798 59945
rect 108966 59144 109258 59945
rect 109426 59144 109810 59945
rect 109978 59144 110270 59945
rect 110438 59144 110822 59945
rect 110990 59144 111282 59945
rect 111450 59144 111834 59945
rect 112002 59144 112294 59945
rect 112462 59144 112754 59945
rect 112922 59144 113306 59945
rect 113474 59144 113766 59945
rect 113934 59144 114318 59945
rect 114486 59144 114778 59945
rect 114946 59144 115330 59945
rect 115498 59144 115790 59945
rect 115958 59144 116342 59945
rect 116510 59144 116802 59945
rect 116970 59144 117354 59945
rect 117522 59144 117814 59945
rect 117982 59144 118366 59945
rect 118534 59144 118826 59945
rect 118994 59144 119378 59945
rect 119546 59144 119838 59945
rect 120006 59144 120298 59945
rect 120466 59144 120850 59945
rect 121018 59144 121310 59945
rect 121478 59144 121862 59945
rect 122030 59144 122322 59945
rect 122490 59144 122874 59945
rect 123042 59144 123334 59945
rect 123502 59144 123886 59945
rect 124054 59144 124346 59945
rect 124514 59144 124898 59945
rect 125066 59144 125358 59945
rect 125526 59144 125910 59945
rect 126078 59144 126370 59945
rect 126538 59144 126922 59945
rect 127090 59144 127382 59945
rect 127550 59144 127934 59945
rect 128102 59144 128394 59945
rect 128562 59144 128854 59945
rect 129022 59144 129406 59945
rect 129574 59144 129866 59945
rect 130034 59144 130418 59945
rect 130586 59144 130878 59945
rect 131046 59144 131430 59945
rect 131598 59144 131890 59945
rect 132058 59144 132442 59945
rect 132610 59144 132902 59945
rect 133070 59144 133454 59945
rect 133622 59144 133914 59945
rect 134082 59144 134466 59945
rect 134634 59144 134926 59945
rect 135094 59144 135478 59945
rect 135646 59144 135938 59945
rect 136106 59144 136398 59945
rect 136566 59144 136950 59945
rect 137118 59144 137410 59945
rect 137578 59144 137962 59945
rect 138130 59144 138422 59945
rect 138590 59144 138974 59945
rect 139142 59144 139434 59945
rect 139602 59144 139986 59945
rect 140154 59144 140446 59945
rect 140614 59144 140998 59945
rect 141166 59144 141458 59945
rect 141626 59144 142010 59945
rect 142178 59144 142470 59945
rect 142638 59144 143022 59945
rect 143190 59144 143482 59945
rect 143650 59144 144034 59945
rect 144202 59144 144494 59945
rect 144662 59144 144954 59945
rect 145122 59144 145506 59945
rect 145674 59144 145966 59945
rect 146134 59144 146518 59945
rect 146686 59144 146978 59945
rect 147146 59144 147530 59945
rect 147698 59144 147990 59945
rect 148158 59144 148542 59945
rect 148710 59144 149002 59945
rect 149170 59144 149554 59945
rect 149722 59144 150014 59945
rect 150182 59144 150566 59945
rect 150734 59144 151026 59945
rect 151194 59144 151578 59945
rect 151746 59144 152038 59945
rect 152206 59144 152498 59945
rect 152666 59144 153050 59945
rect 153218 59144 153510 59945
rect 153678 59144 154062 59945
rect 154230 59144 154522 59945
rect 154690 59144 155074 59945
rect 155242 59144 155534 59945
rect 155702 59144 156086 59945
rect 156254 59144 156546 59945
rect 156714 59144 157098 59945
rect 157266 59144 157558 59945
rect 157726 59144 158110 59945
rect 158278 59144 158570 59945
rect 158738 59144 159122 59945
rect 159290 59144 159582 59945
rect 204 303 159680 59144
<< metal3 >>
rect 0 59576 800 59696
rect 0 59032 800 59152
rect 0 58488 800 58608
rect 0 57944 800 58064
rect 0 57400 800 57520
rect 0 56856 800 56976
rect 0 56312 800 56432
rect 0 55768 800 55888
rect 0 55224 800 55344
rect 0 54680 800 54800
rect 0 54136 800 54256
rect 0 53592 800 53712
rect 0 52912 800 53032
rect 0 52368 800 52488
rect 0 51824 800 51944
rect 0 51280 800 51400
rect 0 50736 800 50856
rect 0 50192 800 50312
rect 0 49648 800 49768
rect 0 49104 800 49224
rect 0 48560 800 48680
rect 0 48016 800 48136
rect 0 47472 800 47592
rect 0 46928 800 47048
rect 0 46248 800 46368
rect 0 45704 800 45824
rect 0 45160 800 45280
rect 0 44616 800 44736
rect 0 44072 800 44192
rect 0 43528 800 43648
rect 0 42984 800 43104
rect 0 42440 800 42560
rect 0 41896 800 42016
rect 0 41352 800 41472
rect 0 40808 800 40928
rect 0 40264 800 40384
rect 0 39584 800 39704
rect 0 39040 800 39160
rect 0 38496 800 38616
rect 0 37952 800 38072
rect 0 37408 800 37528
rect 0 36864 800 36984
rect 0 36320 800 36440
rect 0 35776 800 35896
rect 0 35232 800 35352
rect 0 34688 800 34808
rect 0 34144 800 34264
rect 0 33600 800 33720
rect 0 32920 800 33040
rect 0 32376 800 32496
rect 0 31832 800 31952
rect 0 31288 800 31408
rect 0 30744 800 30864
rect 0 30200 800 30320
rect 0 29656 800 29776
rect 0 29112 800 29232
rect 0 28568 800 28688
rect 0 28024 800 28144
rect 0 27480 800 27600
rect 0 26936 800 27056
rect 0 26256 800 26376
rect 0 25712 800 25832
rect 0 25168 800 25288
rect 0 24624 800 24744
rect 0 24080 800 24200
rect 0 23536 800 23656
rect 0 22992 800 23112
rect 0 22448 800 22568
rect 0 21904 800 22024
rect 0 21360 800 21480
rect 0 20816 800 20936
rect 0 20272 800 20392
rect 0 19592 800 19712
rect 0 19048 800 19168
rect 0 18504 800 18624
rect 0 17960 800 18080
rect 0 17416 800 17536
rect 0 16872 800 16992
rect 0 16328 800 16448
rect 0 15784 800 15904
rect 0 15240 800 15360
rect 0 14696 800 14816
rect 0 14152 800 14272
rect 0 13608 800 13728
rect 0 12928 800 13048
rect 0 12384 800 12504
rect 0 11840 800 11960
rect 0 11296 800 11416
rect 0 10752 800 10872
rect 0 10208 800 10328
rect 0 9664 800 9784
rect 0 9120 800 9240
rect 0 8576 800 8696
rect 0 8032 800 8152
rect 0 7488 800 7608
rect 0 6944 800 7064
rect 0 6264 800 6384
rect 0 5720 800 5840
rect 0 5176 800 5296
rect 0 4632 800 4752
rect 0 4088 800 4208
rect 0 3544 800 3664
rect 0 3000 800 3120
rect 0 2456 800 2576
rect 0 1912 800 2032
rect 0 1368 800 1488
rect 0 824 800 944
rect 0 280 800 400
<< obsm3 >>
rect 800 59776 158128 59941
rect 880 59496 158128 59776
rect 800 59232 158128 59496
rect 880 58952 158128 59232
rect 800 58688 158128 58952
rect 880 58408 158128 58688
rect 800 58144 158128 58408
rect 880 57864 158128 58144
rect 800 57600 158128 57864
rect 880 57320 158128 57600
rect 800 57056 158128 57320
rect 880 56776 158128 57056
rect 800 56512 158128 56776
rect 880 56232 158128 56512
rect 800 55968 158128 56232
rect 880 55688 158128 55968
rect 800 55424 158128 55688
rect 880 55144 158128 55424
rect 800 54880 158128 55144
rect 880 54600 158128 54880
rect 800 54336 158128 54600
rect 880 54056 158128 54336
rect 800 53792 158128 54056
rect 880 53512 158128 53792
rect 800 53112 158128 53512
rect 880 52832 158128 53112
rect 800 52568 158128 52832
rect 880 52288 158128 52568
rect 800 52024 158128 52288
rect 880 51744 158128 52024
rect 800 51480 158128 51744
rect 880 51200 158128 51480
rect 800 50936 158128 51200
rect 880 50656 158128 50936
rect 800 50392 158128 50656
rect 880 50112 158128 50392
rect 800 49848 158128 50112
rect 880 49568 158128 49848
rect 800 49304 158128 49568
rect 880 49024 158128 49304
rect 800 48760 158128 49024
rect 880 48480 158128 48760
rect 800 48216 158128 48480
rect 880 47936 158128 48216
rect 800 47672 158128 47936
rect 880 47392 158128 47672
rect 800 47128 158128 47392
rect 880 46848 158128 47128
rect 800 46448 158128 46848
rect 880 46168 158128 46448
rect 800 45904 158128 46168
rect 880 45624 158128 45904
rect 800 45360 158128 45624
rect 880 45080 158128 45360
rect 800 44816 158128 45080
rect 880 44536 158128 44816
rect 800 44272 158128 44536
rect 880 43992 158128 44272
rect 800 43728 158128 43992
rect 880 43448 158128 43728
rect 800 43184 158128 43448
rect 880 42904 158128 43184
rect 800 42640 158128 42904
rect 880 42360 158128 42640
rect 800 42096 158128 42360
rect 880 41816 158128 42096
rect 800 41552 158128 41816
rect 880 41272 158128 41552
rect 800 41008 158128 41272
rect 880 40728 158128 41008
rect 800 40464 158128 40728
rect 880 40184 158128 40464
rect 800 39784 158128 40184
rect 880 39504 158128 39784
rect 800 39240 158128 39504
rect 880 38960 158128 39240
rect 800 38696 158128 38960
rect 880 38416 158128 38696
rect 800 38152 158128 38416
rect 880 37872 158128 38152
rect 800 37608 158128 37872
rect 880 37328 158128 37608
rect 800 37064 158128 37328
rect 880 36784 158128 37064
rect 800 36520 158128 36784
rect 880 36240 158128 36520
rect 800 35976 158128 36240
rect 880 35696 158128 35976
rect 800 35432 158128 35696
rect 880 35152 158128 35432
rect 800 34888 158128 35152
rect 880 34608 158128 34888
rect 800 34344 158128 34608
rect 880 34064 158128 34344
rect 800 33800 158128 34064
rect 880 33520 158128 33800
rect 800 33120 158128 33520
rect 880 32840 158128 33120
rect 800 32576 158128 32840
rect 880 32296 158128 32576
rect 800 32032 158128 32296
rect 880 31752 158128 32032
rect 800 31488 158128 31752
rect 880 31208 158128 31488
rect 800 30944 158128 31208
rect 880 30664 158128 30944
rect 800 30400 158128 30664
rect 880 30120 158128 30400
rect 800 29856 158128 30120
rect 880 29576 158128 29856
rect 800 29312 158128 29576
rect 880 29032 158128 29312
rect 800 28768 158128 29032
rect 880 28488 158128 28768
rect 800 28224 158128 28488
rect 880 27944 158128 28224
rect 800 27680 158128 27944
rect 880 27400 158128 27680
rect 800 27136 158128 27400
rect 880 26856 158128 27136
rect 800 26456 158128 26856
rect 880 26176 158128 26456
rect 800 25912 158128 26176
rect 880 25632 158128 25912
rect 800 25368 158128 25632
rect 880 25088 158128 25368
rect 800 24824 158128 25088
rect 880 24544 158128 24824
rect 800 24280 158128 24544
rect 880 24000 158128 24280
rect 800 23736 158128 24000
rect 880 23456 158128 23736
rect 800 23192 158128 23456
rect 880 22912 158128 23192
rect 800 22648 158128 22912
rect 880 22368 158128 22648
rect 800 22104 158128 22368
rect 880 21824 158128 22104
rect 800 21560 158128 21824
rect 880 21280 158128 21560
rect 800 21016 158128 21280
rect 880 20736 158128 21016
rect 800 20472 158128 20736
rect 880 20192 158128 20472
rect 800 19792 158128 20192
rect 880 19512 158128 19792
rect 800 19248 158128 19512
rect 880 18968 158128 19248
rect 800 18704 158128 18968
rect 880 18424 158128 18704
rect 800 18160 158128 18424
rect 880 17880 158128 18160
rect 800 17616 158128 17880
rect 880 17336 158128 17616
rect 800 17072 158128 17336
rect 880 16792 158128 17072
rect 800 16528 158128 16792
rect 880 16248 158128 16528
rect 800 15984 158128 16248
rect 880 15704 158128 15984
rect 800 15440 158128 15704
rect 880 15160 158128 15440
rect 800 14896 158128 15160
rect 880 14616 158128 14896
rect 800 14352 158128 14616
rect 880 14072 158128 14352
rect 800 13808 158128 14072
rect 880 13528 158128 13808
rect 800 13128 158128 13528
rect 880 12848 158128 13128
rect 800 12584 158128 12848
rect 880 12304 158128 12584
rect 800 12040 158128 12304
rect 880 11760 158128 12040
rect 800 11496 158128 11760
rect 880 11216 158128 11496
rect 800 10952 158128 11216
rect 880 10672 158128 10952
rect 800 10408 158128 10672
rect 880 10128 158128 10408
rect 800 9864 158128 10128
rect 880 9584 158128 9864
rect 800 9320 158128 9584
rect 880 9040 158128 9320
rect 800 8776 158128 9040
rect 880 8496 158128 8776
rect 800 8232 158128 8496
rect 880 7952 158128 8232
rect 800 7688 158128 7952
rect 880 7408 158128 7688
rect 800 7144 158128 7408
rect 880 6864 158128 7144
rect 800 6464 158128 6864
rect 880 6184 158128 6464
rect 800 5920 158128 6184
rect 880 5640 158128 5920
rect 800 5376 158128 5640
rect 880 5096 158128 5376
rect 800 4832 158128 5096
rect 880 4552 158128 4832
rect 800 4288 158128 4552
rect 880 4008 158128 4288
rect 800 3744 158128 4008
rect 880 3464 158128 3744
rect 800 3200 158128 3464
rect 880 2920 158128 3200
rect 800 2656 158128 2920
rect 880 2376 158128 2656
rect 800 2112 158128 2376
rect 880 1832 158128 2112
rect 800 1568 158128 1832
rect 880 1288 158128 1568
rect 800 1024 158128 1288
rect 880 744 158128 1024
rect 800 480 158128 744
rect 880 307 158128 480
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
rect 65648 2128 65968 57712
rect 81008 2128 81328 57712
rect 96368 2128 96688 57712
rect 111728 2128 112048 57712
rect 127088 2128 127408 57712
rect 142448 2128 142768 57712
rect 157808 2128 158128 57712
<< obsm4 >>
rect 2267 57792 151925 59941
rect 2267 26827 4128 57792
rect 4608 26827 19488 57792
rect 19968 26827 34848 57792
rect 35328 26827 50208 57792
rect 50688 26827 65568 57792
rect 66048 26827 80928 57792
rect 81408 26827 96288 57792
rect 96768 26827 111648 57792
rect 112128 26827 127008 57792
rect 127488 26827 142368 57792
rect 142848 26827 151925 57792
<< labels >>
rlabel metal3 s 0 280 800 400 6 CLK
port 1 nsew signal input
rlabel metal3 s 0 824 800 944 6 RST_N
port 2 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 cpu_ack_o
port 3 nsew signal output
rlabel metal3 s 0 4632 800 4752 6 cpu_adr_i[0]
port 4 nsew signal input
rlabel metal3 s 0 23536 800 23656 6 cpu_adr_i[10]
port 5 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 cpu_adr_i[11]
port 6 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 cpu_adr_i[12]
port 7 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 cpu_adr_i[13]
port 8 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 cpu_adr_i[14]
port 9 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 cpu_adr_i[15]
port 10 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 cpu_adr_i[16]
port 11 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 cpu_adr_i[17]
port 12 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 cpu_adr_i[18]
port 13 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 cpu_adr_i[19]
port 14 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 cpu_adr_i[1]
port 15 nsew signal input
rlabel metal3 s 0 40264 800 40384 6 cpu_adr_i[20]
port 16 nsew signal input
rlabel metal3 s 0 41896 800 42016 6 cpu_adr_i[21]
port 17 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 cpu_adr_i[22]
port 18 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 cpu_adr_i[23]
port 19 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 cpu_adr_i[24]
port 20 nsew signal input
rlabel metal3 s 0 48560 800 48680 6 cpu_adr_i[25]
port 21 nsew signal input
rlabel metal3 s 0 50192 800 50312 6 cpu_adr_i[26]
port 22 nsew signal input
rlabel metal3 s 0 51824 800 51944 6 cpu_adr_i[27]
port 23 nsew signal input
rlabel metal3 s 0 53592 800 53712 6 cpu_adr_i[28]
port 24 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 cpu_adr_i[29]
port 25 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 cpu_adr_i[2]
port 26 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 cpu_adr_i[30]
port 27 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 cpu_adr_i[31]
port 28 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 cpu_adr_i[3]
port 29 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 cpu_adr_i[4]
port 30 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 cpu_adr_i[5]
port 31 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 cpu_adr_i[6]
port 32 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 cpu_adr_i[7]
port 33 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 cpu_adr_i[8]
port 34 nsew signal input
rlabel metal3 s 0 21904 800 22024 6 cpu_adr_i[9]
port 35 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 cpu_cyc_i
port 36 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 cpu_dat_i[0]
port 37 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 cpu_dat_i[10]
port 38 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 cpu_dat_i[11]
port 39 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 cpu_dat_i[12]
port 40 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 cpu_dat_i[13]
port 41 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 cpu_dat_i[14]
port 42 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 cpu_dat_i[15]
port 43 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 cpu_dat_i[16]
port 44 nsew signal input
rlabel metal3 s 0 35776 800 35896 6 cpu_dat_i[17]
port 45 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 cpu_dat_i[18]
port 46 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 cpu_dat_i[19]
port 47 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 cpu_dat_i[1]
port 48 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 cpu_dat_i[20]
port 49 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 cpu_dat_i[21]
port 50 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 cpu_dat_i[22]
port 51 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 cpu_dat_i[23]
port 52 nsew signal input
rlabel metal3 s 0 47472 800 47592 6 cpu_dat_i[24]
port 53 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 cpu_dat_i[25]
port 54 nsew signal input
rlabel metal3 s 0 50736 800 50856 6 cpu_dat_i[26]
port 55 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 cpu_dat_i[27]
port 56 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 cpu_dat_i[28]
port 57 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 cpu_dat_i[29]
port 58 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 cpu_dat_i[2]
port 59 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 cpu_dat_i[30]
port 60 nsew signal input
rlabel metal3 s 0 59032 800 59152 6 cpu_dat_i[31]
port 61 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 cpu_dat_i[3]
port 62 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 cpu_dat_i[4]
port 63 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 cpu_dat_i[5]
port 64 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 cpu_dat_i[6]
port 65 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 cpu_dat_i[7]
port 66 nsew signal input
rlabel metal3 s 0 20816 800 20936 6 cpu_dat_i[8]
port 67 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 cpu_dat_i[9]
port 68 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 cpu_dat_o[0]
port 69 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 cpu_dat_o[10]
port 70 nsew signal output
rlabel metal3 s 0 26256 800 26376 6 cpu_dat_o[11]
port 71 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 cpu_dat_o[12]
port 72 nsew signal output
rlabel metal3 s 0 29656 800 29776 6 cpu_dat_o[13]
port 73 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 cpu_dat_o[14]
port 74 nsew signal output
rlabel metal3 s 0 32920 800 33040 6 cpu_dat_o[15]
port 75 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 cpu_dat_o[16]
port 76 nsew signal output
rlabel metal3 s 0 36320 800 36440 6 cpu_dat_o[17]
port 77 nsew signal output
rlabel metal3 s 0 37952 800 38072 6 cpu_dat_o[18]
port 78 nsew signal output
rlabel metal3 s 0 39584 800 39704 6 cpu_dat_o[19]
port 79 nsew signal output
rlabel metal3 s 0 8032 800 8152 6 cpu_dat_o[1]
port 80 nsew signal output
rlabel metal3 s 0 41352 800 41472 6 cpu_dat_o[20]
port 81 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 cpu_dat_o[21]
port 82 nsew signal output
rlabel metal3 s 0 44616 800 44736 6 cpu_dat_o[22]
port 83 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 cpu_dat_o[23]
port 84 nsew signal output
rlabel metal3 s 0 48016 800 48136 6 cpu_dat_o[24]
port 85 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 cpu_dat_o[25]
port 86 nsew signal output
rlabel metal3 s 0 51280 800 51400 6 cpu_dat_o[26]
port 87 nsew signal output
rlabel metal3 s 0 52912 800 53032 6 cpu_dat_o[27]
port 88 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 cpu_dat_o[28]
port 89 nsew signal output
rlabel metal3 s 0 56312 800 56432 6 cpu_dat_o[29]
port 90 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 cpu_dat_o[2]
port 91 nsew signal output
rlabel metal3 s 0 57944 800 58064 6 cpu_dat_o[30]
port 92 nsew signal output
rlabel metal3 s 0 59576 800 59696 6 cpu_dat_o[31]
port 93 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 cpu_dat_o[3]
port 94 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 cpu_dat_o[4]
port 95 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 cpu_dat_o[5]
port 96 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 cpu_dat_o[6]
port 97 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 cpu_dat_o[7]
port 98 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 cpu_dat_o[8]
port 99 nsew signal output
rlabel metal3 s 0 22992 800 23112 6 cpu_dat_o[9]
port 100 nsew signal output
rlabel metal3 s 0 2456 800 2576 6 cpu_err_o
port 101 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 cpu_rty_o
port 102 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 cpu_sel_i[0]
port 103 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 cpu_sel_i[1]
port 104 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 cpu_sel_i[2]
port 105 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 cpu_sel_i[3]
port 106 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 cpu_stb_i
port 107 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 cpu_we_i
port 108 nsew signal input
rlabel metal2 s 53470 59200 53526 60000 6 gpio_ack_i
port 109 nsew signal input
rlabel metal2 s 56506 59200 56562 60000 6 gpio_adr_o[0]
port 110 nsew signal output
rlabel metal2 s 73618 59200 73674 60000 6 gpio_adr_o[10]
port 111 nsew signal output
rlabel metal2 s 75090 59200 75146 60000 6 gpio_adr_o[11]
port 112 nsew signal output
rlabel metal2 s 76654 59200 76710 60000 6 gpio_adr_o[12]
port 113 nsew signal output
rlabel metal2 s 78126 59200 78182 60000 6 gpio_adr_o[13]
port 114 nsew signal output
rlabel metal2 s 79690 59200 79746 60000 6 gpio_adr_o[14]
port 115 nsew signal output
rlabel metal2 s 81162 59200 81218 60000 6 gpio_adr_o[15]
port 116 nsew signal output
rlabel metal2 s 82634 59200 82690 60000 6 gpio_adr_o[16]
port 117 nsew signal output
rlabel metal2 s 84198 59200 84254 60000 6 gpio_adr_o[17]
port 118 nsew signal output
rlabel metal2 s 85670 59200 85726 60000 6 gpio_adr_o[18]
port 119 nsew signal output
rlabel metal2 s 87234 59200 87290 60000 6 gpio_adr_o[19]
port 120 nsew signal output
rlabel metal2 s 58530 59200 58586 60000 6 gpio_adr_o[1]
port 121 nsew signal output
rlabel metal2 s 88706 59200 88762 60000 6 gpio_adr_o[20]
port 122 nsew signal output
rlabel metal2 s 90178 59200 90234 60000 6 gpio_adr_o[21]
port 123 nsew signal output
rlabel metal2 s 91742 59200 91798 60000 6 gpio_adr_o[22]
port 124 nsew signal output
rlabel metal2 s 93214 59200 93270 60000 6 gpio_adr_o[23]
port 125 nsew signal output
rlabel metal2 s 94778 59200 94834 60000 6 gpio_adr_o[24]
port 126 nsew signal output
rlabel metal2 s 96250 59200 96306 60000 6 gpio_adr_o[25]
port 127 nsew signal output
rlabel metal2 s 97722 59200 97778 60000 6 gpio_adr_o[26]
port 128 nsew signal output
rlabel metal2 s 99286 59200 99342 60000 6 gpio_adr_o[27]
port 129 nsew signal output
rlabel metal2 s 100758 59200 100814 60000 6 gpio_adr_o[28]
port 130 nsew signal output
rlabel metal2 s 102322 59200 102378 60000 6 gpio_adr_o[29]
port 131 nsew signal output
rlabel metal2 s 60554 59200 60610 60000 6 gpio_adr_o[2]
port 132 nsew signal output
rlabel metal2 s 103794 59200 103850 60000 6 gpio_adr_o[30]
port 133 nsew signal output
rlabel metal2 s 105266 59200 105322 60000 6 gpio_adr_o[31]
port 134 nsew signal output
rlabel metal2 s 62578 59200 62634 60000 6 gpio_adr_o[3]
port 135 nsew signal output
rlabel metal2 s 64510 59200 64566 60000 6 gpio_adr_o[4]
port 136 nsew signal output
rlabel metal2 s 66074 59200 66130 60000 6 gpio_adr_o[5]
port 137 nsew signal output
rlabel metal2 s 67546 59200 67602 60000 6 gpio_adr_o[6]
port 138 nsew signal output
rlabel metal2 s 69110 59200 69166 60000 6 gpio_adr_o[7]
port 139 nsew signal output
rlabel metal2 s 70582 59200 70638 60000 6 gpio_adr_o[8]
port 140 nsew signal output
rlabel metal2 s 72146 59200 72202 60000 6 gpio_adr_o[9]
port 141 nsew signal output
rlabel metal2 s 54022 59200 54078 60000 6 gpio_cyc_o
port 142 nsew signal output
rlabel metal2 s 56966 59200 57022 60000 6 gpio_dat_i[0]
port 143 nsew signal input
rlabel metal2 s 74078 59200 74134 60000 6 gpio_dat_i[10]
port 144 nsew signal input
rlabel metal2 s 75642 59200 75698 60000 6 gpio_dat_i[11]
port 145 nsew signal input
rlabel metal2 s 77114 59200 77170 60000 6 gpio_dat_i[12]
port 146 nsew signal input
rlabel metal2 s 78678 59200 78734 60000 6 gpio_dat_i[13]
port 147 nsew signal input
rlabel metal2 s 80150 59200 80206 60000 6 gpio_dat_i[14]
port 148 nsew signal input
rlabel metal2 s 81622 59200 81678 60000 6 gpio_dat_i[15]
port 149 nsew signal input
rlabel metal2 s 83186 59200 83242 60000 6 gpio_dat_i[16]
port 150 nsew signal input
rlabel metal2 s 84658 59200 84714 60000 6 gpio_dat_i[17]
port 151 nsew signal input
rlabel metal2 s 86222 59200 86278 60000 6 gpio_dat_i[18]
port 152 nsew signal input
rlabel metal2 s 87694 59200 87750 60000 6 gpio_dat_i[19]
port 153 nsew signal input
rlabel metal2 s 58990 59200 59046 60000 6 gpio_dat_i[1]
port 154 nsew signal input
rlabel metal2 s 89166 59200 89222 60000 6 gpio_dat_i[20]
port 155 nsew signal input
rlabel metal2 s 90730 59200 90786 60000 6 gpio_dat_i[21]
port 156 nsew signal input
rlabel metal2 s 92202 59200 92258 60000 6 gpio_dat_i[22]
port 157 nsew signal input
rlabel metal2 s 93766 59200 93822 60000 6 gpio_dat_i[23]
port 158 nsew signal input
rlabel metal2 s 95238 59200 95294 60000 6 gpio_dat_i[24]
port 159 nsew signal input
rlabel metal2 s 96710 59200 96766 60000 6 gpio_dat_i[25]
port 160 nsew signal input
rlabel metal2 s 98274 59200 98330 60000 6 gpio_dat_i[26]
port 161 nsew signal input
rlabel metal2 s 99746 59200 99802 60000 6 gpio_dat_i[27]
port 162 nsew signal input
rlabel metal2 s 101310 59200 101366 60000 6 gpio_dat_i[28]
port 163 nsew signal input
rlabel metal2 s 102782 59200 102838 60000 6 gpio_dat_i[29]
port 164 nsew signal input
rlabel metal2 s 61014 59200 61070 60000 6 gpio_dat_i[2]
port 165 nsew signal input
rlabel metal2 s 104254 59200 104310 60000 6 gpio_dat_i[30]
port 166 nsew signal input
rlabel metal2 s 105818 59200 105874 60000 6 gpio_dat_i[31]
port 167 nsew signal input
rlabel metal2 s 63038 59200 63094 60000 6 gpio_dat_i[3]
port 168 nsew signal input
rlabel metal2 s 65062 59200 65118 60000 6 gpio_dat_i[4]
port 169 nsew signal input
rlabel metal2 s 66534 59200 66590 60000 6 gpio_dat_i[5]
port 170 nsew signal input
rlabel metal2 s 68098 59200 68154 60000 6 gpio_dat_i[6]
port 171 nsew signal input
rlabel metal2 s 69570 59200 69626 60000 6 gpio_dat_i[7]
port 172 nsew signal input
rlabel metal2 s 71134 59200 71190 60000 6 gpio_dat_i[8]
port 173 nsew signal input
rlabel metal2 s 72606 59200 72662 60000 6 gpio_dat_i[9]
port 174 nsew signal input
rlabel metal2 s 57518 59200 57574 60000 6 gpio_dat_o[0]
port 175 nsew signal output
rlabel metal2 s 74630 59200 74686 60000 6 gpio_dat_o[10]
port 176 nsew signal output
rlabel metal2 s 76102 59200 76158 60000 6 gpio_dat_o[11]
port 177 nsew signal output
rlabel metal2 s 77666 59200 77722 60000 6 gpio_dat_o[12]
port 178 nsew signal output
rlabel metal2 s 79138 59200 79194 60000 6 gpio_dat_o[13]
port 179 nsew signal output
rlabel metal2 s 80610 59200 80666 60000 6 gpio_dat_o[14]
port 180 nsew signal output
rlabel metal2 s 82174 59200 82230 60000 6 gpio_dat_o[15]
port 181 nsew signal output
rlabel metal2 s 83646 59200 83702 60000 6 gpio_dat_o[16]
port 182 nsew signal output
rlabel metal2 s 85210 59200 85266 60000 6 gpio_dat_o[17]
port 183 nsew signal output
rlabel metal2 s 86682 59200 86738 60000 6 gpio_dat_o[18]
port 184 nsew signal output
rlabel metal2 s 88154 59200 88210 60000 6 gpio_dat_o[19]
port 185 nsew signal output
rlabel metal2 s 59542 59200 59598 60000 6 gpio_dat_o[1]
port 186 nsew signal output
rlabel metal2 s 89718 59200 89774 60000 6 gpio_dat_o[20]
port 187 nsew signal output
rlabel metal2 s 91190 59200 91246 60000 6 gpio_dat_o[21]
port 188 nsew signal output
rlabel metal2 s 92754 59200 92810 60000 6 gpio_dat_o[22]
port 189 nsew signal output
rlabel metal2 s 94226 59200 94282 60000 6 gpio_dat_o[23]
port 190 nsew signal output
rlabel metal2 s 95790 59200 95846 60000 6 gpio_dat_o[24]
port 191 nsew signal output
rlabel metal2 s 97262 59200 97318 60000 6 gpio_dat_o[25]
port 192 nsew signal output
rlabel metal2 s 98734 59200 98790 60000 6 gpio_dat_o[26]
port 193 nsew signal output
rlabel metal2 s 100298 59200 100354 60000 6 gpio_dat_o[27]
port 194 nsew signal output
rlabel metal2 s 101770 59200 101826 60000 6 gpio_dat_o[28]
port 195 nsew signal output
rlabel metal2 s 103334 59200 103390 60000 6 gpio_dat_o[29]
port 196 nsew signal output
rlabel metal2 s 61566 59200 61622 60000 6 gpio_dat_o[2]
port 197 nsew signal output
rlabel metal2 s 104806 59200 104862 60000 6 gpio_dat_o[30]
port 198 nsew signal output
rlabel metal2 s 106278 59200 106334 60000 6 gpio_dat_o[31]
port 199 nsew signal output
rlabel metal2 s 63590 59200 63646 60000 6 gpio_dat_o[3]
port 200 nsew signal output
rlabel metal2 s 65522 59200 65578 60000 6 gpio_dat_o[4]
port 201 nsew signal output
rlabel metal2 s 67086 59200 67142 60000 6 gpio_dat_o[5]
port 202 nsew signal output
rlabel metal2 s 68558 59200 68614 60000 6 gpio_dat_o[6]
port 203 nsew signal output
rlabel metal2 s 70122 59200 70178 60000 6 gpio_dat_o[7]
port 204 nsew signal output
rlabel metal2 s 71594 59200 71650 60000 6 gpio_dat_o[8]
port 205 nsew signal output
rlabel metal2 s 73066 59200 73122 60000 6 gpio_dat_o[9]
port 206 nsew signal output
rlabel metal2 s 54482 59200 54538 60000 6 gpio_err_i
port 207 nsew signal input
rlabel metal2 s 55034 59200 55090 60000 6 gpio_rty_i
port 208 nsew signal input
rlabel metal2 s 57978 59200 58034 60000 6 gpio_sel_o[0]
port 209 nsew signal output
rlabel metal2 s 60002 59200 60058 60000 6 gpio_sel_o[1]
port 210 nsew signal output
rlabel metal2 s 62026 59200 62082 60000 6 gpio_sel_o[2]
port 211 nsew signal output
rlabel metal2 s 64050 59200 64106 60000 6 gpio_sel_o[3]
port 212 nsew signal output
rlabel metal2 s 55494 59200 55550 60000 6 gpio_stb_o
port 213 nsew signal output
rlabel metal2 s 56046 59200 56102 60000 6 gpio_we_o
port 214 nsew signal output
rlabel metal2 s 106830 59200 106886 60000 6 ksc_ack_i
port 215 nsew signal input
rlabel metal2 s 109866 59200 109922 60000 6 ksc_adr_o[0]
port 216 nsew signal output
rlabel metal2 s 126978 59200 127034 60000 6 ksc_adr_o[10]
port 217 nsew signal output
rlabel metal2 s 128450 59200 128506 60000 6 ksc_adr_o[11]
port 218 nsew signal output
rlabel metal2 s 129922 59200 129978 60000 6 ksc_adr_o[12]
port 219 nsew signal output
rlabel metal2 s 131486 59200 131542 60000 6 ksc_adr_o[13]
port 220 nsew signal output
rlabel metal2 s 132958 59200 133014 60000 6 ksc_adr_o[14]
port 221 nsew signal output
rlabel metal2 s 134522 59200 134578 60000 6 ksc_adr_o[15]
port 222 nsew signal output
rlabel metal2 s 135994 59200 136050 60000 6 ksc_adr_o[16]
port 223 nsew signal output
rlabel metal2 s 137466 59200 137522 60000 6 ksc_adr_o[17]
port 224 nsew signal output
rlabel metal2 s 139030 59200 139086 60000 6 ksc_adr_o[18]
port 225 nsew signal output
rlabel metal2 s 140502 59200 140558 60000 6 ksc_adr_o[19]
port 226 nsew signal output
rlabel metal2 s 111890 59200 111946 60000 6 ksc_adr_o[1]
port 227 nsew signal output
rlabel metal2 s 142066 59200 142122 60000 6 ksc_adr_o[20]
port 228 nsew signal output
rlabel metal2 s 143538 59200 143594 60000 6 ksc_adr_o[21]
port 229 nsew signal output
rlabel metal2 s 145010 59200 145066 60000 6 ksc_adr_o[22]
port 230 nsew signal output
rlabel metal2 s 146574 59200 146630 60000 6 ksc_adr_o[23]
port 231 nsew signal output
rlabel metal2 s 148046 59200 148102 60000 6 ksc_adr_o[24]
port 232 nsew signal output
rlabel metal2 s 149610 59200 149666 60000 6 ksc_adr_o[25]
port 233 nsew signal output
rlabel metal2 s 151082 59200 151138 60000 6 ksc_adr_o[26]
port 234 nsew signal output
rlabel metal2 s 152554 59200 152610 60000 6 ksc_adr_o[27]
port 235 nsew signal output
rlabel metal2 s 154118 59200 154174 60000 6 ksc_adr_o[28]
port 236 nsew signal output
rlabel metal2 s 155590 59200 155646 60000 6 ksc_adr_o[29]
port 237 nsew signal output
rlabel metal2 s 113822 59200 113878 60000 6 ksc_adr_o[2]
port 238 nsew signal output
rlabel metal2 s 157154 59200 157210 60000 6 ksc_adr_o[30]
port 239 nsew signal output
rlabel metal2 s 158626 59200 158682 60000 6 ksc_adr_o[31]
port 240 nsew signal output
rlabel metal2 s 115846 59200 115902 60000 6 ksc_adr_o[3]
port 241 nsew signal output
rlabel metal2 s 117870 59200 117926 60000 6 ksc_adr_o[4]
port 242 nsew signal output
rlabel metal2 s 119434 59200 119490 60000 6 ksc_adr_o[5]
port 243 nsew signal output
rlabel metal2 s 120906 59200 120962 60000 6 ksc_adr_o[6]
port 244 nsew signal output
rlabel metal2 s 122378 59200 122434 60000 6 ksc_adr_o[7]
port 245 nsew signal output
rlabel metal2 s 123942 59200 123998 60000 6 ksc_adr_o[8]
port 246 nsew signal output
rlabel metal2 s 125414 59200 125470 60000 6 ksc_adr_o[9]
port 247 nsew signal output
rlabel metal2 s 107290 59200 107346 60000 6 ksc_cyc_o
port 248 nsew signal output
rlabel metal2 s 110326 59200 110382 60000 6 ksc_dat_i[0]
port 249 nsew signal input
rlabel metal2 s 127438 59200 127494 60000 6 ksc_dat_i[10]
port 250 nsew signal input
rlabel metal2 s 128910 59200 128966 60000 6 ksc_dat_i[11]
port 251 nsew signal input
rlabel metal2 s 130474 59200 130530 60000 6 ksc_dat_i[12]
port 252 nsew signal input
rlabel metal2 s 131946 59200 132002 60000 6 ksc_dat_i[13]
port 253 nsew signal input
rlabel metal2 s 133510 59200 133566 60000 6 ksc_dat_i[14]
port 254 nsew signal input
rlabel metal2 s 134982 59200 135038 60000 6 ksc_dat_i[15]
port 255 nsew signal input
rlabel metal2 s 136454 59200 136510 60000 6 ksc_dat_i[16]
port 256 nsew signal input
rlabel metal2 s 138018 59200 138074 60000 6 ksc_dat_i[17]
port 257 nsew signal input
rlabel metal2 s 139490 59200 139546 60000 6 ksc_dat_i[18]
port 258 nsew signal input
rlabel metal2 s 141054 59200 141110 60000 6 ksc_dat_i[19]
port 259 nsew signal input
rlabel metal2 s 112350 59200 112406 60000 6 ksc_dat_i[1]
port 260 nsew signal input
rlabel metal2 s 142526 59200 142582 60000 6 ksc_dat_i[20]
port 261 nsew signal input
rlabel metal2 s 144090 59200 144146 60000 6 ksc_dat_i[21]
port 262 nsew signal input
rlabel metal2 s 145562 59200 145618 60000 6 ksc_dat_i[22]
port 263 nsew signal input
rlabel metal2 s 147034 59200 147090 60000 6 ksc_dat_i[23]
port 264 nsew signal input
rlabel metal2 s 148598 59200 148654 60000 6 ksc_dat_i[24]
port 265 nsew signal input
rlabel metal2 s 150070 59200 150126 60000 6 ksc_dat_i[25]
port 266 nsew signal input
rlabel metal2 s 151634 59200 151690 60000 6 ksc_dat_i[26]
port 267 nsew signal input
rlabel metal2 s 153106 59200 153162 60000 6 ksc_dat_i[27]
port 268 nsew signal input
rlabel metal2 s 154578 59200 154634 60000 6 ksc_dat_i[28]
port 269 nsew signal input
rlabel metal2 s 156142 59200 156198 60000 6 ksc_dat_i[29]
port 270 nsew signal input
rlabel metal2 s 114374 59200 114430 60000 6 ksc_dat_i[2]
port 271 nsew signal input
rlabel metal2 s 157614 59200 157670 60000 6 ksc_dat_i[30]
port 272 nsew signal input
rlabel metal2 s 159178 59200 159234 60000 6 ksc_dat_i[31]
port 273 nsew signal input
rlabel metal2 s 116398 59200 116454 60000 6 ksc_dat_i[3]
port 274 nsew signal input
rlabel metal2 s 118422 59200 118478 60000 6 ksc_dat_i[4]
port 275 nsew signal input
rlabel metal2 s 119894 59200 119950 60000 6 ksc_dat_i[5]
port 276 nsew signal input
rlabel metal2 s 121366 59200 121422 60000 6 ksc_dat_i[6]
port 277 nsew signal input
rlabel metal2 s 122930 59200 122986 60000 6 ksc_dat_i[7]
port 278 nsew signal input
rlabel metal2 s 124402 59200 124458 60000 6 ksc_dat_i[8]
port 279 nsew signal input
rlabel metal2 s 125966 59200 126022 60000 6 ksc_dat_i[9]
port 280 nsew signal input
rlabel metal2 s 110878 59200 110934 60000 6 ksc_dat_o[0]
port 281 nsew signal output
rlabel metal2 s 127990 59200 128046 60000 6 ksc_dat_o[10]
port 282 nsew signal output
rlabel metal2 s 129462 59200 129518 60000 6 ksc_dat_o[11]
port 283 nsew signal output
rlabel metal2 s 130934 59200 130990 60000 6 ksc_dat_o[12]
port 284 nsew signal output
rlabel metal2 s 132498 59200 132554 60000 6 ksc_dat_o[13]
port 285 nsew signal output
rlabel metal2 s 133970 59200 134026 60000 6 ksc_dat_o[14]
port 286 nsew signal output
rlabel metal2 s 135534 59200 135590 60000 6 ksc_dat_o[15]
port 287 nsew signal output
rlabel metal2 s 137006 59200 137062 60000 6 ksc_dat_o[16]
port 288 nsew signal output
rlabel metal2 s 138478 59200 138534 60000 6 ksc_dat_o[17]
port 289 nsew signal output
rlabel metal2 s 140042 59200 140098 60000 6 ksc_dat_o[18]
port 290 nsew signal output
rlabel metal2 s 141514 59200 141570 60000 6 ksc_dat_o[19]
port 291 nsew signal output
rlabel metal2 s 112810 59200 112866 60000 6 ksc_dat_o[1]
port 292 nsew signal output
rlabel metal2 s 143078 59200 143134 60000 6 ksc_dat_o[20]
port 293 nsew signal output
rlabel metal2 s 144550 59200 144606 60000 6 ksc_dat_o[21]
port 294 nsew signal output
rlabel metal2 s 146022 59200 146078 60000 6 ksc_dat_o[22]
port 295 nsew signal output
rlabel metal2 s 147586 59200 147642 60000 6 ksc_dat_o[23]
port 296 nsew signal output
rlabel metal2 s 149058 59200 149114 60000 6 ksc_dat_o[24]
port 297 nsew signal output
rlabel metal2 s 150622 59200 150678 60000 6 ksc_dat_o[25]
port 298 nsew signal output
rlabel metal2 s 152094 59200 152150 60000 6 ksc_dat_o[26]
port 299 nsew signal output
rlabel metal2 s 153566 59200 153622 60000 6 ksc_dat_o[27]
port 300 nsew signal output
rlabel metal2 s 155130 59200 155186 60000 6 ksc_dat_o[28]
port 301 nsew signal output
rlabel metal2 s 156602 59200 156658 60000 6 ksc_dat_o[29]
port 302 nsew signal output
rlabel metal2 s 114834 59200 114890 60000 6 ksc_dat_o[2]
port 303 nsew signal output
rlabel metal2 s 158166 59200 158222 60000 6 ksc_dat_o[30]
port 304 nsew signal output
rlabel metal2 s 159638 59200 159694 60000 6 ksc_dat_o[31]
port 305 nsew signal output
rlabel metal2 s 116858 59200 116914 60000 6 ksc_dat_o[3]
port 306 nsew signal output
rlabel metal2 s 118882 59200 118938 60000 6 ksc_dat_o[4]
port 307 nsew signal output
rlabel metal2 s 120354 59200 120410 60000 6 ksc_dat_o[5]
port 308 nsew signal output
rlabel metal2 s 121918 59200 121974 60000 6 ksc_dat_o[6]
port 309 nsew signal output
rlabel metal2 s 123390 59200 123446 60000 6 ksc_dat_o[7]
port 310 nsew signal output
rlabel metal2 s 124954 59200 125010 60000 6 ksc_dat_o[8]
port 311 nsew signal output
rlabel metal2 s 126426 59200 126482 60000 6 ksc_dat_o[9]
port 312 nsew signal output
rlabel metal2 s 107842 59200 107898 60000 6 ksc_err_i
port 313 nsew signal input
rlabel metal2 s 108302 59200 108358 60000 6 ksc_rty_i
port 314 nsew signal input
rlabel metal2 s 111338 59200 111394 60000 6 ksc_sel_o[0]
port 315 nsew signal output
rlabel metal2 s 113362 59200 113418 60000 6 ksc_sel_o[1]
port 316 nsew signal output
rlabel metal2 s 115386 59200 115442 60000 6 ksc_sel_o[2]
port 317 nsew signal output
rlabel metal2 s 117410 59200 117466 60000 6 ksc_sel_o[3]
port 318 nsew signal output
rlabel metal2 s 108854 59200 108910 60000 6 ksc_stb_o
port 319 nsew signal output
rlabel metal2 s 109314 59200 109370 60000 6 ksc_we_o
port 320 nsew signal output
rlabel metal2 s 202 59200 258 60000 6 spi_ack_i
port 321 nsew signal input
rlabel metal2 s 3146 59200 3202 60000 6 spi_adr_o[0]
port 322 nsew signal output
rlabel metal2 s 20258 59200 20314 60000 6 spi_adr_o[10]
port 323 nsew signal output
rlabel metal2 s 21822 59200 21878 60000 6 spi_adr_o[11]
port 324 nsew signal output
rlabel metal2 s 23294 59200 23350 60000 6 spi_adr_o[12]
port 325 nsew signal output
rlabel metal2 s 24766 59200 24822 60000 6 spi_adr_o[13]
port 326 nsew signal output
rlabel metal2 s 26330 59200 26386 60000 6 spi_adr_o[14]
port 327 nsew signal output
rlabel metal2 s 27802 59200 27858 60000 6 spi_adr_o[15]
port 328 nsew signal output
rlabel metal2 s 29366 59200 29422 60000 6 spi_adr_o[16]
port 329 nsew signal output
rlabel metal2 s 30838 59200 30894 60000 6 spi_adr_o[17]
port 330 nsew signal output
rlabel metal2 s 32310 59200 32366 60000 6 spi_adr_o[18]
port 331 nsew signal output
rlabel metal2 s 33874 59200 33930 60000 6 spi_adr_o[19]
port 332 nsew signal output
rlabel metal2 s 5170 59200 5226 60000 6 spi_adr_o[1]
port 333 nsew signal output
rlabel metal2 s 35346 59200 35402 60000 6 spi_adr_o[20]
port 334 nsew signal output
rlabel metal2 s 36910 59200 36966 60000 6 spi_adr_o[21]
port 335 nsew signal output
rlabel metal2 s 38382 59200 38438 60000 6 spi_adr_o[22]
port 336 nsew signal output
rlabel metal2 s 39946 59200 40002 60000 6 spi_adr_o[23]
port 337 nsew signal output
rlabel metal2 s 41418 59200 41474 60000 6 spi_adr_o[24]
port 338 nsew signal output
rlabel metal2 s 42890 59200 42946 60000 6 spi_adr_o[25]
port 339 nsew signal output
rlabel metal2 s 44454 59200 44510 60000 6 spi_adr_o[26]
port 340 nsew signal output
rlabel metal2 s 45926 59200 45982 60000 6 spi_adr_o[27]
port 341 nsew signal output
rlabel metal2 s 47490 59200 47546 60000 6 spi_adr_o[28]
port 342 nsew signal output
rlabel metal2 s 48962 59200 49018 60000 6 spi_adr_o[29]
port 343 nsew signal output
rlabel metal2 s 7194 59200 7250 60000 6 spi_adr_o[2]
port 344 nsew signal output
rlabel metal2 s 50434 59200 50490 60000 6 spi_adr_o[30]
port 345 nsew signal output
rlabel metal2 s 51998 59200 52054 60000 6 spi_adr_o[31]
port 346 nsew signal output
rlabel metal2 s 9218 59200 9274 60000 6 spi_adr_o[3]
port 347 nsew signal output
rlabel metal2 s 11242 59200 11298 60000 6 spi_adr_o[4]
port 348 nsew signal output
rlabel metal2 s 12714 59200 12770 60000 6 spi_adr_o[5]
port 349 nsew signal output
rlabel metal2 s 14278 59200 14334 60000 6 spi_adr_o[6]
port 350 nsew signal output
rlabel metal2 s 15750 59200 15806 60000 6 spi_adr_o[7]
port 351 nsew signal output
rlabel metal2 s 17222 59200 17278 60000 6 spi_adr_o[8]
port 352 nsew signal output
rlabel metal2 s 18786 59200 18842 60000 6 spi_adr_o[9]
port 353 nsew signal output
rlabel metal2 s 662 59200 718 60000 6 spi_cyc_o
port 354 nsew signal output
rlabel metal2 s 3698 59200 3754 60000 6 spi_dat_i[0]
port 355 nsew signal input
rlabel metal2 s 20810 59200 20866 60000 6 spi_dat_i[10]
port 356 nsew signal input
rlabel metal2 s 22282 59200 22338 60000 6 spi_dat_i[11]
port 357 nsew signal input
rlabel metal2 s 23846 59200 23902 60000 6 spi_dat_i[12]
port 358 nsew signal input
rlabel metal2 s 25318 59200 25374 60000 6 spi_dat_i[13]
port 359 nsew signal input
rlabel metal2 s 26790 59200 26846 60000 6 spi_dat_i[14]
port 360 nsew signal input
rlabel metal2 s 28354 59200 28410 60000 6 spi_dat_i[15]
port 361 nsew signal input
rlabel metal2 s 29826 59200 29882 60000 6 spi_dat_i[16]
port 362 nsew signal input
rlabel metal2 s 31390 59200 31446 60000 6 spi_dat_i[17]
port 363 nsew signal input
rlabel metal2 s 32862 59200 32918 60000 6 spi_dat_i[18]
port 364 nsew signal input
rlabel metal2 s 34334 59200 34390 60000 6 spi_dat_i[19]
port 365 nsew signal input
rlabel metal2 s 5722 59200 5778 60000 6 spi_dat_i[1]
port 366 nsew signal input
rlabel metal2 s 35898 59200 35954 60000 6 spi_dat_i[20]
port 367 nsew signal input
rlabel metal2 s 37370 59200 37426 60000 6 spi_dat_i[21]
port 368 nsew signal input
rlabel metal2 s 38934 59200 38990 60000 6 spi_dat_i[22]
port 369 nsew signal input
rlabel metal2 s 40406 59200 40462 60000 6 spi_dat_i[23]
port 370 nsew signal input
rlabel metal2 s 41878 59200 41934 60000 6 spi_dat_i[24]
port 371 nsew signal input
rlabel metal2 s 43442 59200 43498 60000 6 spi_dat_i[25]
port 372 nsew signal input
rlabel metal2 s 44914 59200 44970 60000 6 spi_dat_i[26]
port 373 nsew signal input
rlabel metal2 s 46478 59200 46534 60000 6 spi_dat_i[27]
port 374 nsew signal input
rlabel metal2 s 47950 59200 48006 60000 6 spi_dat_i[28]
port 375 nsew signal input
rlabel metal2 s 49422 59200 49478 60000 6 spi_dat_i[29]
port 376 nsew signal input
rlabel metal2 s 7746 59200 7802 60000 6 spi_dat_i[2]
port 377 nsew signal input
rlabel metal2 s 50986 59200 51042 60000 6 spi_dat_i[30]
port 378 nsew signal input
rlabel metal2 s 52458 59200 52514 60000 6 spi_dat_i[31]
port 379 nsew signal input
rlabel metal2 s 9678 59200 9734 60000 6 spi_dat_i[3]
port 380 nsew signal input
rlabel metal2 s 11702 59200 11758 60000 6 spi_dat_i[4]
port 381 nsew signal input
rlabel metal2 s 13266 59200 13322 60000 6 spi_dat_i[5]
port 382 nsew signal input
rlabel metal2 s 14738 59200 14794 60000 6 spi_dat_i[6]
port 383 nsew signal input
rlabel metal2 s 16210 59200 16266 60000 6 spi_dat_i[7]
port 384 nsew signal input
rlabel metal2 s 17774 59200 17830 60000 6 spi_dat_i[8]
port 385 nsew signal input
rlabel metal2 s 19246 59200 19302 60000 6 spi_dat_i[9]
port 386 nsew signal input
rlabel metal2 s 4158 59200 4214 60000 6 spi_dat_o[0]
port 387 nsew signal output
rlabel metal2 s 21270 59200 21326 60000 6 spi_dat_o[10]
port 388 nsew signal output
rlabel metal2 s 22834 59200 22890 60000 6 spi_dat_o[11]
port 389 nsew signal output
rlabel metal2 s 24306 59200 24362 60000 6 spi_dat_o[12]
port 390 nsew signal output
rlabel metal2 s 25778 59200 25834 60000 6 spi_dat_o[13]
port 391 nsew signal output
rlabel metal2 s 27342 59200 27398 60000 6 spi_dat_o[14]
port 392 nsew signal output
rlabel metal2 s 28814 59200 28870 60000 6 spi_dat_o[15]
port 393 nsew signal output
rlabel metal2 s 30378 59200 30434 60000 6 spi_dat_o[16]
port 394 nsew signal output
rlabel metal2 s 31850 59200 31906 60000 6 spi_dat_o[17]
port 395 nsew signal output
rlabel metal2 s 33322 59200 33378 60000 6 spi_dat_o[18]
port 396 nsew signal output
rlabel metal2 s 34886 59200 34942 60000 6 spi_dat_o[19]
port 397 nsew signal output
rlabel metal2 s 6182 59200 6238 60000 6 spi_dat_o[1]
port 398 nsew signal output
rlabel metal2 s 36358 59200 36414 60000 6 spi_dat_o[20]
port 399 nsew signal output
rlabel metal2 s 37922 59200 37978 60000 6 spi_dat_o[21]
port 400 nsew signal output
rlabel metal2 s 39394 59200 39450 60000 6 spi_dat_o[22]
port 401 nsew signal output
rlabel metal2 s 40866 59200 40922 60000 6 spi_dat_o[23]
port 402 nsew signal output
rlabel metal2 s 42430 59200 42486 60000 6 spi_dat_o[24]
port 403 nsew signal output
rlabel metal2 s 43902 59200 43958 60000 6 spi_dat_o[25]
port 404 nsew signal output
rlabel metal2 s 45466 59200 45522 60000 6 spi_dat_o[26]
port 405 nsew signal output
rlabel metal2 s 46938 59200 46994 60000 6 spi_dat_o[27]
port 406 nsew signal output
rlabel metal2 s 48410 59200 48466 60000 6 spi_dat_o[28]
port 407 nsew signal output
rlabel metal2 s 49974 59200 50030 60000 6 spi_dat_o[29]
port 408 nsew signal output
rlabel metal2 s 8206 59200 8262 60000 6 spi_dat_o[2]
port 409 nsew signal output
rlabel metal2 s 51446 59200 51502 60000 6 spi_dat_o[30]
port 410 nsew signal output
rlabel metal2 s 53010 59200 53066 60000 6 spi_dat_o[31]
port 411 nsew signal output
rlabel metal2 s 10230 59200 10286 60000 6 spi_dat_o[3]
port 412 nsew signal output
rlabel metal2 s 12254 59200 12310 60000 6 spi_dat_o[4]
port 413 nsew signal output
rlabel metal2 s 13726 59200 13782 60000 6 spi_dat_o[5]
port 414 nsew signal output
rlabel metal2 s 15290 59200 15346 60000 6 spi_dat_o[6]
port 415 nsew signal output
rlabel metal2 s 16762 59200 16818 60000 6 spi_dat_o[7]
port 416 nsew signal output
rlabel metal2 s 18234 59200 18290 60000 6 spi_dat_o[8]
port 417 nsew signal output
rlabel metal2 s 19798 59200 19854 60000 6 spi_dat_o[9]
port 418 nsew signal output
rlabel metal2 s 1122 59200 1178 60000 6 spi_err_i
port 419 nsew signal input
rlabel metal2 s 1674 59200 1730 60000 6 spi_rty_i
port 420 nsew signal input
rlabel metal2 s 4710 59200 4766 60000 6 spi_sel_o[0]
port 421 nsew signal output
rlabel metal2 s 6734 59200 6790 60000 6 spi_sel_o[1]
port 422 nsew signal output
rlabel metal2 s 8666 59200 8722 60000 6 spi_sel_o[2]
port 423 nsew signal output
rlabel metal2 s 10690 59200 10746 60000 6 spi_sel_o[3]
port 424 nsew signal output
rlabel metal2 s 2134 59200 2190 60000 6 spi_stb_o
port 425 nsew signal output
rlabel metal2 s 2686 59200 2742 60000 6 spi_we_o
port 426 nsew signal output
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 427 nsew power input
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 427 nsew power input
rlabel metal4 s 65648 2128 65968 57712 6 vccd1
port 427 nsew power input
rlabel metal4 s 96368 2128 96688 57712 6 vccd1
port 427 nsew power input
rlabel metal4 s 127088 2128 127408 57712 6 vccd1
port 427 nsew power input
rlabel metal4 s 157808 2128 158128 57712 6 vccd1
port 427 nsew power input
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 428 nsew ground input
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 428 nsew ground input
rlabel metal4 s 81008 2128 81328 57712 6 vssd1
port 428 nsew ground input
rlabel metal4 s 111728 2128 112048 57712 6 vssd1
port 428 nsew ground input
rlabel metal4 s 142448 2128 142768 57712 6 vssd1
port 428 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 160000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17939068
string GDS_FILE /home/q3k/sky130/qf105/openlane/mkQF100Fabric/runs/mkQF100Fabric/results/finishing/mkQF100Fabric.magic.gds
string GDS_START 912122
<< end >>

