VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mkQF100Fabric
  CLASS BLOCK ;
  FOREIGN mkQF100Fabric ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 300.000 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END CLK
  PIN RST_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END RST_N
  PIN cpu_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END cpu_ack_o
  PIN cpu_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END cpu_adr_i[0]
  PIN cpu_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END cpu_adr_i[10]
  PIN cpu_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END cpu_adr_i[11]
  PIN cpu_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END cpu_adr_i[12]
  PIN cpu_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END cpu_adr_i[13]
  PIN cpu_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END cpu_adr_i[14]
  PIN cpu_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END cpu_adr_i[15]
  PIN cpu_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END cpu_adr_i[16]
  PIN cpu_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
    END
  END cpu_adr_i[17]
  PIN cpu_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END cpu_adr_i[18]
  PIN cpu_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END cpu_adr_i[19]
  PIN cpu_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END cpu_adr_i[1]
  PIN cpu_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END cpu_adr_i[20]
  PIN cpu_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END cpu_adr_i[21]
  PIN cpu_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END cpu_adr_i[22]
  PIN cpu_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END cpu_adr_i[23]
  PIN cpu_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END cpu_adr_i[24]
  PIN cpu_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.800 4.000 243.400 ;
    END
  END cpu_adr_i[25]
  PIN cpu_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.960 4.000 251.560 ;
    END
  END cpu_adr_i[26]
  PIN cpu_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END cpu_adr_i[27]
  PIN cpu_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END cpu_adr_i[28]
  PIN cpu_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END cpu_adr_i[29]
  PIN cpu_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END cpu_adr_i[2]
  PIN cpu_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END cpu_adr_i[30]
  PIN cpu_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END cpu_adr_i[31]
  PIN cpu_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END cpu_adr_i[3]
  PIN cpu_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END cpu_adr_i[4]
  PIN cpu_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END cpu_adr_i[5]
  PIN cpu_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END cpu_adr_i[6]
  PIN cpu_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END cpu_adr_i[7]
  PIN cpu_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END cpu_adr_i[8]
  PIN cpu_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END cpu_adr_i[9]
  PIN cpu_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END cpu_cyc_i
  PIN cpu_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END cpu_dat_i[0]
  PIN cpu_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END cpu_dat_i[10]
  PIN cpu_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END cpu_dat_i[11]
  PIN cpu_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END cpu_dat_i[12]
  PIN cpu_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END cpu_dat_i[13]
  PIN cpu_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END cpu_dat_i[14]
  PIN cpu_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END cpu_dat_i[15]
  PIN cpu_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END cpu_dat_i[16]
  PIN cpu_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END cpu_dat_i[17]
  PIN cpu_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END cpu_dat_i[18]
  PIN cpu_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END cpu_dat_i[19]
  PIN cpu_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END cpu_dat_i[1]
  PIN cpu_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END cpu_dat_i[20]
  PIN cpu_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END cpu_dat_i[21]
  PIN cpu_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END cpu_dat_i[22]
  PIN cpu_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END cpu_dat_i[23]
  PIN cpu_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END cpu_dat_i[24]
  PIN cpu_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END cpu_dat_i[25]
  PIN cpu_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.680 4.000 254.280 ;
    END
  END cpu_dat_i[26]
  PIN cpu_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END cpu_dat_i[27]
  PIN cpu_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END cpu_dat_i[28]
  PIN cpu_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END cpu_dat_i[29]
  PIN cpu_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END cpu_dat_i[2]
  PIN cpu_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END cpu_dat_i[30]
  PIN cpu_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END cpu_dat_i[31]
  PIN cpu_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END cpu_dat_i[3]
  PIN cpu_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END cpu_dat_i[4]
  PIN cpu_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END cpu_dat_i[5]
  PIN cpu_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END cpu_dat_i[6]
  PIN cpu_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END cpu_dat_i[7]
  PIN cpu_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 4.000 104.680 ;
    END
  END cpu_dat_i[8]
  PIN cpu_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END cpu_dat_i[9]
  PIN cpu_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END cpu_dat_o[0]
  PIN cpu_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END cpu_dat_o[10]
  PIN cpu_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END cpu_dat_o[11]
  PIN cpu_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END cpu_dat_o[12]
  PIN cpu_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END cpu_dat_o[13]
  PIN cpu_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END cpu_dat_o[14]
  PIN cpu_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END cpu_dat_o[15]
  PIN cpu_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END cpu_dat_o[16]
  PIN cpu_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.600 4.000 182.200 ;
    END
  END cpu_dat_o[17]
  PIN cpu_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.760 4.000 190.360 ;
    END
  END cpu_dat_o[18]
  PIN cpu_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END cpu_dat_o[19]
  PIN cpu_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END cpu_dat_o[1]
  PIN cpu_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END cpu_dat_o[20]
  PIN cpu_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END cpu_dat_o[21]
  PIN cpu_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END cpu_dat_o[22]
  PIN cpu_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END cpu_dat_o[23]
  PIN cpu_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END cpu_dat_o[24]
  PIN cpu_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END cpu_dat_o[25]
  PIN cpu_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.400 4.000 257.000 ;
    END
  END cpu_dat_o[26]
  PIN cpu_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END cpu_dat_o[27]
  PIN cpu_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END cpu_dat_o[28]
  PIN cpu_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END cpu_dat_o[29]
  PIN cpu_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END cpu_dat_o[2]
  PIN cpu_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END cpu_dat_o[30]
  PIN cpu_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END cpu_dat_o[31]
  PIN cpu_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END cpu_dat_o[3]
  PIN cpu_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END cpu_dat_o[4]
  PIN cpu_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END cpu_dat_o[5]
  PIN cpu_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END cpu_dat_o[6]
  PIN cpu_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END cpu_dat_o[7]
  PIN cpu_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END cpu_dat_o[8]
  PIN cpu_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END cpu_dat_o[9]
  PIN cpu_err_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END cpu_err_o
  PIN cpu_rty_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END cpu_rty_o
  PIN cpu_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END cpu_sel_i[0]
  PIN cpu_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END cpu_sel_i[1]
  PIN cpu_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END cpu_sel_i[2]
  PIN cpu_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END cpu_sel_i[3]
  PIN cpu_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END cpu_stb_i
  PIN cpu_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END cpu_we_i
  PIN gpio_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 296.000 251.070 300.000 ;
    END
  END gpio_ack_i
  PIN gpio_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 296.000 265.330 300.000 ;
    END
  END gpio_adr_o[0]
  PIN gpio_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 296.000 345.370 300.000 ;
    END
  END gpio_adr_o[10]
  PIN gpio_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 296.000 352.270 300.000 ;
    END
  END gpio_adr_o[11]
  PIN gpio_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 296.000 359.630 300.000 ;
    END
  END gpio_adr_o[12]
  PIN gpio_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 296.000 366.530 300.000 ;
    END
  END gpio_adr_o[13]
  PIN gpio_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 296.000 373.890 300.000 ;
    END
  END gpio_adr_o[14]
  PIN gpio_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 296.000 380.790 300.000 ;
    END
  END gpio_adr_o[15]
  PIN gpio_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.410 296.000 387.690 300.000 ;
    END
  END gpio_adr_o[16]
  PIN gpio_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 296.000 395.050 300.000 ;
    END
  END gpio_adr_o[17]
  PIN gpio_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 296.000 401.950 300.000 ;
    END
  END gpio_adr_o[18]
  PIN gpio_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 296.000 409.310 300.000 ;
    END
  END gpio_adr_o[19]
  PIN gpio_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 296.000 274.530 300.000 ;
    END
  END gpio_adr_o[1]
  PIN gpio_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 296.000 416.210 300.000 ;
    END
  END gpio_adr_o[20]
  PIN gpio_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 296.000 423.110 300.000 ;
    END
  END gpio_adr_o[21]
  PIN gpio_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 296.000 430.470 300.000 ;
    END
  END gpio_adr_o[22]
  PIN gpio_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 296.000 437.370 300.000 ;
    END
  END gpio_adr_o[23]
  PIN gpio_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 296.000 444.270 300.000 ;
    END
  END gpio_adr_o[24]
  PIN gpio_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 296.000 451.630 300.000 ;
    END
  END gpio_adr_o[25]
  PIN gpio_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 296.000 458.530 300.000 ;
    END
  END gpio_adr_o[26]
  PIN gpio_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 296.000 465.890 300.000 ;
    END
  END gpio_adr_o[27]
  PIN gpio_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 296.000 472.790 300.000 ;
    END
  END gpio_adr_o[28]
  PIN gpio_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 296.000 479.690 300.000 ;
    END
  END gpio_adr_o[29]
  PIN gpio_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 296.000 284.190 300.000 ;
    END
  END gpio_adr_o[2]
  PIN gpio_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 296.000 487.050 300.000 ;
    END
  END gpio_adr_o[30]
  PIN gpio_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.670 296.000 493.950 300.000 ;
    END
  END gpio_adr_o[31]
  PIN gpio_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 296.000 293.390 300.000 ;
    END
  END gpio_adr_o[3]
  PIN gpio_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 296.000 303.050 300.000 ;
    END
  END gpio_adr_o[4]
  PIN gpio_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 296.000 309.950 300.000 ;
    END
  END gpio_adr_o[5]
  PIN gpio_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 296.000 317.310 300.000 ;
    END
  END gpio_adr_o[6]
  PIN gpio_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 296.000 324.210 300.000 ;
    END
  END gpio_adr_o[7]
  PIN gpio_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 296.000 331.110 300.000 ;
    END
  END gpio_adr_o[8]
  PIN gpio_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 296.000 338.470 300.000 ;
    END
  END gpio_adr_o[9]
  PIN gpio_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 296.000 253.370 300.000 ;
    END
  END gpio_cyc_o
  PIN gpio_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 296.000 267.630 300.000 ;
    END
  END gpio_dat_i[0]
  PIN gpio_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 296.000 347.670 300.000 ;
    END
  END gpio_dat_i[10]
  PIN gpio_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 296.000 355.030 300.000 ;
    END
  END gpio_dat_i[11]
  PIN gpio_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 296.000 361.930 300.000 ;
    END
  END gpio_dat_i[12]
  PIN gpio_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 296.000 368.830 300.000 ;
    END
  END gpio_dat_i[13]
  PIN gpio_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.910 296.000 376.190 300.000 ;
    END
  END gpio_dat_i[14]
  PIN gpio_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 296.000 383.090 300.000 ;
    END
  END gpio_dat_i[15]
  PIN gpio_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 296.000 390.450 300.000 ;
    END
  END gpio_dat_i[16]
  PIN gpio_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 296.000 397.350 300.000 ;
    END
  END gpio_dat_i[17]
  PIN gpio_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 296.000 404.250 300.000 ;
    END
  END gpio_dat_i[18]
  PIN gpio_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 296.000 411.610 300.000 ;
    END
  END gpio_dat_i[19]
  PIN gpio_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 296.000 276.830 300.000 ;
    END
  END gpio_dat_i[1]
  PIN gpio_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 296.000 418.510 300.000 ;
    END
  END gpio_dat_i[20]
  PIN gpio_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 296.000 425.410 300.000 ;
    END
  END gpio_dat_i[21]
  PIN gpio_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 296.000 432.770 300.000 ;
    END
  END gpio_dat_i[22]
  PIN gpio_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 296.000 439.670 300.000 ;
    END
  END gpio_dat_i[23]
  PIN gpio_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 296.000 447.030 300.000 ;
    END
  END gpio_dat_i[24]
  PIN gpio_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 296.000 453.930 300.000 ;
    END
  END gpio_dat_i[25]
  PIN gpio_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 296.000 460.830 300.000 ;
    END
  END gpio_dat_i[26]
  PIN gpio_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 296.000 468.190 300.000 ;
    END
  END gpio_dat_i[27]
  PIN gpio_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 296.000 475.090 300.000 ;
    END
  END gpio_dat_i[28]
  PIN gpio_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 296.000 481.990 300.000 ;
    END
  END gpio_dat_i[29]
  PIN gpio_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 296.000 286.490 300.000 ;
    END
  END gpio_dat_i[2]
  PIN gpio_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 296.000 489.350 300.000 ;
    END
  END gpio_dat_i[30]
  PIN gpio_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 296.000 496.250 300.000 ;
    END
  END gpio_dat_i[31]
  PIN gpio_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 296.000 295.690 300.000 ;
    END
  END gpio_dat_i[3]
  PIN gpio_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 296.000 305.350 300.000 ;
    END
  END gpio_dat_i[4]
  PIN gpio_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 296.000 312.250 300.000 ;
    END
  END gpio_dat_i[5]
  PIN gpio_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 296.000 319.610 300.000 ;
    END
  END gpio_dat_i[6]
  PIN gpio_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 296.000 326.510 300.000 ;
    END
  END gpio_dat_i[7]
  PIN gpio_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 296.000 333.410 300.000 ;
    END
  END gpio_dat_i[8]
  PIN gpio_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 296.000 340.770 300.000 ;
    END
  END gpio_dat_i[9]
  PIN gpio_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 296.000 269.930 300.000 ;
    END
  END gpio_dat_o[0]
  PIN gpio_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 296.000 349.970 300.000 ;
    END
  END gpio_dat_o[10]
  PIN gpio_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 296.000 357.330 300.000 ;
    END
  END gpio_dat_o[11]
  PIN gpio_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 296.000 364.230 300.000 ;
    END
  END gpio_dat_o[12]
  PIN gpio_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 296.000 371.130 300.000 ;
    END
  END gpio_dat_o[13]
  PIN gpio_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 296.000 378.490 300.000 ;
    END
  END gpio_dat_o[14]
  PIN gpio_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 296.000 385.390 300.000 ;
    END
  END gpio_dat_o[15]
  PIN gpio_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 296.000 392.750 300.000 ;
    END
  END gpio_dat_o[16]
  PIN gpio_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 296.000 399.650 300.000 ;
    END
  END gpio_dat_o[17]
  PIN gpio_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 296.000 406.550 300.000 ;
    END
  END gpio_dat_o[18]
  PIN gpio_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 296.000 413.910 300.000 ;
    END
  END gpio_dat_o[19]
  PIN gpio_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 296.000 279.590 300.000 ;
    END
  END gpio_dat_o[1]
  PIN gpio_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 296.000 420.810 300.000 ;
    END
  END gpio_dat_o[20]
  PIN gpio_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 296.000 428.170 300.000 ;
    END
  END gpio_dat_o[21]
  PIN gpio_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 296.000 435.070 300.000 ;
    END
  END gpio_dat_o[22]
  PIN gpio_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 296.000 441.970 300.000 ;
    END
  END gpio_dat_o[23]
  PIN gpio_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 296.000 449.330 300.000 ;
    END
  END gpio_dat_o[24]
  PIN gpio_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 296.000 456.230 300.000 ;
    END
  END gpio_dat_o[25]
  PIN gpio_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 296.000 463.130 300.000 ;
    END
  END gpio_dat_o[26]
  PIN gpio_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 296.000 470.490 300.000 ;
    END
  END gpio_dat_o[27]
  PIN gpio_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 296.000 477.390 300.000 ;
    END
  END gpio_dat_o[28]
  PIN gpio_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 296.000 484.750 300.000 ;
    END
  END gpio_dat_o[29]
  PIN gpio_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 296.000 288.790 300.000 ;
    END
  END gpio_dat_o[2]
  PIN gpio_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 296.000 491.650 300.000 ;
    END
  END gpio_dat_o[30]
  PIN gpio_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.270 296.000 498.550 300.000 ;
    END
  END gpio_dat_o[31]
  PIN gpio_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 296.000 298.450 300.000 ;
    END
  END gpio_dat_o[3]
  PIN gpio_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 296.000 307.650 300.000 ;
    END
  END gpio_dat_o[4]
  PIN gpio_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 296.000 314.550 300.000 ;
    END
  END gpio_dat_o[5]
  PIN gpio_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 296.000 321.910 300.000 ;
    END
  END gpio_dat_o[6]
  PIN gpio_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 296.000 328.810 300.000 ;
    END
  END gpio_dat_o[7]
  PIN gpio_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 296.000 336.170 300.000 ;
    END
  END gpio_dat_o[8]
  PIN gpio_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 296.000 343.070 300.000 ;
    END
  END gpio_dat_o[9]
  PIN gpio_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 296.000 255.670 300.000 ;
    END
  END gpio_err_i
  PIN gpio_rty_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 296.000 257.970 300.000 ;
    END
  END gpio_rty_i
  PIN gpio_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 296.000 272.230 300.000 ;
    END
  END gpio_sel_o[0]
  PIN gpio_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 296.000 281.890 300.000 ;
    END
  END gpio_sel_o[1]
  PIN gpio_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 296.000 291.090 300.000 ;
    END
  END gpio_sel_o[2]
  PIN gpio_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 296.000 300.750 300.000 ;
    END
  END gpio_sel_o[3]
  PIN gpio_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 296.000 260.730 300.000 ;
    END
  END gpio_stb_o
  PIN gpio_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 296.000 263.030 300.000 ;
    END
  END gpio_we_o
  PIN spi_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 296.000 1.290 300.000 ;
    END
  END spi_ack_i
  PIN spi_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 296.000 15.090 300.000 ;
    END
  END spi_adr_o[0]
  PIN spi_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 296.000 95.590 300.000 ;
    END
  END spi_adr_o[10]
  PIN spi_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 296.000 102.490 300.000 ;
    END
  END spi_adr_o[11]
  PIN spi_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 296.000 109.390 300.000 ;
    END
  END spi_adr_o[12]
  PIN spi_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 296.000 116.750 300.000 ;
    END
  END spi_adr_o[13]
  PIN spi_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 296.000 123.650 300.000 ;
    END
  END spi_adr_o[14]
  PIN spi_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 296.000 131.010 300.000 ;
    END
  END spi_adr_o[15]
  PIN spi_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 296.000 137.910 300.000 ;
    END
  END spi_adr_o[16]
  PIN spi_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 296.000 144.810 300.000 ;
    END
  END spi_adr_o[17]
  PIN spi_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 296.000 152.170 300.000 ;
    END
  END spi_adr_o[18]
  PIN spi_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 296.000 159.070 300.000 ;
    END
  END spi_adr_o[19]
  PIN spi_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 296.000 24.750 300.000 ;
    END
  END spi_adr_o[1]
  PIN spi_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 296.000 165.970 300.000 ;
    END
  END spi_adr_o[20]
  PIN spi_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 296.000 173.330 300.000 ;
    END
  END spi_adr_o[21]
  PIN spi_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 296.000 180.230 300.000 ;
    END
  END spi_adr_o[22]
  PIN spi_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 296.000 187.590 300.000 ;
    END
  END spi_adr_o[23]
  PIN spi_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 296.000 194.490 300.000 ;
    END
  END spi_adr_o[24]
  PIN spi_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 296.000 201.390 300.000 ;
    END
  END spi_adr_o[25]
  PIN spi_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 296.000 208.750 300.000 ;
    END
  END spi_adr_o[26]
  PIN spi_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 296.000 215.650 300.000 ;
    END
  END spi_adr_o[27]
  PIN spi_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 296.000 222.550 300.000 ;
    END
  END spi_adr_o[28]
  PIN spi_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 296.000 229.910 300.000 ;
    END
  END spi_adr_o[29]
  PIN spi_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 296.000 33.950 300.000 ;
    END
  END spi_adr_o[2]
  PIN spi_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 296.000 236.810 300.000 ;
    END
  END spi_adr_o[30]
  PIN spi_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 296.000 244.170 300.000 ;
    END
  END spi_adr_o[31]
  PIN spi_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 296.000 43.610 300.000 ;
    END
  END spi_adr_o[3]
  PIN spi_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 296.000 52.810 300.000 ;
    END
  END spi_adr_o[4]
  PIN spi_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 296.000 60.170 300.000 ;
    END
  END spi_adr_o[5]
  PIN spi_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 296.000 67.070 300.000 ;
    END
  END spi_adr_o[6]
  PIN spi_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 296.000 73.970 300.000 ;
    END
  END spi_adr_o[7]
  PIN spi_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 296.000 81.330 300.000 ;
    END
  END spi_adr_o[8]
  PIN spi_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 296.000 88.230 300.000 ;
    END
  END spi_adr_o[9]
  PIN spi_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 296.000 3.590 300.000 ;
    END
  END spi_cyc_o
  PIN spi_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 296.000 17.390 300.000 ;
    END
  END spi_dat_i[0]
  PIN spi_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 296.000 97.890 300.000 ;
    END
  END spi_dat_i[10]
  PIN spi_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 296.000 104.790 300.000 ;
    END
  END spi_dat_i[11]
  PIN spi_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 296.000 111.690 300.000 ;
    END
  END spi_dat_i[12]
  PIN spi_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 296.000 119.050 300.000 ;
    END
  END spi_dat_i[13]
  PIN spi_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 296.000 125.950 300.000 ;
    END
  END spi_dat_i[14]
  PIN spi_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 296.000 133.310 300.000 ;
    END
  END spi_dat_i[15]
  PIN spi_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 296.000 140.210 300.000 ;
    END
  END spi_dat_i[16]
  PIN spi_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 296.000 147.110 300.000 ;
    END
  END spi_dat_i[17]
  PIN spi_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 296.000 154.470 300.000 ;
    END
  END spi_dat_i[18]
  PIN spi_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 296.000 161.370 300.000 ;
    END
  END spi_dat_i[19]
  PIN spi_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 296.000 27.050 300.000 ;
    END
  END spi_dat_i[1]
  PIN spi_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 296.000 168.730 300.000 ;
    END
  END spi_dat_i[20]
  PIN spi_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 296.000 175.630 300.000 ;
    END
  END spi_dat_i[21]
  PIN spi_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 296.000 182.530 300.000 ;
    END
  END spi_dat_i[22]
  PIN spi_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 296.000 189.890 300.000 ;
    END
  END spi_dat_i[23]
  PIN spi_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 296.000 196.790 300.000 ;
    END
  END spi_dat_i[24]
  PIN spi_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 296.000 203.690 300.000 ;
    END
  END spi_dat_i[25]
  PIN spi_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 296.000 211.050 300.000 ;
    END
  END spi_dat_i[26]
  PIN spi_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 296.000 217.950 300.000 ;
    END
  END spi_dat_i[27]
  PIN spi_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 296.000 225.310 300.000 ;
    END
  END spi_dat_i[28]
  PIN spi_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 296.000 232.210 300.000 ;
    END
  END spi_dat_i[29]
  PIN spi_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 296.000 36.250 300.000 ;
    END
  END spi_dat_i[2]
  PIN spi_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 296.000 239.110 300.000 ;
    END
  END spi_dat_i[30]
  PIN spi_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 296.000 246.470 300.000 ;
    END
  END spi_dat_i[31]
  PIN spi_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 296.000 45.910 300.000 ;
    END
  END spi_dat_i[3]
  PIN spi_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 296.000 55.110 300.000 ;
    END
  END spi_dat_i[4]
  PIN spi_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 296.000 62.470 300.000 ;
    END
  END spi_dat_i[5]
  PIN spi_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 296.000 69.370 300.000 ;
    END
  END spi_dat_i[6]
  PIN spi_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 296.000 76.730 300.000 ;
    END
  END spi_dat_i[7]
  PIN spi_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 296.000 83.630 300.000 ;
    END
  END spi_dat_i[8]
  PIN spi_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 296.000 90.530 300.000 ;
    END
  END spi_dat_i[9]
  PIN spi_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 296.000 20.150 300.000 ;
    END
  END spi_dat_o[0]
  PIN spi_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 296.000 100.190 300.000 ;
    END
  END spi_dat_o[10]
  PIN spi_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 296.000 107.090 300.000 ;
    END
  END spi_dat_o[11]
  PIN spi_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 296.000 114.450 300.000 ;
    END
  END spi_dat_o[12]
  PIN spi_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 296.000 121.350 300.000 ;
    END
  END spi_dat_o[13]
  PIN spi_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 296.000 128.250 300.000 ;
    END
  END spi_dat_o[14]
  PIN spi_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 296.000 135.610 300.000 ;
    END
  END spi_dat_o[15]
  PIN spi_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 296.000 142.510 300.000 ;
    END
  END spi_dat_o[16]
  PIN spi_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 296.000 149.870 300.000 ;
    END
  END spi_dat_o[17]
  PIN spi_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 296.000 156.770 300.000 ;
    END
  END spi_dat_o[18]
  PIN spi_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 296.000 163.670 300.000 ;
    END
  END spi_dat_o[19]
  PIN spi_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 296.000 29.350 300.000 ;
    END
  END spi_dat_o[1]
  PIN spi_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 296.000 171.030 300.000 ;
    END
  END spi_dat_o[20]
  PIN spi_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 296.000 177.930 300.000 ;
    END
  END spi_dat_o[21]
  PIN spi_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 296.000 184.830 300.000 ;
    END
  END spi_dat_o[22]
  PIN spi_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 296.000 192.190 300.000 ;
    END
  END spi_dat_o[23]
  PIN spi_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 296.000 199.090 300.000 ;
    END
  END spi_dat_o[24]
  PIN spi_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 296.000 206.450 300.000 ;
    END
  END spi_dat_o[25]
  PIN spi_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 296.000 213.350 300.000 ;
    END
  END spi_dat_o[26]
  PIN spi_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 296.000 220.250 300.000 ;
    END
  END spi_dat_o[27]
  PIN spi_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 296.000 227.610 300.000 ;
    END
  END spi_dat_o[28]
  PIN spi_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 296.000 234.510 300.000 ;
    END
  END spi_dat_o[29]
  PIN spi_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 296.000 39.010 300.000 ;
    END
  END spi_dat_o[2]
  PIN spi_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 296.000 241.410 300.000 ;
    END
  END spi_dat_o[30]
  PIN spi_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 296.000 248.770 300.000 ;
    END
  END spi_dat_o[31]
  PIN spi_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 296.000 48.210 300.000 ;
    END
  END spi_dat_o[3]
  PIN spi_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 296.000 57.870 300.000 ;
    END
  END spi_dat_o[4]
  PIN spi_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 296.000 64.770 300.000 ;
    END
  END spi_dat_o[5]
  PIN spi_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 296.000 71.670 300.000 ;
    END
  END spi_dat_o[6]
  PIN spi_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 296.000 79.030 300.000 ;
    END
  END spi_dat_o[7]
  PIN spi_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 296.000 85.930 300.000 ;
    END
  END spi_dat_o[8]
  PIN spi_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 296.000 92.830 300.000 ;
    END
  END spi_dat_o[9]
  PIN spi_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 296.000 5.890 300.000 ;
    END
  END spi_err_i
  PIN spi_rty_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 296.000 8.190 300.000 ;
    END
  END spi_rty_i
  PIN spi_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 296.000 22.450 300.000 ;
    END
  END spi_sel_o[0]
  PIN spi_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 296.000 31.650 300.000 ;
    END
  END spi_sel_o[1]
  PIN spi_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 296.000 41.310 300.000 ;
    END
  END spi_sel_o[2]
  PIN spi_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 296.000 50.510 300.000 ;
    END
  END spi_sel_o[3]
  PIN spi_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 296.000 10.490 300.000 ;
    END
  END spi_stb_o
  PIN spi_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 296.000 12.790 300.000 ;
    END
  END spi_we_o
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 288.560 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 288.405 ;
      LAYER met1 ;
        RECT 0.990 6.500 498.570 291.000 ;
      LAYER met2 ;
        RECT 1.570 295.720 3.030 298.365 ;
        RECT 3.870 295.720 5.330 298.365 ;
        RECT 6.170 295.720 7.630 298.365 ;
        RECT 8.470 295.720 9.930 298.365 ;
        RECT 10.770 295.720 12.230 298.365 ;
        RECT 13.070 295.720 14.530 298.365 ;
        RECT 15.370 295.720 16.830 298.365 ;
        RECT 17.670 295.720 19.590 298.365 ;
        RECT 20.430 295.720 21.890 298.365 ;
        RECT 22.730 295.720 24.190 298.365 ;
        RECT 25.030 295.720 26.490 298.365 ;
        RECT 27.330 295.720 28.790 298.365 ;
        RECT 29.630 295.720 31.090 298.365 ;
        RECT 31.930 295.720 33.390 298.365 ;
        RECT 34.230 295.720 35.690 298.365 ;
        RECT 36.530 295.720 38.450 298.365 ;
        RECT 39.290 295.720 40.750 298.365 ;
        RECT 41.590 295.720 43.050 298.365 ;
        RECT 43.890 295.720 45.350 298.365 ;
        RECT 46.190 295.720 47.650 298.365 ;
        RECT 48.490 295.720 49.950 298.365 ;
        RECT 50.790 295.720 52.250 298.365 ;
        RECT 53.090 295.720 54.550 298.365 ;
        RECT 55.390 295.720 57.310 298.365 ;
        RECT 58.150 295.720 59.610 298.365 ;
        RECT 60.450 295.720 61.910 298.365 ;
        RECT 62.750 295.720 64.210 298.365 ;
        RECT 65.050 295.720 66.510 298.365 ;
        RECT 67.350 295.720 68.810 298.365 ;
        RECT 69.650 295.720 71.110 298.365 ;
        RECT 71.950 295.720 73.410 298.365 ;
        RECT 74.250 295.720 76.170 298.365 ;
        RECT 77.010 295.720 78.470 298.365 ;
        RECT 79.310 295.720 80.770 298.365 ;
        RECT 81.610 295.720 83.070 298.365 ;
        RECT 83.910 295.720 85.370 298.365 ;
        RECT 86.210 295.720 87.670 298.365 ;
        RECT 88.510 295.720 89.970 298.365 ;
        RECT 90.810 295.720 92.270 298.365 ;
        RECT 93.110 295.720 95.030 298.365 ;
        RECT 95.870 295.720 97.330 298.365 ;
        RECT 98.170 295.720 99.630 298.365 ;
        RECT 100.470 295.720 101.930 298.365 ;
        RECT 102.770 295.720 104.230 298.365 ;
        RECT 105.070 295.720 106.530 298.365 ;
        RECT 107.370 295.720 108.830 298.365 ;
        RECT 109.670 295.720 111.130 298.365 ;
        RECT 111.970 295.720 113.890 298.365 ;
        RECT 114.730 295.720 116.190 298.365 ;
        RECT 117.030 295.720 118.490 298.365 ;
        RECT 119.330 295.720 120.790 298.365 ;
        RECT 121.630 295.720 123.090 298.365 ;
        RECT 123.930 295.720 125.390 298.365 ;
        RECT 126.230 295.720 127.690 298.365 ;
        RECT 128.530 295.720 130.450 298.365 ;
        RECT 131.290 295.720 132.750 298.365 ;
        RECT 133.590 295.720 135.050 298.365 ;
        RECT 135.890 295.720 137.350 298.365 ;
        RECT 138.190 295.720 139.650 298.365 ;
        RECT 140.490 295.720 141.950 298.365 ;
        RECT 142.790 295.720 144.250 298.365 ;
        RECT 145.090 295.720 146.550 298.365 ;
        RECT 147.390 295.720 149.310 298.365 ;
        RECT 150.150 295.720 151.610 298.365 ;
        RECT 152.450 295.720 153.910 298.365 ;
        RECT 154.750 295.720 156.210 298.365 ;
        RECT 157.050 295.720 158.510 298.365 ;
        RECT 159.350 295.720 160.810 298.365 ;
        RECT 161.650 295.720 163.110 298.365 ;
        RECT 163.950 295.720 165.410 298.365 ;
        RECT 166.250 295.720 168.170 298.365 ;
        RECT 169.010 295.720 170.470 298.365 ;
        RECT 171.310 295.720 172.770 298.365 ;
        RECT 173.610 295.720 175.070 298.365 ;
        RECT 175.910 295.720 177.370 298.365 ;
        RECT 178.210 295.720 179.670 298.365 ;
        RECT 180.510 295.720 181.970 298.365 ;
        RECT 182.810 295.720 184.270 298.365 ;
        RECT 185.110 295.720 187.030 298.365 ;
        RECT 187.870 295.720 189.330 298.365 ;
        RECT 190.170 295.720 191.630 298.365 ;
        RECT 192.470 295.720 193.930 298.365 ;
        RECT 194.770 295.720 196.230 298.365 ;
        RECT 197.070 295.720 198.530 298.365 ;
        RECT 199.370 295.720 200.830 298.365 ;
        RECT 201.670 295.720 203.130 298.365 ;
        RECT 203.970 295.720 205.890 298.365 ;
        RECT 206.730 295.720 208.190 298.365 ;
        RECT 209.030 295.720 210.490 298.365 ;
        RECT 211.330 295.720 212.790 298.365 ;
        RECT 213.630 295.720 215.090 298.365 ;
        RECT 215.930 295.720 217.390 298.365 ;
        RECT 218.230 295.720 219.690 298.365 ;
        RECT 220.530 295.720 221.990 298.365 ;
        RECT 222.830 295.720 224.750 298.365 ;
        RECT 225.590 295.720 227.050 298.365 ;
        RECT 227.890 295.720 229.350 298.365 ;
        RECT 230.190 295.720 231.650 298.365 ;
        RECT 232.490 295.720 233.950 298.365 ;
        RECT 234.790 295.720 236.250 298.365 ;
        RECT 237.090 295.720 238.550 298.365 ;
        RECT 239.390 295.720 240.850 298.365 ;
        RECT 241.690 295.720 243.610 298.365 ;
        RECT 244.450 295.720 245.910 298.365 ;
        RECT 246.750 295.720 248.210 298.365 ;
        RECT 249.050 295.720 250.510 298.365 ;
        RECT 251.350 295.720 252.810 298.365 ;
        RECT 253.650 295.720 255.110 298.365 ;
        RECT 255.950 295.720 257.410 298.365 ;
        RECT 258.250 295.720 260.170 298.365 ;
        RECT 261.010 295.720 262.470 298.365 ;
        RECT 263.310 295.720 264.770 298.365 ;
        RECT 265.610 295.720 267.070 298.365 ;
        RECT 267.910 295.720 269.370 298.365 ;
        RECT 270.210 295.720 271.670 298.365 ;
        RECT 272.510 295.720 273.970 298.365 ;
        RECT 274.810 295.720 276.270 298.365 ;
        RECT 277.110 295.720 279.030 298.365 ;
        RECT 279.870 295.720 281.330 298.365 ;
        RECT 282.170 295.720 283.630 298.365 ;
        RECT 284.470 295.720 285.930 298.365 ;
        RECT 286.770 295.720 288.230 298.365 ;
        RECT 289.070 295.720 290.530 298.365 ;
        RECT 291.370 295.720 292.830 298.365 ;
        RECT 293.670 295.720 295.130 298.365 ;
        RECT 295.970 295.720 297.890 298.365 ;
        RECT 298.730 295.720 300.190 298.365 ;
        RECT 301.030 295.720 302.490 298.365 ;
        RECT 303.330 295.720 304.790 298.365 ;
        RECT 305.630 295.720 307.090 298.365 ;
        RECT 307.930 295.720 309.390 298.365 ;
        RECT 310.230 295.720 311.690 298.365 ;
        RECT 312.530 295.720 313.990 298.365 ;
        RECT 314.830 295.720 316.750 298.365 ;
        RECT 317.590 295.720 319.050 298.365 ;
        RECT 319.890 295.720 321.350 298.365 ;
        RECT 322.190 295.720 323.650 298.365 ;
        RECT 324.490 295.720 325.950 298.365 ;
        RECT 326.790 295.720 328.250 298.365 ;
        RECT 329.090 295.720 330.550 298.365 ;
        RECT 331.390 295.720 332.850 298.365 ;
        RECT 333.690 295.720 335.610 298.365 ;
        RECT 336.450 295.720 337.910 298.365 ;
        RECT 338.750 295.720 340.210 298.365 ;
        RECT 341.050 295.720 342.510 298.365 ;
        RECT 343.350 295.720 344.810 298.365 ;
        RECT 345.650 295.720 347.110 298.365 ;
        RECT 347.950 295.720 349.410 298.365 ;
        RECT 350.250 295.720 351.710 298.365 ;
        RECT 352.550 295.720 354.470 298.365 ;
        RECT 355.310 295.720 356.770 298.365 ;
        RECT 357.610 295.720 359.070 298.365 ;
        RECT 359.910 295.720 361.370 298.365 ;
        RECT 362.210 295.720 363.670 298.365 ;
        RECT 364.510 295.720 365.970 298.365 ;
        RECT 366.810 295.720 368.270 298.365 ;
        RECT 369.110 295.720 370.570 298.365 ;
        RECT 371.410 295.720 373.330 298.365 ;
        RECT 374.170 295.720 375.630 298.365 ;
        RECT 376.470 295.720 377.930 298.365 ;
        RECT 378.770 295.720 380.230 298.365 ;
        RECT 381.070 295.720 382.530 298.365 ;
        RECT 383.370 295.720 384.830 298.365 ;
        RECT 385.670 295.720 387.130 298.365 ;
        RECT 387.970 295.720 389.890 298.365 ;
        RECT 390.730 295.720 392.190 298.365 ;
        RECT 393.030 295.720 394.490 298.365 ;
        RECT 395.330 295.720 396.790 298.365 ;
        RECT 397.630 295.720 399.090 298.365 ;
        RECT 399.930 295.720 401.390 298.365 ;
        RECT 402.230 295.720 403.690 298.365 ;
        RECT 404.530 295.720 405.990 298.365 ;
        RECT 406.830 295.720 408.750 298.365 ;
        RECT 409.590 295.720 411.050 298.365 ;
        RECT 411.890 295.720 413.350 298.365 ;
        RECT 414.190 295.720 415.650 298.365 ;
        RECT 416.490 295.720 417.950 298.365 ;
        RECT 418.790 295.720 420.250 298.365 ;
        RECT 421.090 295.720 422.550 298.365 ;
        RECT 423.390 295.720 424.850 298.365 ;
        RECT 425.690 295.720 427.610 298.365 ;
        RECT 428.450 295.720 429.910 298.365 ;
        RECT 430.750 295.720 432.210 298.365 ;
        RECT 433.050 295.720 434.510 298.365 ;
        RECT 435.350 295.720 436.810 298.365 ;
        RECT 437.650 295.720 439.110 298.365 ;
        RECT 439.950 295.720 441.410 298.365 ;
        RECT 442.250 295.720 443.710 298.365 ;
        RECT 444.550 295.720 446.470 298.365 ;
        RECT 447.310 295.720 448.770 298.365 ;
        RECT 449.610 295.720 451.070 298.365 ;
        RECT 451.910 295.720 453.370 298.365 ;
        RECT 454.210 295.720 455.670 298.365 ;
        RECT 456.510 295.720 457.970 298.365 ;
        RECT 458.810 295.720 460.270 298.365 ;
        RECT 461.110 295.720 462.570 298.365 ;
        RECT 463.410 295.720 465.330 298.365 ;
        RECT 466.170 295.720 467.630 298.365 ;
        RECT 468.470 295.720 469.930 298.365 ;
        RECT 470.770 295.720 472.230 298.365 ;
        RECT 473.070 295.720 474.530 298.365 ;
        RECT 475.370 295.720 476.830 298.365 ;
        RECT 477.670 295.720 479.130 298.365 ;
        RECT 479.970 295.720 481.430 298.365 ;
        RECT 482.270 295.720 484.190 298.365 ;
        RECT 485.030 295.720 486.490 298.365 ;
        RECT 487.330 295.720 488.790 298.365 ;
        RECT 489.630 295.720 491.090 298.365 ;
        RECT 491.930 295.720 493.390 298.365 ;
        RECT 494.230 295.720 495.690 298.365 ;
        RECT 496.530 295.720 497.990 298.365 ;
        RECT 1.020 1.515 498.540 295.720 ;
      LAYER met3 ;
        RECT 4.400 297.480 489.835 298.345 ;
        RECT 4.000 296.160 489.835 297.480 ;
        RECT 4.400 294.760 489.835 296.160 ;
        RECT 4.000 293.440 489.835 294.760 ;
        RECT 4.400 292.040 489.835 293.440 ;
        RECT 4.000 290.720 489.835 292.040 ;
        RECT 4.400 289.320 489.835 290.720 ;
        RECT 4.000 288.000 489.835 289.320 ;
        RECT 4.400 286.600 489.835 288.000 ;
        RECT 4.000 285.280 489.835 286.600 ;
        RECT 4.400 283.880 489.835 285.280 ;
        RECT 4.000 282.560 489.835 283.880 ;
        RECT 4.400 281.160 489.835 282.560 ;
        RECT 4.000 279.840 489.835 281.160 ;
        RECT 4.400 278.440 489.835 279.840 ;
        RECT 4.000 277.120 489.835 278.440 ;
        RECT 4.400 275.720 489.835 277.120 ;
        RECT 4.000 274.400 489.835 275.720 ;
        RECT 4.400 273.000 489.835 274.400 ;
        RECT 4.000 271.680 489.835 273.000 ;
        RECT 4.400 270.280 489.835 271.680 ;
        RECT 4.000 268.960 489.835 270.280 ;
        RECT 4.400 267.560 489.835 268.960 ;
        RECT 4.000 265.560 489.835 267.560 ;
        RECT 4.400 264.160 489.835 265.560 ;
        RECT 4.000 262.840 489.835 264.160 ;
        RECT 4.400 261.440 489.835 262.840 ;
        RECT 4.000 260.120 489.835 261.440 ;
        RECT 4.400 258.720 489.835 260.120 ;
        RECT 4.000 257.400 489.835 258.720 ;
        RECT 4.400 256.000 489.835 257.400 ;
        RECT 4.000 254.680 489.835 256.000 ;
        RECT 4.400 253.280 489.835 254.680 ;
        RECT 4.000 251.960 489.835 253.280 ;
        RECT 4.400 250.560 489.835 251.960 ;
        RECT 4.000 249.240 489.835 250.560 ;
        RECT 4.400 247.840 489.835 249.240 ;
        RECT 4.000 246.520 489.835 247.840 ;
        RECT 4.400 245.120 489.835 246.520 ;
        RECT 4.000 243.800 489.835 245.120 ;
        RECT 4.400 242.400 489.835 243.800 ;
        RECT 4.000 241.080 489.835 242.400 ;
        RECT 4.400 239.680 489.835 241.080 ;
        RECT 4.000 238.360 489.835 239.680 ;
        RECT 4.400 236.960 489.835 238.360 ;
        RECT 4.000 235.640 489.835 236.960 ;
        RECT 4.400 234.240 489.835 235.640 ;
        RECT 4.000 232.240 489.835 234.240 ;
        RECT 4.400 230.840 489.835 232.240 ;
        RECT 4.000 229.520 489.835 230.840 ;
        RECT 4.400 228.120 489.835 229.520 ;
        RECT 4.000 226.800 489.835 228.120 ;
        RECT 4.400 225.400 489.835 226.800 ;
        RECT 4.000 224.080 489.835 225.400 ;
        RECT 4.400 222.680 489.835 224.080 ;
        RECT 4.000 221.360 489.835 222.680 ;
        RECT 4.400 219.960 489.835 221.360 ;
        RECT 4.000 218.640 489.835 219.960 ;
        RECT 4.400 217.240 489.835 218.640 ;
        RECT 4.000 215.920 489.835 217.240 ;
        RECT 4.400 214.520 489.835 215.920 ;
        RECT 4.000 213.200 489.835 214.520 ;
        RECT 4.400 211.800 489.835 213.200 ;
        RECT 4.000 210.480 489.835 211.800 ;
        RECT 4.400 209.080 489.835 210.480 ;
        RECT 4.000 207.760 489.835 209.080 ;
        RECT 4.400 206.360 489.835 207.760 ;
        RECT 4.000 205.040 489.835 206.360 ;
        RECT 4.400 203.640 489.835 205.040 ;
        RECT 4.000 202.320 489.835 203.640 ;
        RECT 4.400 200.920 489.835 202.320 ;
        RECT 4.000 198.920 489.835 200.920 ;
        RECT 4.400 197.520 489.835 198.920 ;
        RECT 4.000 196.200 489.835 197.520 ;
        RECT 4.400 194.800 489.835 196.200 ;
        RECT 4.000 193.480 489.835 194.800 ;
        RECT 4.400 192.080 489.835 193.480 ;
        RECT 4.000 190.760 489.835 192.080 ;
        RECT 4.400 189.360 489.835 190.760 ;
        RECT 4.000 188.040 489.835 189.360 ;
        RECT 4.400 186.640 489.835 188.040 ;
        RECT 4.000 185.320 489.835 186.640 ;
        RECT 4.400 183.920 489.835 185.320 ;
        RECT 4.000 182.600 489.835 183.920 ;
        RECT 4.400 181.200 489.835 182.600 ;
        RECT 4.000 179.880 489.835 181.200 ;
        RECT 4.400 178.480 489.835 179.880 ;
        RECT 4.000 177.160 489.835 178.480 ;
        RECT 4.400 175.760 489.835 177.160 ;
        RECT 4.000 174.440 489.835 175.760 ;
        RECT 4.400 173.040 489.835 174.440 ;
        RECT 4.000 171.720 489.835 173.040 ;
        RECT 4.400 170.320 489.835 171.720 ;
        RECT 4.000 169.000 489.835 170.320 ;
        RECT 4.400 167.600 489.835 169.000 ;
        RECT 4.000 165.600 489.835 167.600 ;
        RECT 4.400 164.200 489.835 165.600 ;
        RECT 4.000 162.880 489.835 164.200 ;
        RECT 4.400 161.480 489.835 162.880 ;
        RECT 4.000 160.160 489.835 161.480 ;
        RECT 4.400 158.760 489.835 160.160 ;
        RECT 4.000 157.440 489.835 158.760 ;
        RECT 4.400 156.040 489.835 157.440 ;
        RECT 4.000 154.720 489.835 156.040 ;
        RECT 4.400 153.320 489.835 154.720 ;
        RECT 4.000 152.000 489.835 153.320 ;
        RECT 4.400 150.600 489.835 152.000 ;
        RECT 4.000 149.280 489.835 150.600 ;
        RECT 4.400 147.880 489.835 149.280 ;
        RECT 4.000 146.560 489.835 147.880 ;
        RECT 4.400 145.160 489.835 146.560 ;
        RECT 4.000 143.840 489.835 145.160 ;
        RECT 4.400 142.440 489.835 143.840 ;
        RECT 4.000 141.120 489.835 142.440 ;
        RECT 4.400 139.720 489.835 141.120 ;
        RECT 4.000 138.400 489.835 139.720 ;
        RECT 4.400 137.000 489.835 138.400 ;
        RECT 4.000 135.680 489.835 137.000 ;
        RECT 4.400 134.280 489.835 135.680 ;
        RECT 4.000 132.280 489.835 134.280 ;
        RECT 4.400 130.880 489.835 132.280 ;
        RECT 4.000 129.560 489.835 130.880 ;
        RECT 4.400 128.160 489.835 129.560 ;
        RECT 4.000 126.840 489.835 128.160 ;
        RECT 4.400 125.440 489.835 126.840 ;
        RECT 4.000 124.120 489.835 125.440 ;
        RECT 4.400 122.720 489.835 124.120 ;
        RECT 4.000 121.400 489.835 122.720 ;
        RECT 4.400 120.000 489.835 121.400 ;
        RECT 4.000 118.680 489.835 120.000 ;
        RECT 4.400 117.280 489.835 118.680 ;
        RECT 4.000 115.960 489.835 117.280 ;
        RECT 4.400 114.560 489.835 115.960 ;
        RECT 4.000 113.240 489.835 114.560 ;
        RECT 4.400 111.840 489.835 113.240 ;
        RECT 4.000 110.520 489.835 111.840 ;
        RECT 4.400 109.120 489.835 110.520 ;
        RECT 4.000 107.800 489.835 109.120 ;
        RECT 4.400 106.400 489.835 107.800 ;
        RECT 4.000 105.080 489.835 106.400 ;
        RECT 4.400 103.680 489.835 105.080 ;
        RECT 4.000 102.360 489.835 103.680 ;
        RECT 4.400 100.960 489.835 102.360 ;
        RECT 4.000 98.960 489.835 100.960 ;
        RECT 4.400 97.560 489.835 98.960 ;
        RECT 4.000 96.240 489.835 97.560 ;
        RECT 4.400 94.840 489.835 96.240 ;
        RECT 4.000 93.520 489.835 94.840 ;
        RECT 4.400 92.120 489.835 93.520 ;
        RECT 4.000 90.800 489.835 92.120 ;
        RECT 4.400 89.400 489.835 90.800 ;
        RECT 4.000 88.080 489.835 89.400 ;
        RECT 4.400 86.680 489.835 88.080 ;
        RECT 4.000 85.360 489.835 86.680 ;
        RECT 4.400 83.960 489.835 85.360 ;
        RECT 4.000 82.640 489.835 83.960 ;
        RECT 4.400 81.240 489.835 82.640 ;
        RECT 4.000 79.920 489.835 81.240 ;
        RECT 4.400 78.520 489.835 79.920 ;
        RECT 4.000 77.200 489.835 78.520 ;
        RECT 4.400 75.800 489.835 77.200 ;
        RECT 4.000 74.480 489.835 75.800 ;
        RECT 4.400 73.080 489.835 74.480 ;
        RECT 4.000 71.760 489.835 73.080 ;
        RECT 4.400 70.360 489.835 71.760 ;
        RECT 4.000 69.040 489.835 70.360 ;
        RECT 4.400 67.640 489.835 69.040 ;
        RECT 4.000 65.640 489.835 67.640 ;
        RECT 4.400 64.240 489.835 65.640 ;
        RECT 4.000 62.920 489.835 64.240 ;
        RECT 4.400 61.520 489.835 62.920 ;
        RECT 4.000 60.200 489.835 61.520 ;
        RECT 4.400 58.800 489.835 60.200 ;
        RECT 4.000 57.480 489.835 58.800 ;
        RECT 4.400 56.080 489.835 57.480 ;
        RECT 4.000 54.760 489.835 56.080 ;
        RECT 4.400 53.360 489.835 54.760 ;
        RECT 4.000 52.040 489.835 53.360 ;
        RECT 4.400 50.640 489.835 52.040 ;
        RECT 4.000 49.320 489.835 50.640 ;
        RECT 4.400 47.920 489.835 49.320 ;
        RECT 4.000 46.600 489.835 47.920 ;
        RECT 4.400 45.200 489.835 46.600 ;
        RECT 4.000 43.880 489.835 45.200 ;
        RECT 4.400 42.480 489.835 43.880 ;
        RECT 4.000 41.160 489.835 42.480 ;
        RECT 4.400 39.760 489.835 41.160 ;
        RECT 4.000 38.440 489.835 39.760 ;
        RECT 4.400 37.040 489.835 38.440 ;
        RECT 4.000 35.720 489.835 37.040 ;
        RECT 4.400 34.320 489.835 35.720 ;
        RECT 4.000 32.320 489.835 34.320 ;
        RECT 4.400 30.920 489.835 32.320 ;
        RECT 4.000 29.600 489.835 30.920 ;
        RECT 4.400 28.200 489.835 29.600 ;
        RECT 4.000 26.880 489.835 28.200 ;
        RECT 4.400 25.480 489.835 26.880 ;
        RECT 4.000 24.160 489.835 25.480 ;
        RECT 4.400 22.760 489.835 24.160 ;
        RECT 4.000 21.440 489.835 22.760 ;
        RECT 4.400 20.040 489.835 21.440 ;
        RECT 4.000 18.720 489.835 20.040 ;
        RECT 4.400 17.320 489.835 18.720 ;
        RECT 4.000 16.000 489.835 17.320 ;
        RECT 4.400 14.600 489.835 16.000 ;
        RECT 4.000 13.280 489.835 14.600 ;
        RECT 4.400 11.880 489.835 13.280 ;
        RECT 4.000 10.560 489.835 11.880 ;
        RECT 4.400 9.160 489.835 10.560 ;
        RECT 4.000 7.840 489.835 9.160 ;
        RECT 4.400 6.440 489.835 7.840 ;
        RECT 4.000 5.120 489.835 6.440 ;
        RECT 4.400 3.720 489.835 5.120 ;
        RECT 4.000 2.400 489.835 3.720 ;
        RECT 4.400 1.535 489.835 2.400 ;
      LAYER met4 ;
        RECT 7.655 288.960 388.865 291.545 ;
        RECT 7.655 15.815 20.640 288.960 ;
        RECT 23.040 15.815 97.440 288.960 ;
        RECT 99.840 15.815 174.240 288.960 ;
        RECT 176.640 15.815 251.040 288.960 ;
        RECT 253.440 15.815 327.840 288.960 ;
        RECT 330.240 15.815 388.865 288.960 ;
  END
END mkQF100Fabric
END LIBRARY

