* NGSPICE file created from mkQF100Fabric.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__fakediode_2 abstract view
.subckt sky130_ef_sc_hd__fakediode_2 DIODE VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

.subckt mkQF100Fabric CLK RST_N VGND VPWR cpu_ack_o cpu_adr_i[0] cpu_adr_i[10] cpu_adr_i[11]
+ cpu_adr_i[12] cpu_adr_i[13] cpu_adr_i[14] cpu_adr_i[15] cpu_adr_i[16] cpu_adr_i[17]
+ cpu_adr_i[18] cpu_adr_i[19] cpu_adr_i[1] cpu_adr_i[20] cpu_adr_i[21] cpu_adr_i[22]
+ cpu_adr_i[23] cpu_adr_i[24] cpu_adr_i[25] cpu_adr_i[26] cpu_adr_i[27] cpu_adr_i[28]
+ cpu_adr_i[29] cpu_adr_i[2] cpu_adr_i[30] cpu_adr_i[31] cpu_adr_i[3] cpu_adr_i[4]
+ cpu_adr_i[5] cpu_adr_i[6] cpu_adr_i[7] cpu_adr_i[8] cpu_adr_i[9] cpu_cyc_i cpu_dat_i[0]
+ cpu_dat_i[10] cpu_dat_i[11] cpu_dat_i[12] cpu_dat_i[13] cpu_dat_i[14] cpu_dat_i[15]
+ cpu_dat_i[16] cpu_dat_i[17] cpu_dat_i[18] cpu_dat_i[19] cpu_dat_i[1] cpu_dat_i[20]
+ cpu_dat_i[21] cpu_dat_i[22] cpu_dat_i[23] cpu_dat_i[24] cpu_dat_i[25] cpu_dat_i[26]
+ cpu_dat_i[27] cpu_dat_i[28] cpu_dat_i[29] cpu_dat_i[2] cpu_dat_i[30] cpu_dat_i[31]
+ cpu_dat_i[3] cpu_dat_i[4] cpu_dat_i[5] cpu_dat_i[6] cpu_dat_i[7] cpu_dat_i[8] cpu_dat_i[9]
+ cpu_dat_o[0] cpu_dat_o[10] cpu_dat_o[11] cpu_dat_o[12] cpu_dat_o[13] cpu_dat_o[14]
+ cpu_dat_o[15] cpu_dat_o[16] cpu_dat_o[17] cpu_dat_o[18] cpu_dat_o[19] cpu_dat_o[1]
+ cpu_dat_o[20] cpu_dat_o[21] cpu_dat_o[22] cpu_dat_o[23] cpu_dat_o[24] cpu_dat_o[25]
+ cpu_dat_o[26] cpu_dat_o[27] cpu_dat_o[28] cpu_dat_o[29] cpu_dat_o[2] cpu_dat_o[30]
+ cpu_dat_o[31] cpu_dat_o[3] cpu_dat_o[4] cpu_dat_o[5] cpu_dat_o[6] cpu_dat_o[7] cpu_dat_o[8]
+ cpu_dat_o[9] cpu_err_o cpu_rty_o cpu_sel_i[0] cpu_sel_i[1] cpu_sel_i[2] cpu_sel_i[3]
+ cpu_stb_i cpu_we_i spi_ack_i spi_adr_o[0] spi_adr_o[10] spi_adr_o[11] spi_adr_o[12]
+ spi_adr_o[13] spi_adr_o[14] spi_adr_o[15] spi_adr_o[16] spi_adr_o[17] spi_adr_o[18]
+ spi_adr_o[19] spi_adr_o[1] spi_adr_o[20] spi_adr_o[21] spi_adr_o[22] spi_adr_o[23]
+ spi_adr_o[24] spi_adr_o[25] spi_adr_o[26] spi_adr_o[27] spi_adr_o[28] spi_adr_o[29]
+ spi_adr_o[2] spi_adr_o[30] spi_adr_o[31] spi_adr_o[3] spi_adr_o[4] spi_adr_o[5]
+ spi_adr_o[6] spi_adr_o[7] spi_adr_o[8] spi_adr_o[9] spi_cyc_o spi_dat_i[0] spi_dat_i[10]
+ spi_dat_i[11] spi_dat_i[12] spi_dat_i[13] spi_dat_i[14] spi_dat_i[15] spi_dat_i[16]
+ spi_dat_i[17] spi_dat_i[18] spi_dat_i[19] spi_dat_i[1] spi_dat_i[20] spi_dat_i[21]
+ spi_dat_i[22] spi_dat_i[23] spi_dat_i[24] spi_dat_i[25] spi_dat_i[26] spi_dat_i[27]
+ spi_dat_i[28] spi_dat_i[29] spi_dat_i[2] spi_dat_i[30] spi_dat_i[31] spi_dat_i[3]
+ spi_dat_i[4] spi_dat_i[5] spi_dat_i[6] spi_dat_i[7] spi_dat_i[8] spi_dat_i[9] spi_dat_o[0]
+ spi_dat_o[10] spi_dat_o[11] spi_dat_o[12] spi_dat_o[13] spi_dat_o[14] spi_dat_o[15]
+ spi_dat_o[16] spi_dat_o[17] spi_dat_o[18] spi_dat_o[19] spi_dat_o[1] spi_dat_o[20]
+ spi_dat_o[21] spi_dat_o[22] spi_dat_o[23] spi_dat_o[24] spi_dat_o[25] spi_dat_o[26]
+ spi_dat_o[27] spi_dat_o[28] spi_dat_o[29] spi_dat_o[2] spi_dat_o[30] spi_dat_o[31]
+ spi_dat_o[3] spi_dat_o[4] spi_dat_o[5] spi_dat_o[6] spi_dat_o[7] spi_dat_o[8] spi_dat_o[9]
+ spi_err_i spi_rty_i spi_sel_o[0] spi_sel_o[1] spi_sel_o[2] spi_sel_o[3] spi_stb_o
+ spi_we_o
XANTENNA__2479__B1 _2119_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2106_ _2915_/Q _1914_/X _2058_/X _2523_/A VGND VGND VPWR VPWR _2624_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2037_ _2903_/Q _2018_/X _1994_/X _2508_/A VGND VGND VPWR VPWR _2610_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2651__B1 _2650_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2939_ _2946_/CLK _2939_/D VGND VGND VPWR VPWR _2939_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2403__B1 _1545_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1611__D1 _1611_/D1 VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2190__A _2190_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1757__A2 _1756_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1534__A _1534_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1693__A1 _1692_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input92_A spi_dat_i[26] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1709__A _1709_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1748__A2 _1689_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output179_A _2017_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1444__A _1444_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_6_CLK clkbuf_1_0_0_CLK/X VGND VGND VPWR VPWR _2946_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_49_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1684__A1 _1645_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2476__A3 _1528_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2275__A _2275_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2397__C1 _2231_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2724_ _2745_/CLK _2724_/D VGND VGND VPWR VPWR _2724_/Q sky130_fd_sc_hd__dfxtp_1
X_2655_ _2939_/Q _2649_/X _2650_/X VGND VGND VPWR VPWR _2939_/D sky130_fd_sc_hd__a21o_1
X_1606_ _1702_/A VGND VGND VPWR VPWR _1606_/X sky130_fd_sc_hd__buf_2
X_2586_ _2586_/A _2593_/B VGND VGND VPWR VPWR _2884_/D sky130_fd_sc_hd__nor2_1
X_1537_ _1902_/A _1530_/X _1533_/X _1536_/X input74/X VGND VGND VPWR VPWR _1537_/Y
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA__1354__A _1354_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1468_ _2949_/A _1531_/A _1467_/X VGND VGND VPWR VPWR _1616_/A sky130_fd_sc_hd__a21oi_4
X_1399_ _2772_/Q _1428_/A _1398_/Y _1431_/A VGND VGND VPWR VPWR _1509_/B sky130_fd_sc_hd__o211ai_2
XFILLER_41_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1675__A1 _1670_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1801__B _2128_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2185__A _2185_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1454__A_N _1409_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1427__A1 _1815_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1978__A2 _1961_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2632__B _2632_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1529__A _1562_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2124__S _2124_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2388__C1 _2365_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1363__B1 _1362_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1414__D _1414_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1666__A1 _1664_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2672__CLK _2920_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1418__A1 _1803_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1430__C _1454_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2542__B _2542_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2379__C1 _2231_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2034__S _2034_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2394__A2 _1785_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2440_ _1662_/X _1666_/Y _2436_/X _2431_/X VGND VGND VPWR VPWR _2792_/D sky130_fd_sc_hd__o211a_1
XFILLER_64_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2371_ _2371_/A VGND VGND VPWR VPWR _2759_/D sky130_fd_sc_hd__clkbuf_1
X_1322_ _1479_/A _1319_/Y _1321_/Y VGND VGND VPWR VPWR _2552_/A sky130_fd_sc_hd__o21ai_2
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1902__A _1902_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2082__A1 input52/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2707_ _2776_/CLK _2707_/D VGND VGND VPWR VPWR _2707_/Q sky130_fd_sc_hd__dfxtp_1
X_2638_ _2638_/A _2638_/B VGND VGND VPWR VPWR _2929_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1345__B1 _2761_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2569_ _1504_/Y _1327_/Y _2552_/B VGND VGND VPWR VPWR _2873_/D sky130_fd_sc_hd__a21o_1
XFILLER_59_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2695__CLK _2703_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1648__A1 _2181_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2346__C _2370_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2073__A1 _2839_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2339__C_N _2329_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1584__B1 _2675_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input55_A cpu_dat_i[28] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1336__B1 _1335_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2101__A2_N _2064_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1639__A1 _1576_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output211_A _1485_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2116__A2_N _1914_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1940_ _1945_/A _2591_/A VGND VGND VPWR VPWR _1940_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2553__A _2553_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1871_ _1871_/A VGND VGND VPWR VPWR _1871_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1811__B2 _2921_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1811__A1 _1807_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2272__B _2272_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2703__D _2703_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2367__A2 _1457_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1575__B1 _2780_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2423_ _1603_/X _1607_/Y _2416_/X _2405_/X VGND VGND VPWR VPWR _2784_/D sky130_fd_sc_hd__o211a_1
X_2354_ _2354_/A VGND VGND VPWR VPWR _2754_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1335__C _1335_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2524__C1 _2514_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1305_ _2366_/B _1422_/A _1354_/A _1353_/A VGND VGND VPWR VPWR _1306_/A sky130_fd_sc_hd__nand4_4
XFILLER_9_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2285_ _2285_/A VGND VGND VPWR VPWR _2725_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1632__A _1632_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2055__A1 _2836_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2182__B _2194_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1802__A1 _2850_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1566__B1 _1564_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1807__A _1807_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2515__C1 _2514_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2638__A _2638_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1542__A _1568_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2710__CLK _2873_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2860__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1717__A _1717_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1557__B1 _1473_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output161_A _1906_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1436__B _1454_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1309__B1 _2774_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2548__A _2548_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1452__A _1452_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2070_ _2075_/A _2615_/A VGND VGND VPWR VPWR _2070_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2267__B _2267_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_11_CLK_A clkbuf_1_1_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2037__B2 _2508_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2283__A _2283_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1923_ _2816_/Q _2353_/A _1922_/X VGND VGND VPWR VPWR _1923_/Y sky130_fd_sc_hd__o21ai_1
X_1854_ _2753_/Q input33/X _2127_/S VGND VGND VPWR VPWR _2350_/A sky130_fd_sc_hd__mux2_1
XANTENNA__1627__A _1699_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1785_ _2744_/Q input2/X _1785_/S VGND VGND VPWR VPWR _2330_/B sky130_fd_sc_hd__mux2_1
XFILLER_7_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2406_ _1520_/X _1550_/Y _2577_/A _2405_/X VGND VGND VPWR VPWR _2778_/D sky130_fd_sc_hd__o211a_1
XFILLER_58_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1720__B1 _1702_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2337_ _2337_/A _2355_/B _2337_/C VGND VGND VPWR VPWR _2338_/A sky130_fd_sc_hd__and3_1
XANTENNA__1362__A _1362_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2512__A2 _2506_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2177__B _2194_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2268_ _2268_/A VGND VGND VPWR VPWR _2718_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1512__D _1512_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2199_ _2199_/A _2216_/B VGND VGND VPWR VPWR _2200_/A sky130_fd_sc_hd__or2_1
XANTENNA__2733__CLK _2834_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2193__A _2193_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2028__A1 input42/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2883__CLK _2925_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2579__A2 _2401_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1787__A0 _2330_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2132__S _2132_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1847__A2_N _1792_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2368__A _2368_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1711__B1 _1709_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input18_A cpu_adr_i[24] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1490__A2 _1488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1570_ _1567_/X _1569_/X _2673_/Q VGND VGND VPWR VPWR _2158_/B sky130_fd_sc_hd__o21ai_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1950__B1 _1949_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1987__A1_N _2895_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2278__A _2278_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2756__CLK _2880_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2122_ _1859_/X _1853_/X _2582_/A VGND VGND VPWR VPWR _2122_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_6_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1910__A _1910_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2053_ _2731_/Q input47/X _2077_/S VGND VGND VPWR VPWR _2298_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1481__A2 _1788_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1769__B1 _1564_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1906_ _1906_/A VGND VGND VPWR VPWR _1906_/X sky130_fd_sc_hd__clkbuf_1
X_2886_ _2917_/CLK _2886_/D VGND VGND VPWR VPWR _2886_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2430__A1 _2427_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1837_ _2344_/B _2855_/Q _2124_/S VGND VGND VPWR VPWR _2542_/B sky130_fd_sc_hd__mux2_1
X_1768_ _1558_/X _1559_/X _2808_/Q VGND VGND VPWR VPWR _1768_/X sky130_fd_sc_hd__o21a_1
X_1699_ _1699_/A VGND VGND VPWR VPWR _1699_/X sky130_fd_sc_hd__buf_4
XANTENNA__1941__A0 _2714_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1820__A _2109_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2635__B _2639_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2127__S _2127_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2421__A1 _2412_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2370__B _2391_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2801__D _2801_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2779__CLK _2816_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1417__D _1417_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2010__A1_N _2899_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output124_A _1733_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2545__B _2545_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1448__C1 _1287_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2740_ _2834_/CLK _2740_/D VGND VGND VPWR VPWR _2740_/Q sky130_fd_sc_hd__dfxtp_1
X_2671_ _2929_/CLK _2671_/D VGND VGND VPWR VPWR _2671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1622_ _1619_/Y _1621_/Y _1606_/X VGND VGND VPWR VPWR _1622_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__2711__D _2711_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1905__A _1911_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1553_ _1551_/Y _1482_/Y _1552_/Y VGND VGND VPWR VPWR _1553_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__1923__B1 _1922_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1484_ _2076_/A VGND VGND VPWR VPWR _1945_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2479__A1 _2812_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1640__A _1712_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2105_ _2845_/Q _2251_/A _2104_/X VGND VGND VPWR VPWR _2523_/A sky130_fd_sc_hd__o21ai_2
XFILLER_35_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2036_ _2833_/Q _2033_/X _2035_/X VGND VGND VPWR VPWR _2508_/A sky130_fd_sc_hd__o21ai_1
XFILLER_63_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1552__B1_N _2704_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2100__B1 _2099_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2651__A1 _2937_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2938_ _2946_/CLK _2938_/D VGND VGND VPWR VPWR _2938_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2403__A1 _2706_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2403__B2 _1467_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1611__C1 _1565_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2190__B _2194_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2921__CLK _2925_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2869_ _2873_/CLK _2869_/D VGND VGND VPWR VPWR _2869_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1815__A _1815_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1534__B _1534_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1693__A2 _1640_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2381__A _2381_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input85_A spi_dat_i[1] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1602__C1 _1595_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1381__A1 _1379_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1669__C1 _1668_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1684__A2 _1657_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2556__A _2573_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2706__D _2706_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2944__CLK _2946_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2291__A _2296_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2723_ _2745_/CLK _2723_/D VGND VGND VPWR VPWR _2723_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2397__B1 _1309_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2149__B1 _2140_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2654_ _2654_/A VGND VGND VPWR VPWR _2938_/D sky130_fd_sc_hd__clkbuf_1
X_1605_ _2152_/B _1543_/X _2678_/Q VGND VGND VPWR VPWR _1605_/Y sky130_fd_sc_hd__o21ai_1
X_2585_ _2632_/A _2585_/B VGND VGND VPWR VPWR _2883_/D sky130_fd_sc_hd__nand2_1
X_1536_ _1710_/A VGND VGND VPWR VPWR _1536_/X sky130_fd_sc_hd__buf_2
XANTENNA__1635__A _1707_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1467_ _2705_/Q VGND VGND VPWR VPWR _1467_/X sky130_fd_sc_hd__buf_2
X_1398_ input22/X _1429_/A _1447_/C _1447_/D VGND VGND VPWR VPWR _1398_/Y sky130_fd_sc_hd__nand4b_1
XFILLER_27_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1675__A2 _1674_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1370__A _1370_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1801__C _2332_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2185__B _2185_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2019_ _2019_/A VGND VGND VPWR VPWR _2072_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__1427__A2 _1426_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2388__B1 _1329_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1363__A1 _2868_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2817__CLK _2920_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2376__A _2376_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1666__A2 _1665_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1418__A2 _1788_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1430__D _1454_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2379__B1 _1496_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output191_A _2086_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1455__A _1500_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2370_ _2370_/A _2391_/B _2370_/C VGND VGND VPWR VPWR _2371_/A sky130_fd_sc_hd__and3_1
XANTENNA__2551__B1 _2415_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1321_ _1424_/A _1380_/A _2861_/Q VGND VGND VPWR VPWR _1321_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_49_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2286__A _2296_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2706_ _2929_/CLK _2706_/D VGND VGND VPWR VPWR _2706_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput210 _2949_/X VGND VGND VPWR VPWR spi_stb_o sky130_fd_sc_hd__buf_2
X_2637_ _2637_/A _2639_/B VGND VGND VPWR VPWR _2928_/D sky130_fd_sc_hd__nor2_1
XANTENNA__1365__A _2869_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1345__A1 _1307_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2568_ _2401_/C _2358_/X _2384_/A _1503_/Y _2558_/X VGND VGND VPWR VPWR _2872_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_59_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2499_ _2826_/Q _2493_/X _1990_/X _2488_/X VGND VGND VPWR VPWR _2826_/D sky130_fd_sc_hd__o211a_1
X_1519_ _1682_/A VGND VGND VPWR VPWR _1519_/X sky130_fd_sc_hd__buf_2
XFILLER_56_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1648__A2 _2181_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2073__A2 _2033_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1584__A1 _1567_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1336__A1 _2880_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input48_A cpu_dat_i[21] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1639__A2 _1588_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output204_A _1980_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1870_ _1878_/A _2931_/Q VGND VGND VPWR VPWR _1871_/A sky130_fd_sc_hd__and2_1
XANTENNA__1811__A2 _2534_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1575__A1 _1517_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2422_ _2408_/X _2410_/X _2421_/Y VGND VGND VPWR VPWR _2783_/D sky130_fd_sc_hd__o21ai_1
X_2353_ _2353_/A _2353_/B _2352_/X VGND VGND VPWR VPWR _2354_/A sky130_fd_sc_hd__or3b_1
XANTENNA__2524__B1 _2109_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1913__A _1913_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1304_ _1304_/A VGND VGND VPWR VPWR _1422_/A sky130_fd_sc_hd__buf_2
X_2284_ _2284_/A _2284_/B _2289_/C VGND VGND VPWR VPWR _2285_/A sky130_fd_sc_hd__and3_1
XFILLER_49_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2055__A2 _2025_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1802__A2 _2474_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2460__C1 _2451_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1999_ _2011_/A _2602_/A VGND VGND VPWR VPWR _1999_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__1566__A1 _1561_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2515__B1 _2067_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2638__B _2638_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2654__A _2654_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input102_A spi_dat_i[6] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2306__C_N _2305_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2804__D _2804_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1557__A1 _1520_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1309__A1 _1307_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1436__C _1454_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output154_A _1890_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2548__B _2548_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2714__D _2714_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1922_ _2364_/A _2358_/A _2249_/A VGND VGND VPWR VPWR _1922_/X sky130_fd_sc_hd__or3_1
X_1853_ _1853_/A VGND VGND VPWR VPWR _1853_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__2685__CLK _2839_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1908__A _1908_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1784_ _2113_/S VGND VGND VPWR VPWR _1785_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_6_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2405_ _2451_/A VGND VGND VPWR VPWR _2405_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1525__A1_N _1504_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1720__A1 _2203_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2336_ _2526_/A VGND VGND VPWR VPWR _2355_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1362__B _1362_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2267_ _2272_/A _2267_/B _2257_/X VGND VGND VPWR VPWR _2268_/A sky130_fd_sc_hd__or3b_1
XFILLER_38_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2198_ _2198_/A VGND VGND VPWR VPWR _2216_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_25_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2474__A _2474_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2193__B _2193_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1787__A1 _2849_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1818__A _2027_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2649__A _2649_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1711__A1 _1651_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2368__B _2368_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2384__A _2384_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1447__B _1454_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1950__A1 _2820_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1463__A _2706_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2121_ _2882_/Q _1530_/X _1840_/X _2120_/Y VGND VGND VPWR VPWR _2582_/A sky130_fd_sc_hd__a2bb2o_2
XANTENNA__2709__D _2709_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2052_ _2075_/A _2612_/A VGND VGND VPWR VPWR _2052_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2294__A _2294_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1481__A3 _1803_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1769__A1 _1723_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1905_ _1911_/A _2667_/Q VGND VGND VPWR VPWR _1906_/A sky130_fd_sc_hd__and2_1
XANTENNA__1638__A _1710_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2885_ _2925_/CLK _2885_/D VGND VGND VPWR VPWR _2885_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2430__A2 _2428_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1836_ _2750_/Q input30/X _1860_/S VGND VGND VPWR VPWR _2344_/B sky130_fd_sc_hd__mux2_1
X_1767_ _1763_/X _1766_/Y _1632_/A _1633_/A VGND VGND VPWR VPWR _1767_/X sky130_fd_sc_hd__o211a_1
X_1698_ _1698_/A VGND VGND VPWR VPWR _1698_/X sky130_fd_sc_hd__buf_4
XANTENNA__1941__A1 input60/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2700__CLK _2703_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2319_ _2319_/A VGND VGND VPWR VPWR _2739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1820__B _1865_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2850__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2406__C1 _2405_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1548__A _1548_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2421__A2 _2168_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2370__C _2370_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_leaf_10_CLK_A clkbuf_1_1_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2069__A2_N _2064_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input30_A cpu_adr_i[6] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output117_A _1688_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1448__B1 _1447_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2670_ _2670_/CLK _2670_/D VGND VGND VPWR VPWR _2670_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2053__S _2077_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1621_ _1620_/X _1543_/X _2680_/Q VGND VGND VPWR VPWR _1621_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2723__CLK _2745_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1552_ _1744_/A _1568_/A _2704_/Q VGND VGND VPWR VPWR _1552_/Y sky130_fd_sc_hd__o21bai_1
XANTENNA__1923__A1 _2816_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1905__B _2667_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1483_ _1778_/A _1807_/A _1482_/Y VGND VGND VPWR VPWR _2076_/A sky130_fd_sc_hd__a21o_4
XANTENNA__2289__A _2289_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2479__A2 _2475_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2873__CLK _2873_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1687__B1 _1630_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2104_ _2114_/A _2114_/B _2320_/B VGND VGND VPWR VPWR _2104_/X sky130_fd_sc_hd__or3_1
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2035_ _2035_/A _2072_/B _2291_/B VGND VGND VPWR VPWR _2035_/X sky130_fd_sc_hd__or3_1
XANTENNA__1439__B1 _2874_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2100__A1 _2844_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2651__A2 _2649_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2937_ _2946_/CLK _2937_/D VGND VGND VPWR VPWR _2937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2403__A2 _2529_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2902__D _2902_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1611__B1 _1564_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2868_ _2873_/CLK _2868_/D VGND VGND VPWR VPWR _2868_/Q sky130_fd_sc_hd__dfxtp_1
X_2799_ _2809_/CLK _2799_/D VGND VGND VPWR VPWR _2799_/Q sky130_fd_sc_hd__dfxtp_1
X_1819_ _2747_/Q input27/X _2108_/S VGND VGND VPWR VPWR _2337_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2199__A _2199_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1678__B1 _2688_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2627__C1 _2626_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2947__212 VGND VGND VPWR VPWR _2947__212/HI cpu_err_o sky130_fd_sc_hd__conb_1
XFILLER_60_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2662__A _2665_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1850__A0 _2348_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2812__D _2812_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1602__B1 _1593_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2746__CLK _2925_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input78_A spi_dat_i[13] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2896__CLK _2917_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1381__A2 _1488_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1924__A1_N _2886_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1669__B1 _1667_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2556__B _2556_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2048__S _2093_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1939__A1_N _2888_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2291__B _2291_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2722_ _2745_/CLK _2722_/D VGND VGND VPWR VPWR _2722_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2722__D _2722_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2397__A1 _1301_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2149__A1 _2669_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2653_ _2665_/A _2938_/Q _2653_/C VGND VGND VPWR VPWR _2654_/A sky130_fd_sc_hd__and3_1
XANTENNA__1916__A _2058_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1604_ _1576_/X _1588_/X _1533_/X _1536_/X _1604_/D1 VGND VGND VPWR VPWR _1604_/Y
+ sky130_fd_sc_hd__o2111ai_2
X_2584_ _2618_/A VGND VGND VPWR VPWR _2632_/A sky130_fd_sc_hd__clkbuf_2
X_1535_ _1699_/A VGND VGND VPWR VPWR _1710_/A sky130_fd_sc_hd__buf_2
X_1466_ input73/X _1465_/X _2705_/Q VGND VGND VPWR VPWR _1531_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__1651__A _1723_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1397_ _2865_/Q _1287_/X _1396_/Y VGND VGND VPWR VPWR _2560_/B sky130_fd_sc_hd__o21ai_2
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1370__B _1409_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2018_ _2233_/A VGND VGND VPWR VPWR _2018_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2085__B1 _2058_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2769__CLK _2776_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2388__A1 _2366_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1596__C1 _1595_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1826__A _2243_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1363__A2 _1324_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2657__A _2657_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1561__A _1717_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2807__D _2807_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1418__A3 _1803_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1823__B1 _2631_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2392__A _2392_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2379__A1 _1367_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output184_A _2052_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1455__B _1455_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1320_ _1400_/A _1401_/A _1422_/A VGND VGND VPWR VPWR _1380_/A sky130_fd_sc_hd__o21a_2
XANTENNA__2551__A1 _1528_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2717__D _2717_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2286__B _2286_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2911__CLK _2915_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1504__B1_N _2873_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2705_ _2929_/CLK _2705_/D VGND VGND VPWR VPWR _2705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput200 _1952_/Y VGND VGND VPWR VPWR spi_dat_o[4] sky130_fd_sc_hd__buf_2
X_2636_ _2638_/A _2636_/B VGND VGND VPWR VPWR _2927_/D sky130_fd_sc_hd__nand2_1
Xoutput211 _1485_/Y VGND VGND VPWR VPWR spi_we_o sky130_fd_sc_hd__buf_2
XANTENNA__1345__A2 _1308_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2567_ _1493_/Y _1339_/Y _2552_/B VGND VGND VPWR VPWR _2871_/D sky130_fd_sc_hd__a21o_1
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2498_ _2498_/A _2508_/B VGND VGND VPWR VPWR _2825_/D sky130_fd_sc_hd__nand2_1
X_1518_ _1616_/A VGND VGND VPWR VPWR _1682_/A sky130_fd_sc_hd__buf_2
XFILLER_59_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2477__A _2531_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1449_ _1449_/A _1449_/B VGND VGND VPWR VPWR _1508_/C sky130_fd_sc_hd__nand2_1
XFILLER_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1502__C1 _1311_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1805__B1 _1802_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1584__A2 _1569_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1556__A _1740_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1336__A2 _1324_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1741__C1 _1740_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2934__CLK _2946_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1291__A _1291_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1575__A2 _1519_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1490__B1_N _2880_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2421_ _2412_/X _2168_/A _1597_/X VGND VGND VPWR VPWR _2421_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__2524__A1 _2846_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2352_ _2352_/A VGND VGND VPWR VPWR _2352_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2283_ _2283_/A VGND VGND VPWR VPWR _2724_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2297__A _2297_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1303_ _1400_/A VGND VGND VPWR VPWR _2366_/B sky130_fd_sc_hd__clkinv_2
XFILLER_49_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2460__B1 _2456_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1998_ _2897_/Q _1953_/X _1994_/X _2500_/A VGND VGND VPWR VPWR _2602_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__2807__CLK _2809_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2910__D _2910_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1566__A2 _2064_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1376__A _1376_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2258__C_N _2257_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2619_ _2619_/A _2626_/B VGND VGND VPWR VPWR _2911_/D sky130_fd_sc_hd__nand2_1
XANTENNA__2515__A1 _2838_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2000__A _2064_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1286__A _1343_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2820__D _2820_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1557__A2 _1550_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input60_A cpu_dat_i[3] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1436__D _1454_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1309__A2 _1308_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output147_A _1877_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1493__A1 _1445_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2442__B1 _2441_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1921_ _2711_/Q input35/X _2132_/S VGND VGND VPWR VPWR _2249_/A sky130_fd_sc_hd__mux2_1
X_1852_ _1830_/X _1824_/X _2636_/B VGND VGND VPWR VPWR _1852_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__2580__A _2580_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2730__D _2730_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1783_ _2047_/A VGND VGND VPWR VPWR _2113_/S sky130_fd_sc_hd__buf_4
X_2404_ _2395_/A _2366_/A _2231_/A _1469_/Y _2403_/Y VGND VGND VPWR VPWR _2777_/D
+ sky130_fd_sc_hd__o2111a_1
X_2335_ _2335_/A VGND VGND VPWR VPWR _2746_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1720__A2 _2203_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2266_ _2266_/A VGND VGND VPWR VPWR _2717_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1362__C _1362_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2197_ _2197_/A _2197_/B VGND VGND VPWR VPWR _2199_/A sky130_fd_sc_hd__nand2_1
XFILLER_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2905__D _2905_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2490__A _2490_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1711__A2 _1663_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2665__A _2665_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2384__B _2391_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2815__D _2815_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2424__B1 _1610_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2573__C_N _2415_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1447__C _1447_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1744__A _1744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1950__A2 _2353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2120_ _2812_/Q _1841_/X _2119_/X VGND VGND VPWR VPWR _2120_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2051_ _2905_/Q _2018_/X _1994_/X _2511_/A VGND VGND VPWR VPWR _2612_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_19_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1466__A1 input73/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2294__B _2308_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2725__D _2725_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1904_ _1904_/A VGND VGND VPWR VPWR _1904_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1769__A2 _2533_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1919__A _2019_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2884_ _2920_/CLK _2884_/D VGND VGND VPWR VPWR _2884_/Q sky130_fd_sc_hd__dfxtp_1
X_1835_ _1830_/X _1824_/X _2633_/A VGND VGND VPWR VPWR _1835_/Y sky130_fd_sc_hd__a21oi_2
X_1766_ _2219_/A _2219_/B _1549_/X VGND VGND VPWR VPWR _1766_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_7_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1697_ _1696_/X _1682_/X _2797_/Q VGND VGND VPWR VPWR _1697_/X sky130_fd_sc_hd__o21a_1
XFILLER_44_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ _2318_/A _2332_/B _2337_/C VGND VGND VPWR VPWR _2319_/A sky130_fd_sc_hd__and3_1
XFILLER_26_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2249_ _2249_/A _2260_/B _2265_/C VGND VGND VPWR VPWR _2250_/A sky130_fd_sc_hd__and3_1
XFILLER_25_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1820__C _2337_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2406__B1 _2577_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1564__A _1698_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1393__B1 _1392_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1283__B _1289_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput100 spi_dat_i[4] VGND VGND VPWR VPWR _1589_/D1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__2675__CLK _2816_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input23_A cpu_adr_i[29] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2395__A _2395_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1448__A1 _2760_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1739__A _1739_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1620_ _1692_/A VGND VGND VPWR VPWR _1620_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1474__A _2671_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1551_ _2949_/A _1698_/A VGND VGND VPWR VPWR _1551_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__1923__A2 _2353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1384__B1 _2769_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1482_ _1807_/A _2527_/B _1481_/X VGND VGND VPWR VPWR _1482_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_4_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2289__B _2308_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_9_CLK clkbuf_1_1_0_CLK/X VGND VGND VPWR VPWR _2915_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1687__A1 _2193_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2103_ _2740_/Q input56/X _2113_/S VGND VGND VPWR VPWR _2320_/B sky130_fd_sc_hd__mux2_1
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2034_ _2728_/Q input43/X _2034_/S VGND VGND VPWR VPWR _2291_/B sky130_fd_sc_hd__mux2_1
XANTENNA__1439__A1 _1815_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2100__A2 _1814_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2936_ _2946_/CLK _2936_/D VGND VGND VPWR VPWR _2936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1611__A1 _1561_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2867_ _2929_/CLK _2867_/D VGND VGND VPWR VPWR _2867_/Q sky130_fd_sc_hd__dfxtp_1
X_1818_ _2027_/A VGND VGND VPWR VPWR _2108_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_11_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2798_ _2840_/CLK _2798_/D VGND VGND VPWR VPWR _2798_/Q sky130_fd_sc_hd__dfxtp_1
X_1749_ _1723_/X _2533_/A _1709_/X _1710_/X input92/X VGND VGND VPWR VPWR _1749_/Y
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA__2572__C1 _2558_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1375__B1 _1374_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2698__CLK _2703_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2199__B _2216_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1678__A1 _1620_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2627__B1 _1481_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2662__B _2944_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1850__A1 _2857_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1559__A _1682_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1602__A1 _1597_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1294__A _1414_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1669__A1 _1662_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1469__A _2811_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2721_ _2745_/CLK _2721_/D VGND VGND VPWR VPWR _2721_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2397__A2 _1457_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2149__A2 _2136_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2652_ _2652_/A VGND VGND VPWR VPWR _2665_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2583_ _1567_/X _1569_/X _2312_/A VGND VGND VPWR VPWR _2618_/A sky130_fd_sc_hd__o21a_4
XANTENNA__1357__B1 _2759_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2840__CLK _2840_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1603_ _1517_/X _1519_/X _2784_/Q VGND VGND VPWR VPWR _1603_/X sky130_fd_sc_hd__o21a_1
X_1534_ _1534_/A _1534_/B input73/X VGND VGND VPWR VPWR _1699_/A sky130_fd_sc_hd__nor3b_4
XANTENNA__2291__C_N _2281_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1932__A _1945_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1465_ _1534_/A _1534_/B VGND VGND VPWR VPWR _1465_/X sky130_fd_sc_hd__or2_4
X_1396_ _2372_/B _2372_/C _1437_/A VGND VGND VPWR VPWR _1396_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__1416__A1_N _1408_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2017_ _2044_/A _2605_/A VGND VGND VPWR VPWR _2017_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2085__B2 _2518_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1379__A _1424_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2913__D _2913_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2919_ _2925_/CLK _2919_/D VGND VGND VPWR VPWR _2919_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2388__A2 _1330_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1596__B1 _1593_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2003__A _2014_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1842__A _2046_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1520__B1 _2778_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2713__CLK _2776_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1823__A1 _1779_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2823__D _2823_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1289__A _1289_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input90_A spi_dat_i[24] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2379__A2 _1457_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2863__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1587__B1 _2782_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output177_A _2006_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1455__C _1455_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2536__C1 _2531_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2551__A2 _1528_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2059__S _2093_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2733__D _2733_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1927__A _2058_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1578__B1 _2674_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2704_ _2929_/CLK _2704_/D VGND VGND VPWR VPWR _2704_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput201 _1959_/Y VGND VGND VPWR VPWR spi_dat_o[5] sky130_fd_sc_hd__buf_2
X_2635_ _2635_/A _2639_/B VGND VGND VPWR VPWR _2926_/D sky130_fd_sc_hd__nor2_1
X_2566_ _2357_/X _2358_/X _2380_/A _1381_/Y _2558_/X VGND VGND VPWR VPWR _2870_/D
+ sky130_fd_sc_hd__o311a_1
XANTENNA__1750__B1 _2698_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2497_ _2510_/A VGND VGND VPWR VPWR _2508_/B sky130_fd_sc_hd__clkbuf_2
X_1517_ _1707_/A VGND VGND VPWR VPWR _1517_/X sky130_fd_sc_hd__buf_2
X_1448_ _2760_/Q _1428_/A _1447_/Y _1287_/X VGND VGND VPWR VPWR _1449_/B sky130_fd_sc_hd__o211ai_1
XFILLER_56_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2908__D _2908_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2736__CLK _2834_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1502__B1 _1406_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1379_ _1424_/A VGND VGND VPWR VPWR _1379_/X sky130_fd_sc_hd__buf_2
XFILLER_64_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2493__A _2493_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2886__CLK _2917_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1805__B2 _1804_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1572__A _1630_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1741__B1 _1739_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2818__D _2818_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2509__C1 _2501_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2420_ _1587_/X _1591_/Y _2416_/X _2405_/X VGND VGND VPWR VPWR _2782_/D sky130_fd_sc_hd__o211a_1
X_2351_ _2351_/A VGND VGND VPWR VPWR _2753_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2759__CLK _2768_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2524__A2 _2519_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1732__B1 _1702_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2282_ _2296_/A _2282_/B _2281_/X VGND VGND VPWR VPWR _2283_/A sky130_fd_sc_hd__or3b_1
X_1302_ _2777_/Q VGND VGND VPWR VPWR _1400_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2085__A1_N _2911_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2728__D _2728_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2460__A1 _1734_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2023__A1_N _2901_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1997_ _2827_/Q _1969_/X _1996_/X VGND VGND VPWR VPWR _2500_/A sky130_fd_sc_hd__o21ai_1
XFILLER_21_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1657__A _1735_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2618_ _2618_/A VGND VGND VPWR VPWR _2626_/B sky130_fd_sc_hd__buf_4
XFILLER_47_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2549_ _2549_/A VGND VGND VPWR VPWR _2859_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2515__A2 _2506_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2488__A _2531_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1487__C1 _1500_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1567__A _1744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2901__CLK _2901_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input53_A cpu_dat_i[26] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2398__A _2398_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1714__B1 _1679_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1503__B1_N _2872_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1493__A2 _1488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1920_ _2113_/S VGND VGND VPWR VPWR _2132_/S sky130_fd_sc_hd__buf_4
XANTENNA__2442__A1 _2427_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1851_ _1807_/X _2545_/B _1789_/X _2927_/Q VGND VGND VPWR VPWR _2636_/B sky130_fd_sc_hd__o22ai_2
XFILLER_30_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1477__A _1477_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1782_ _1807_/A VGND VGND VPWR VPWR _2649_/A sky130_fd_sc_hd__buf_4
XFILLER_11_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2403_ _2706_/Q _2529_/A _1545_/Y _1467_/X VGND VGND VPWR VPWR _2403_/Y sky130_fd_sc_hd__o22ai_1
X_2334_ _2344_/A _2334_/B _2329_/X VGND VGND VPWR VPWR _2335_/A sky130_fd_sc_hd__or3b_1
XANTENNA__1940__A _1945_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2265_ _2265_/A _2284_/B _2265_/C VGND VGND VPWR VPWR _2266_/A sky130_fd_sc_hd__and3_1
X_2196_ _1691_/Y _1693_/Y _2179_/X VGND VGND VPWR VPWR _2690_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__2130__B1 _1840_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2490__B _2495_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2924__CLK _2930_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2921__D _2921_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1944__B1 _1927_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2011__A _2011_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2665__B _2946_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2121__B1 _1840_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2384__C _2399_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2424__A1 _2412_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2831__D _2831_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1297__A _1372_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2188__B1 _2179_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1447__D _1447_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2050_ _2835_/Q _2033_/X _2049_/X VGND VGND VPWR VPWR _2511_/A sky130_fd_sc_hd__o21ai_1
XFILLER_47_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1466__A2 _1465_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2294__C _2313_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2591__A _2591_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1903_ _1911_/A _2946_/Q VGND VGND VPWR VPWR _1904_/A sky130_fd_sc_hd__and2_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1623__C1 _1595_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2883_ _2925_/CLK _2883_/D VGND VGND VPWR VPWR _2883_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2741__D _2741_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1834_ _2924_/Q _1792_/X _1804_/X _1833_/Y VGND VGND VPWR VPWR _2633_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1765_ _1744_/X _1543_/A _2701_/Q VGND VGND VPWR VPWR _2219_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__1935__A _2114_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1696_ _1696_/A VGND VGND VPWR VPWR _1696_/X sky130_fd_sc_hd__clkbuf_2
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ _2362_/A VGND VGND VPWR VPWR _2337_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_57_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2248_ _2248_/A VGND VGND VPWR VPWR _2710_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2916__D _2916_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2103__A0 _2740_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2179_ _2224_/B VGND VGND VPWR VPWR _2179_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2406__A1 _1520_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2006__A _2011_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1845__A _2128_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1393__A1 _1389_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput101 spi_dat_i[5] VGND VGND VPWR VPWR _1598_/D1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__1283__C _1291_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input16_A cpu_adr_i[22] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2395__B _2395_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2826__D _2826_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1448__A2 _1428_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1550_ _1537_/Y _1544_/Y _1549_/X VGND VGND VPWR VPWR _1550_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1384__A1 _1451_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1481_ _1803_/A _1788_/B _1803_/D _2918_/Q VGND VGND VPWR VPWR _1481_/X sky130_fd_sc_hd__a31o_1
XANTENNA__2289__C _2289_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1381__B1_N _2870_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2586__A _2586_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2102_ _2102_/A _2623_/A VGND VGND VPWR VPWR _2102_/Y sky130_fd_sc_hd__nor2_2
XFILLER_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1687__A2 _2193_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2736__D _2736_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2033_ _2033_/A VGND VGND VPWR VPWR _2033_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1439__A2 _1426_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2935_ _2946_/CLK _2935_/D VGND VGND VPWR VPWR _2935_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1611__A2 _1582_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2866_ _2880_/CLK _2866_/D VGND VGND VPWR VPWR _2866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1817_ _2065_/A VGND VGND VPWR VPWR _1865_/B sky130_fd_sc_hd__clkbuf_1
X_2797_ _2839_/CLK _2797_/D VGND VGND VPWR VPWR _2797_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2572__B1 _1408_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1375__A1 _2867_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1748_ _1707_/X _1689_/X _2804_/Q VGND VGND VPWR VPWR _1748_/X sky130_fd_sc_hd__o21a_1
X_1679_ _1702_/A VGND VGND VPWR VPWR _1679_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input8_A cpu_adr_i[15] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1678__A2 _1640_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2627__A1 _1781_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2662__C _2665_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1602__A2 _1601_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1294__B _1354_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1669__A2 _1666_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2792__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output122_A _1721_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2720_ _2745_/CLK _2720_/D VGND VGND VPWR VPWR _2720_/Q sky130_fd_sc_hd__dfxtp_1
X_2651_ _2937_/Q _2649_/X _2650_/X VGND VGND VPWR VPWR _2937_/D sky130_fd_sc_hd__a21o_1
XFILLER_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1485__A _1945_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1602_ _1597_/X _1601_/Y _1593_/X _1595_/X VGND VGND VPWR VPWR _1602_/X sky130_fd_sc_hd__o211a_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2582_ _2582_/A _2593_/B VGND VGND VPWR VPWR _2882_/D sky130_fd_sc_hd__nor2_1
XANTENNA__1357__A1 _1307_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1447__A_N input9/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1533_ _1709_/A VGND VGND VPWR VPWR _1533_/X sky130_fd_sc_hd__buf_2
X_1464_ _1342_/A _1342_/B _1528_/B _1463_/Y VGND VGND VPWR VPWR _1464_/X sky130_fd_sc_hd__o31a_2
XANTENNA__1932__B _2590_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1395_ _1451_/A _1452_/A _2760_/Q VGND VGND VPWR VPWR _2372_/C sky130_fd_sc_hd__o21ai_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2016_ _2900_/Q _2000_/X _1975_/X _2015_/Y VGND VGND VPWR VPWR _2605_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2918_ _2929_/CLK _2918_/D VGND VGND VPWR VPWR _2918_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2388__A3 _2366_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1596__A1 _1587_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2849_ _2925_/CLK _2849_/D VGND VGND VPWR VPWR _2849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2003__B _2054_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1520__A1 _1517_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_opt_2_1_CLK clkbuf_opt_2_1_CLK/A VGND VGND VPWR VPWR clkbuf_opt_2_1_CLK/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_57_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1823__A2 _1781_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1284__B1 _2881_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input83_A spi_dat_i[18] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1587__A1 _1517_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2536__B1 _1820_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2688__CLK _2839_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1578__A1 _2152_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2703_ _2703_/CLK _2703_/D VGND VGND VPWR VPWR _2703_/Q sky130_fd_sc_hd__dfxtp_1
X_2634_ _2638_/A _2634_/B VGND VGND VPWR VPWR _2925_/D sky130_fd_sc_hd__nand2_1
XANTENNA__2104__A _2114_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput202 _1968_/Y VGND VGND VPWR VPWR spi_dat_o[6] sky130_fd_sc_hd__buf_2
X_2565_ _1495_/Y _1497_/Y _2552_/B VGND VGND VPWR VPWR _2869_/D sky130_fd_sc_hd__a21o_1
X_1516_ _1696_/A VGND VGND VPWR VPWR _1707_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__1750__A1 _1692_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2496_ _2824_/Q _2493_/X _1977_/X _2488_/X VGND VGND VPWR VPWR _2824_/D sky130_fd_sc_hd__o211a_1
X_1447_ input9/X _1454_/B _1447_/C _1447_/D VGND VGND VPWR VPWR _1447_/Y sky130_fd_sc_hd__nand4b_1
X_1378_ _1436_/A _1306_/A _1377_/Y VGND VGND VPWR VPWR _2380_/A sky130_fd_sc_hd__o21ai_4
XFILLER_56_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1967__A2_N _1933_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1502__A1 _2879_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2924__D _2924_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2463__C1 _2451_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2014__A _2014_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2949__A _2949_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1853__A _1853_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1741__A1 _1734_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2830__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2834__D _2834_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2509__B1 _2041_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1732__A1 _2207_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2350_ _2350_/A _2355_/B _2370_/C VGND VGND VPWR VPWR _2351_/A sky130_fd_sc_hd__and3_1
X_1301_ _1301_/A VGND VGND VPWR VPWR _1301_/Y sky130_fd_sc_hd__inv_2
X_2281_ _2352_/A VGND VGND VPWR VPWR _2281_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2594__A _2618_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1496__B1 _2764_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2744__D _2744_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2460__A2 _1738_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1996_ _2035_/A _2008_/B _2277_/B VGND VGND VPWR VPWR _1996_/X sky130_fd_sc_hd__or3_1
XFILLER_20_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2005__A2_N _2000_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2617_ _2617_/A _2617_/B VGND VGND VPWR VPWR _2910_/D sky130_fd_sc_hd__nor2_1
XANTENNA__2703__CLK _2703_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2548_ _2548_/A _2548_/B _2537_/X VGND VGND VPWR VPWR _2549_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2919__D _2919_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2479_ _2812_/Q _2475_/X _2119_/X _2525_/B VGND VGND VPWR VPWR _2812_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2853__CLK _2925_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1487__B1 _1377_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2130__A1_N _2884_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2398__B _2398_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1714__A1 _1711_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2829__D _2829_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input46_A cpu_dat_i[1] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1478__A0 _2743_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output202_A _1968_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2442__A2 _2428_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1850_ _2348_/B _2857_/Q _2124_/S VGND VGND VPWR VPWR _2545_/B sky130_fd_sc_hd__mux2_1
XANTENNA__1650__B1 _2790_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1781_ _1853_/A VGND VGND VPWR VPWR _1781_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__2726__CLK _2834_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1402__B1 _1422_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2589__A _2618_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2402_ _2402_/A VGND VGND VPWR VPWR _2776_/D sky130_fd_sc_hd__clkbuf_1
X_2333_ _2333_/A VGND VGND VPWR VPWR _2745_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2363__D1 _2382_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2739__D _2739_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2876__CLK _2880_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1940__B _2591_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2264_ _2312_/A VGND VGND VPWR VPWR _2284_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_2195_ _2195_/A VGND VGND VPWR VPWR _2689_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2130__B2 _2129_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1668__A _1740_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1641__B1 _2682_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1387__B _1387_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1979_ _2894_/Q _1933_/X _1975_/X _1978_/Y VGND VGND VPWR VPWR _2599_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__1944__B2 _2490_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2011__B _2604_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2665__C _2665_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2121__B2 _2120_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input100_A spi_dat_i[4] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2409__C1 _2366_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2424__A2 _2172_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2749__CLK _2768_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2188__A1 _1664_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2899__CLK _2901_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output152_A _1806_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2037__A1_N _2903_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2591__B _2593_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1902_ _1902_/A VGND VGND VPWR VPWR _1911_/A sky130_fd_sc_hd__clkbuf_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1488__A _1488_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1623__B1 _1593_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2882_ _2920_/CLK _2882_/D VGND VGND VPWR VPWR _2882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1833_ _2854_/Q _1814_/X _1832_/X VGND VGND VPWR VPWR _1833_/Y sky130_fd_sc_hd__o21ai_1
X_1764_ _1717_/X _1729_/X _1709_/A _1710_/A input95/X VGND VGND VPWR VPWR _2219_/A
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA__2112__A _2117_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1695_ _1690_/X _1694_/Y _1667_/X _1668_/X VGND VGND VPWR VPWR _1695_/X sky130_fd_sc_hd__o211a_1
XFILLER_44_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2316_ _2316_/A VGND VGND VPWR VPWR _2738_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2247_ _2540_/A _2247_/B _2227_/A VGND VGND VPWR VPWR _2248_/A sky130_fd_sc_hd__or3b_1
XFILLER_54_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2103__A1 input56/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2178_ _2178_/A VGND VGND VPWR VPWR _2681_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1311__C1 _1431_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1862__B1 _1789_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2406__A2 _1550_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2932__D _2932_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1614__B1 _1572_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2006__B _2603_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1845__B _1865_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1393__A2 _1287_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput102 spi_dat_i[6] VGND VGND VPWR VPWR _1604_/D1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2395__C _2395_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1800__S _1970_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1605__B1 _2678_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2842__D _2842_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2030__B1 _2029_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1384__A2 _1452_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1480_ _2327_/A _2848_/Q _2243_/A VGND VGND VPWR VPWR _2527_/B sky130_fd_sc_hd__mux2_1
XFILLER_4_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2586__B _2593_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2101_ _2914_/Q _2064_/X _1804_/X _2100_/Y VGND VGND VPWR VPWR _2623_/A sky130_fd_sc_hd__a2bb2o_4
XFILLER_55_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2032_ _2044_/A _2609_/A VGND VGND VPWR VPWR _2032_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2914__CLK _2920_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1844__A0 _2751_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2752__D _2752_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2934_ _2946_/CLK _2934_/D VGND VGND VPWR VPWR _2934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2107__A _2117_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2865_ _2873_/CLK _2865_/D VGND VGND VPWR VPWR _2865_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1946__A _2076_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1816_ _2114_/A VGND VGND VPWR VPWR _2109_/A sky130_fd_sc_hd__buf_2
X_2796_ _2839_/CLK _2796_/D VGND VGND VPWR VPWR _2796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2572__A1 _2401_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1375__A2 _1343_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1747_ _1742_/X _1746_/Y _1739_/X _1740_/X VGND VGND VPWR VPWR _1747_/X sky130_fd_sc_hd__o211a_1
X_1678_ _1620_/X _1640_/X _2688_/Q VGND VGND VPWR VPWR _1678_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_58_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2927__D _2927_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2627__A2 _2527_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1835__B1 _2633_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2017__A _2044_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1294__C _1294_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2937__CLK _2946_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2837__D _2837_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2079__B1 _2078_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output115_A _1675_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2650_ _2650_/A VGND VGND VPWR VPWR _2650_/X sky130_fd_sc_hd__clkbuf_2
X_1601_ _2167_/A _2167_/B _1572_/X VGND VGND VPWR VPWR _1601_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2581_ _2650_/A VGND VGND VPWR VPWR _2593_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__1357__A2 _1308_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1532_ _1698_/A VGND VGND VPWR VPWR _1709_/A sky130_fd_sc_hd__buf_2
XANTENNA__2597__A _2597_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1762__C1 _1740_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1463_ _2706_/Q VGND VGND VPWR VPWR _1463_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2747__D _2747_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1394_ input9/X _1409_/B VGND VGND VPWR VPWR _2372_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2015_ _2830_/Q _1961_/X _2014_/X VGND VGND VPWR VPWR _2015_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_63_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2917_ _2917_/CLK _2917_/D VGND VGND VPWR VPWR _2917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1596__A2 _1591_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2848_ _2929_/CLK _2848_/D VGND VGND VPWR VPWR _2848_/Q sky130_fd_sc_hd__dfxtp_1
X_2779_ _2816_/CLK _2779_/D VGND VGND VPWR VPWR _2779_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2003__C _2279_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2300__A _2324_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1520__A2 _1519_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1284__A1 _1304_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1587__A2 _1519_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input76_A spi_dat_i[11] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2536__A1 _2852_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_opt_2_1_CLK_A clkbuf_opt_2_1_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_10_CLK clkbuf_1_1_0_CLK/X VGND VGND VPWR VPWR _2901_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2472__B1 _1556_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1578__A2 _1543_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2702_ _2816_/CLK _2702_/D VGND VGND VPWR VPWR _2702_/Q sky130_fd_sc_hd__dfxtp_1
X_2633_ _2633_/A _2639_/B VGND VGND VPWR VPWR _2924_/D sky130_fd_sc_hd__nor2_1
XANTENNA__2104__B _2114_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput203 _1974_/Y VGND VGND VPWR VPWR spi_dat_o[7] sky130_fd_sc_hd__buf_2
X_2564_ _2868_/Q _2540_/X _2554_/X _1362_/Y VGND VGND VPWR VPWR _2868_/D sky130_fd_sc_hd__o211a_1
X_1515_ _1515_/A VGND VGND VPWR VPWR _1696_/A sky130_fd_sc_hd__clkbuf_4
X_2495_ _2495_/A _2495_/B VGND VGND VPWR VPWR _2823_/D sky130_fd_sc_hd__nand2_1
XANTENNA__1750__A2 _1712_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1446_ _1445_/X _1426_/X _2865_/Q VGND VGND VPWR VPWR _1449_/A sky130_fd_sc_hd__o21ai_1
XFILLER_28_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1377_ _1307_/X _1308_/X _2765_/Q VGND VGND VPWR VPWR _1377_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__1499__D1 _1498_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1502__A2 _1444_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2463__B1 _2456_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1671__D1 input80/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2940__D _2940_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2782__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2014__B _2054_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1741__A2 _1738_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2454__B1 _1716_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2206__B1 _2201_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2850__D _2850_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2205__A _2205_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output182_A _2038_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2509__A1 _2834_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1732__A2 _2207_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2280_ _2280_/A VGND VGND VPWR VPWR _2723_/D sky130_fd_sc_hd__clkbuf_1
X_1300_ _2872_/Q _1437_/A _1299_/Y VGND VGND VPWR VPWR _1300_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_1_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1496__A1 _2389_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2445__B1 _2444_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1995_ _2722_/Q input37/X _2034_/S VGND VGND VPWR VPWR _2277_/B sky130_fd_sc_hd__mux2_1
XANTENNA__2760__D _2760_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2616_ _2616_/A _2616_/B VGND VGND VPWR VPWR _2909_/D sky130_fd_sc_hd__nand2_1
XANTENNA__1954__A _2065_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2547_ _2858_/Q _2540_/X _1855_/X _2531_/X VGND VGND VPWR VPWR _2858_/D sky130_fd_sc_hd__o211a_1
XFILLER_47_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2478_ _2510_/A VGND VGND VPWR VPWR _2525_/B sky130_fd_sc_hd__clkbuf_4
X_1429_ _1429_/A VGND VGND VPWR VPWR _1454_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_56_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2935__D _2935_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1487__A1 _2389_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2670__D _2670_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2025__A _2324_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2678__CLK _2901_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1714__A2 _1713_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input39_A cpu_dat_i[13] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1478__A1 input72/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2845__D _2845_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1951__A2_N _1933_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1650__A1 _1635_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1780_ _1807_/A VGND VGND VPWR VPWR _1853_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__1402__A1 _2395_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2401_ _2401_/A _2401_/B _2401_/C VGND VGND VPWR VPWR _2402_/A sky130_fd_sc_hd__and3_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2363__C1 _2386_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2332_ _2332_/A _2332_/B _2337_/C VGND VGND VPWR VPWR _2333_/A sky130_fd_sc_hd__and3_1
XFILLER_57_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2263_ _2263_/A VGND VGND VPWR VPWR _2716_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2194_ _2194_/A _2194_/B VGND VGND VPWR VPWR _2195_/A sky130_fd_sc_hd__or2_1
XFILLER_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2755__D _2755_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2418__B1 _1581_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1949__A _2364_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1641__A1 _1620_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1387__C _1387_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1978_ _2824_/Q _1961_/X _1977_/X VGND VGND VPWR VPWR _1978_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2820__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2409__B1 _2537_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1859__A _1859_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2051__A2_N _2018_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2188__A2 _1665_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1594__A _1740_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_22_CLK_A clkbuf_opt_2_1_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output145_A _1873_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1320__B1 _1422_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1901_ _1901_/A VGND VGND VPWR VPWR _1901_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2881_ _2881_/CLK _2881_/D VGND VGND VPWR VPWR _2881_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1623__A1 _1618_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1832_ _2109_/A _1865_/B _2342_/A VGND VGND VPWR VPWR _1832_/X sky130_fd_sc_hd__or3_1
XANTENNA__2843__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1763_ _1707_/A _1689_/A _2807_/Q VGND VGND VPWR VPWR _1763_/X sky130_fd_sc_hd__o21a_1
X_1694_ _1691_/Y _1693_/Y _1679_/X VGND VGND VPWR VPWR _1694_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__2112__B _2625_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2315_ _2320_/A _2315_/B _2305_/X VGND VGND VPWR VPWR _2316_/A sky130_fd_sc_hd__or3b_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ _2246_/A VGND VGND VPWR VPWR _2709_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2177_ _2177_/A _2194_/B VGND VGND VPWR VPWR _2178_/A sky130_fd_sc_hd__or2_1
XANTENNA__1311__B1 _1309_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1679__A _1702_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1862__A1 _1807_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1862__B2 _2929_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1614__A1 _2171_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1398__B _1429_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1378__B1 _1377_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2303__A _2303_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1845__C _2346_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2575__C1 _1351_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput103 spi_dat_i[7] VGND VGND VPWR VPWR _1611_/D1 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1550__B1 _1549_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2395__D _2395_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2716__CLK _2745_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1998__A1_N _2897_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1605__A1 _2152_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2866__CLK _2880_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1369__B1 _1368_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2213__A _2213_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2566__C1 _2558_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2030__A1 _2832_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2100_ _2844_/Q _1814_/X _2099_/X VGND VGND VPWR VPWR _2100_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2031_ _2902_/Q _2000_/X _1975_/X _2030_/Y VGND VGND VPWR VPWR _2609_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_47_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1844__A1 input31/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1534__C_N input73/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2933_ _2946_/CLK _2933_/D VGND VGND VPWR VPWR _2933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2107__B _2624_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2864_ _2880_/CLK _2864_/D VGND VGND VPWR VPWR _2864_/Q sky130_fd_sc_hd__dfxtp_1
X_1815_ _1815_/A VGND VGND VPWR VPWR _2114_/A sky130_fd_sc_hd__clkbuf_2
X_2795_ _2839_/CLK _2795_/D VGND VGND VPWR VPWR _2795_/Q sky130_fd_sc_hd__dfxtp_1
X_1746_ _2211_/A _2211_/B _1702_/X VGND VGND VPWR VPWR _1746_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__2572__A2 _2358_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1677_ _1651_/X _1663_/X _1637_/X _1638_/X input81/X VGND VGND VPWR VPWR _1677_/Y
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA__1962__A _2114_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2739__CLK _2745_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2229_ _2235_/A VGND VGND VPWR VPWR _2415_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_42_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1835__A1 _1830_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2889__CLK _2920_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2943__D _2943_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2017__B _2605_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2033__A _2033_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1872__A _1878_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1771__B1 _1630_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1294__D _1367_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input21_A cpu_adr_i[27] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2079__A1 _2840_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2208__A _2208_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2853__D _2853_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output108_A _1473_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1600_ _1599_/X _1569_/X _2677_/Q VGND VGND VPWR VPWR _2167_/B sky130_fd_sc_hd__o21ai_1
XFILLER_9_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2580_ _2580_/A VGND VGND VPWR VPWR _2650_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1782__A _1807_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1531_ _1531_/A VGND VGND VPWR VPWR _1698_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1762__B1 _1739_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2597__B _2605_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1462_ _1803_/B _1803_/C _1462_/C _1462_/D VGND VGND VPWR VPWR _1528_/B sky130_fd_sc_hd__nand4_4
X_1393_ _1389_/Y _1287_/X _1392_/Y VGND VGND VPWR VPWR _2556_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__1514__B1 _2811_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2014_ _2014_/A _2054_/B _2284_/A VGND VGND VPWR VPWR _2014_/X sky130_fd_sc_hd__or3_1
XFILLER_24_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2763__D _2763_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2916_ _2920_/CLK _2916_/D VGND VGND VPWR VPWR _2916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1450__C1 _1508_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2847_ _2847_/CLK _2847_/D VGND VGND VPWR VPWR _2847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2778_ _2816_/CLK _2778_/D VGND VGND VPWR VPWR _2778_/Q sky130_fd_sc_hd__dfxtp_1
X_1729_ _1735_/A VGND VGND VPWR VPWR _1729_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__1692__A _1692_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1753__B1 _2805_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2938__D _2938_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1505__B1 _1504_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2673__D _2673_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1284__A2 _1372_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1441__C1 _1444_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2904__CLK _2915_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1992__B1 _1975_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input69_A cpu_sel_i[2] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2536__A2 _2519_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2848__D _2848_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2472__A1 _2408_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2701_ _2703_/CLK _2701_/D VGND VGND VPWR VPWR _2701_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1432__C1 _1444_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2632_ _2632_/A _2632_/B VGND VGND VPWR VPWR _2923_/D sky130_fd_sc_hd__nand2_1
XANTENNA__2104__C _2320_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput204 _1980_/Y VGND VGND VPWR VPWR spi_dat_o[8] sky130_fd_sc_hd__buf_2
X_2563_ _2563_/A VGND VGND VPWR VPWR _2867_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2401__A _2401_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1514_ _1463_/Y _2527_/A _2811_/Q VGND VGND VPWR VPWR _1515_/A sky130_fd_sc_hd__a21o_1
XANTENNA__2758__D _2758_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2494_ _2822_/Q _2493_/X _1965_/X _2488_/X VGND VGND VPWR VPWR _2822_/D sky130_fd_sc_hd__o211a_1
X_1445_ _1445_/A VGND VGND VPWR VPWR _1445_/X sky130_fd_sc_hd__buf_2
XFILLER_56_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1376_ _1376_/A VGND VGND VPWR VPWR _1436_/A sky130_fd_sc_hd__clkinv_2
XANTENNA__1499__C1 _1494_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2463__A1 _1748_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1671__C1 _1627_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2927__CLK _2930_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2014__C _2284_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1726__B1 _1679_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2311__A _2311_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2668__D _2668_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2454__A1 _2453_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2206__A1 _1724_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2509__A2 _2506_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output175_A _1993_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2221__A _2221_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2390__B1 _1455_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2142__B1 _1692_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1496__A2 _1452_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2445__A1 _2427_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1994_ _2058_/A VGND VGND VPWR VPWR _1994_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2615_ _2615_/A _2617_/B VGND VGND VPWR VPWR _2908_/D sky130_fd_sc_hd__nor2_1
XANTENNA__1708__B1 _2798_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2546_ _2546_/A VGND VGND VPWR VPWR _2857_/D sky130_fd_sc_hd__clkbuf_1
X_2477_ _2531_/A VGND VGND VPWR VPWR _2510_/A sky130_fd_sc_hd__buf_4
X_1428_ _1428_/A VGND VGND VPWR VPWR _1477_/A sky130_fd_sc_hd__buf_2
XFILLER_56_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2133__A0 _2247_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1487__A2 _1436_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1359_ _2864_/Q _1343_/X _1358_/Y VGND VGND VPWR VPWR _1423_/C sky130_fd_sc_hd__o21ai_1
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_opt_2_0_CLK_A clkbuf_1_0_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2306__A _2320_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2041__A _2078_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1880__A _1902_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2124__A0 _2241_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2861__D _2861_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2216__A _2216_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1650__A2 _1617_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1402__A2 _2395_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1938__B1 _1937_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2400_ _2400_/A VGND VGND VPWR VPWR _2775_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2363__B1 _1414_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2331_ _2331_/A VGND VGND VPWR VPWR _2744_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2262_ _2272_/A _2262_/B _2257_/X VGND VGND VPWR VPWR _2263_/A sky130_fd_sc_hd__or3b_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2115__B1 _2114_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2193_ _2193_/A _2193_/B VGND VGND VPWR VPWR _2194_/A sky130_fd_sc_hd__nand2_1
XANTENNA__2772__CLK _2776_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1323__D1 _2552_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2418__A1 _2412_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1949__B _1990_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2771__D _2771_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1641__A2 _1640_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1387__D _1387_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1977_ _2014_/A _1990_/B _2270_/A VGND VGND VPWR VPWR _1977_/X sky130_fd_sc_hd__or3_1
XANTENNA__1965__A _2014_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2529_ _2529_/A _2529_/B _2352_/X VGND VGND VPWR VPWR _2530_/A sky130_fd_sc_hd__or3b_1
XANTENNA__2946__D _2946_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2106__B1 _2058_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2409__A1 _2395_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2681__D _2681_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1875__A _1875_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input51_A cpu_dat_i[24] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2795__CLK _2839_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2856__D _2856_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output138_A _1615_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1320__A1 _1400_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1608__C1 _1595_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1900_ _1900_/A _2945_/Q VGND VGND VPWR VPWR _1901_/A sky130_fd_sc_hd__and2_1
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2880_ _2880_/CLK _2880_/D VGND VGND VPWR VPWR _2880_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1623__A2 _1622_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1831_ _2749_/Q input29/X _2108_/S VGND VGND VPWR VPWR _2342_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1762_ _1758_/X _1761_/Y _1739_/X _1740_/X VGND VGND VPWR VPWR _1762_/X sky130_fd_sc_hd__o211a_1
X_1693_ _1692_/X _1640_/X _2690_/Q VGND VGND VPWR VPWR _1693_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2314_ _2314_/A VGND VGND VPWR VPWR _2737_/D sky130_fd_sc_hd__clkbuf_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2111__A2_N _2064_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2245_ _2245_/A _2260_/B _2265_/C VGND VGND VPWR VPWR _2246_/A sky130_fd_sc_hd__and3_1
XANTENNA__2766__D _2766_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2176_ _2198_/A VGND VGND VPWR VPWR _2194_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1311__A1 _1301_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1862__A2 _2548_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1614__A2 _2171_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1398__C _1447_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2668__CLK _2670_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1378__A1 _1436_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2575__B1 _2554_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2303__B _2308_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput104 spi_dat_i[8] VGND VGND VPWR VPWR _1619_/D1 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1550__A1 _1537_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2676__D _2676_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1605__A2 _1543_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input99_A spi_dat_i[3] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1809__S _1860_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1369__A1 _1365_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2566__B1 _1381_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2030__A2 _2025_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1774__D1 input98/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2030_ _2832_/Q _2025_/X _2029_/X VGND VGND VPWR VPWR _2030_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2810__CLK _2881_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2932_ _2946_/CLK _2932_/D VGND VGND VPWR VPWR _2932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2863_ _2929_/CLK _2863_/D VGND VGND VPWR VPWR _2863_/Q sky130_fd_sc_hd__dfxtp_1
X_1814_ _2033_/A VGND VGND VPWR VPWR _1814_/X sky130_fd_sc_hd__buf_2
X_2794_ _2839_/CLK _2794_/D VGND VGND VPWR VPWR _2794_/Q sky130_fd_sc_hd__dfxtp_1
X_1745_ _1744_/X _1685_/X _2697_/Q VGND VGND VPWR VPWR _2211_/B sky130_fd_sc_hd__o21ai_1
XFILLER_8_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2572__A3 _2391_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1676_ _1635_/X _1617_/X _2794_/Q VGND VGND VPWR VPWR _1676_/X sky130_fd_sc_hd__o21a_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2228_ _1551_/Y _1482_/Y _1552_/Y _2386_/D _1572_/X VGND VGND VPWR VPWR _2704_/D
+ sky130_fd_sc_hd__o2111a_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1835__A2 _1824_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2159_ _2198_/A VGND VGND VPWR VPWR _2172_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_leaf_21_CLK_A clkbuf_1_0_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2314__A _2314_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1872__B _2932_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1771__A1 _1769_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2833__CLK _2901_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2079__A2 _2025_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input14_A cpu_adr_i[20] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2208__B _2216_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2224__A _2224_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1530_ _1913_/A VGND VGND VPWR VPWR _1530_/X sky130_fd_sc_hd__buf_2
XANTENNA__1762__A1 _1758_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1857__A2_N _1792_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1461_ _1461_/A _1511_/A _1461_/C VGND VGND VPWR VPWR _1462_/D sky130_fd_sc_hd__nor3_1
X_1392_ _2758_/Q _1428_/A _1391_/Y _1431_/A VGND VGND VPWR VPWR _1392_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_41_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1514__A1 _1463_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2013_ _2725_/Q input40/X _2013_/S VGND VGND VPWR VPWR _2284_/A sky130_fd_sc_hd__mux2_1
XANTENNA__1303__A _1400_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2915_ _2915_/CLK _2915_/D VGND VGND VPWR VPWR _2915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1450__B1 _1392_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2846_ _2881_/CLK _2846_/D VGND VGND VPWR VPWR _2846_/Q sky130_fd_sc_hd__dfxtp_1
X_2777_ _2881_/CLK _2777_/D VGND VGND VPWR VPWR _2777_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2706__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1728_ _1696_/X _1682_/X _2801_/Q VGND VGND VPWR VPWR _1728_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1753__A1 _1696_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1659_ _1599_/X _1612_/X _2685_/Q VGND VGND VPWR VPWR _2185_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__2856__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input6_A cpu_adr_i[13] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1505__A1 _1503_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1505__B2 _1327_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2466__C1 _2451_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2309__A _2309_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2044__A _2044_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1441__B1 _1440_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1992__B2 _1991_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1883__A _1889_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2219__A _2219_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output120_A _1574_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2864__D _2864_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2457__C1 _2451_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2472__A2 _2410_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1680__B1 _1679_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2700_ _2703_/CLK _2700_/D VGND VGND VPWR VPWR _2700_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2729__CLK _2834_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1432__B1 _1430_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2631_ _2631_/A _2631_/B VGND VGND VPWR VPWR _2922_/D sky130_fd_sc_hd__nor2_1
XANTENNA__1793__A _2092_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput205 _1988_/Y VGND VGND VPWR VPWR spi_dat_o[9] sky130_fd_sc_hd__buf_2
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2562_ _2573_/A _2562_/B _2415_/A VGND VGND VPWR VPWR _2563_/A sky130_fd_sc_hd__or3b_1
XFILLER_5_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2401__B _2401_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2879__CLK _2881_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1513_ _1513_/A VGND VGND VPWR VPWR _2527_/A sky130_fd_sc_hd__buf_2
X_2493_ _2493_/A VGND VGND VPWR VPWR _2493_/X sky130_fd_sc_hd__clkbuf_2
X_1444_ _1444_/A VGND VGND VPWR VPWR _1523_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__1499__B1 _1491_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1375_ _2867_/Q _1343_/X _1374_/Y VGND VGND VPWR VPWR _1387_/B sky130_fd_sc_hd__o21ai_1
XFILLER_55_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2774__D _2774_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1968__A _1980_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2463__A2 _1751_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1671__B1 _1626_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2829_ _2901_/CLK _2829_/D VGND VGND VPWR VPWR _2829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1726__A1 _1724_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2039__A _2039_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2684__D _2684_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1878__A _1878_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2454__A2 _2204_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1662__B1 _2792_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2206__A2 _1725_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input81_A spi_dat_i[16] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2859__D _2859_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output168_A _1835_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2390__A1 _2395_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2142__B2 _1859_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2142__A1 _1528_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2445__A2 _2428_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1653__B1 _2684_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1788__A _1803_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1993_ _2011_/A _2601_/A VGND VGND VPWR VPWR _1993_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1405__B1 _2877_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2614_ _2614_/A _2616_/B VGND VGND VPWR VPWR _2907_/D sky130_fd_sc_hd__nand2_1
XANTENNA__2412__A _2453_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2769__D _2769_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1708__A1 _1707_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2545_ _2548_/A _2545_/B _2537_/X VGND VGND VPWR VPWR _2546_/A sky130_fd_sc_hd__or3b_1
X_2476_ _1342_/A _1342_/B _1528_/B _2235_/A VGND VGND VPWR VPWR _2531_/A sky130_fd_sc_hd__o31a_4
X_1427_ _1815_/A _1426_/X _2867_/Q VGND VGND VPWR VPWR _1510_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__2133__A1 _2815_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1358_ _1362_/A _2368_/A _2368_/B VGND VGND VPWR VPWR _1358_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__1487__A3 _1452_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1289_ _1289_/A VGND VGND VPWR VPWR _1353_/A sky130_fd_sc_hd__buf_2
XFILLER_24_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1698__A _1698_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1644__B1 _2789_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2306__B _2306_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2322__A _2322_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2679__D _2679_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2041__B _2054_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1580__C1 _1556_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2124__A1 _2813_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1401__A _1401_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2216__B _2216_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1399__C1 _1431_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1938__A1 _2818_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2363__A1 _2757_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2330_ _2344_/A _2330_/B _2329_/X VGND VGND VPWR VPWR _2331_/A sky130_fd_sc_hd__or3b_1
X_2261_ _2261_/A VGND VGND VPWR VPWR _2715_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2917__CLK _2917_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2115__A1 _2847_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2192_ _1677_/Y _1678_/Y _2179_/X VGND VGND VPWR VPWR _2688_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__1323__C1 _1311_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2418__A2 _2164_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1949__C _2260_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1976_ _2719_/Q input65/X _2013_/S VGND VGND VPWR VPWR _2270_/A sky130_fd_sc_hd__mux2_1
XANTENNA__2051__B1 _1994_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1965__B _1990_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1981__A _2117_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2528_ _2528_/A VGND VGND VPWR VPWR _2848_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2106__B2 _2523_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2459_ _2447_/X _2448_/X _2458_/Y VGND VGND VPWR VPWR _2801_/D sky130_fd_sc_hd__o21ai_1
XFILLER_57_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2409__A2 _2395_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2317__A _2362_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2042__B1 _2041_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2052__A _2075_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1891__A _1902_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input44_A cpu_dat_i[18] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1856__B1 _1855_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1320__A2 _1401_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output200_A _1952_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2872__D _2872_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1608__B1 _1593_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2227__A _2227_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1830_ _1859_/A VGND VGND VPWR VPWR _1830_/X sky130_fd_sc_hd__clkbuf_2
X_1761_ _1759_/Y _1760_/Y _1630_/A VGND VGND VPWR VPWR _1761_/Y sky130_fd_sc_hd__a21oi_1
X_1692_ _1692_/A VGND VGND VPWR VPWR _1692_/X sky130_fd_sc_hd__clkbuf_2
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ _2313_/A _2332_/B _2313_/C VGND VGND VPWR VPWR _2314_/A sky130_fd_sc_hd__and3_1
XFILLER_44_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1306__A _1306_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ _2362_/A VGND VGND VPWR VPWR _2265_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_38_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1847__B1 _1840_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2175_ _2175_/A _2175_/B VGND VGND VPWR VPWR _2177_/A sky130_fd_sc_hd__nand2_1
XFILLER_54_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1311__A2 _1457_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1331__B1_N _2875_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2782__D _2782_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2137__A input1/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1398__D _1447_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1959_ _1980_/A _2595_/A VGND VGND VPWR VPWR _1959_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1378__A2 _1306_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2575__A1 _2878_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2303__C _2313_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2600__A _2600_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput105 spi_dat_i[9] VGND VGND VPWR VPWR _1628_/D1 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1550__A2 _1544_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1838__B1 _1789_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2692__D _2692_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2047__A _2047_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1886__A _1886_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2566__A1 _2357_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1369__A2 _1324_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2015__B1 _2014_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2762__CLK _2764_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1774__C1 _1710_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2510__A _2510_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1825__S _1860_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2867__D _2867_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output150_A _1884_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1829__B1 _2632_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2931_ _2946_/CLK _2931_/D VGND VGND VPWR VPWR _2931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1796__A _2019_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2862_ _2873_/CLK _2862_/D VGND VGND VPWR VPWR _2862_/Q sky130_fd_sc_hd__dfxtp_1
X_1813_ _2092_/A VGND VGND VPWR VPWR _2033_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__2556__C_N _2537_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2793_ _2839_/CLK _2793_/D VGND VGND VPWR VPWR _2793_/Q sky130_fd_sc_hd__dfxtp_1
X_1744_ _1744_/A VGND VGND VPWR VPWR _1744_/X sky130_fd_sc_hd__buf_4
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1675_ _1670_/X _1674_/Y _1667_/X _1668_/X VGND VGND VPWR VPWR _1675_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2777__D _2777_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ _2227_/A VGND VGND VPWR VPWR _2386_/D sky130_fd_sc_hd__buf_4
XFILLER_54_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2158_ _2158_/A _2158_/B VGND VGND VPWR VPWR _2160_/A sky130_fd_sc_hd__nand2_1
XFILLER_26_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2089_ _2842_/Q _1814_/X _2088_/X VGND VGND VPWR VPWR _2089_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_41_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2785__CLK _2816_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1771__A2 _1770_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_22_CLK clkbuf_opt_2_1_CLK/X VGND VGND VPWR VPWR _2768_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2330__A _2344_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2687__D _2687_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2505__A _2505_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2224__B _2224_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output198_A _2117_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1747__C1 _1740_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1762__A2 _1761_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1460_ _2862_/Q _1523_/A _1459_/Y VGND VGND VPWR VPWR _1511_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__2240__A _2251_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_13_CLK clkbuf_opt_3_0_CLK/X VGND VGND VPWR VPWR _2809_/CLK sky130_fd_sc_hd__clkbuf_16
X_1391_ input7/X _1429_/A _1447_/C _1447_/D VGND VGND VPWR VPWR _1391_/Y sky130_fd_sc_hd__nand4b_2
XANTENNA__1514__A2 _2527_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2012_ _2076_/A VGND VGND VPWR VPWR _2044_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2914_ _2920_/CLK _2914_/D VGND VGND VPWR VPWR _2914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2415__A _2415_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1450__A1 _1389_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2845_ _2847_/CLK _2845_/D VGND VGND VPWR VPWR _2845_/Q sky130_fd_sc_hd__dfxtp_1
X_2776_ _2776_/CLK _2776_/D VGND VGND VPWR VPWR _2776_/Q sky130_fd_sc_hd__dfxtp_1
X_1727_ _1722_/X _1726_/Y _1704_/X _1705_/X VGND VGND VPWR VPWR _1727_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2150__A _2647_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1658_ _1645_/X _1657_/X _1626_/X _1627_/X input78/X VGND VGND VPWR VPWR _2185_/A
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA__1753__A2 _1689_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1979__A2_N _1933_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1589_ _1576_/X _1588_/X _1533_/X _1536_/X _1589_/D1 VGND VGND VPWR VPWR _1589_/Y
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA__1505__A2 _1299_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2466__B1 _2456_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2218__B1 _2201_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2325__A _2344_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2044__B _2611_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1441__A1 _2769_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1883__B _2937_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2060__A _2094_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2800__CLK _2809_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2219__B _2219_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2457__B1 _2456_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output113_A _1661_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1680__A1 _1677_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_2_CLK clkbuf_1_0_0_CLK/X VGND VGND VPWR VPWR _2925_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2880__D _2880_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2235__A _2235_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1432__A1 _2762_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2630_ _2632_/A _2630_/B VGND VGND VPWR VPWR _2921_/D sky130_fd_sc_hd__nand2_1
Xoutput206 _2122_/Y VGND VGND VPWR VPWR spi_sel_o[0] sky130_fd_sc_hd__buf_2
X_2561_ _2357_/X _2358_/X _2375_/A _1492_/Y _2558_/X VGND VGND VPWR VPWR _2866_/D
+ sky130_fd_sc_hd__o311a_1
X_2492_ _2492_/A _2495_/B VGND VGND VPWR VPWR _2821_/D sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_20_CLK_A clkbuf_1_0_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1512_ _1512_/A _1512_/B _1512_/C _1512_/D VGND VGND VPWR VPWR _1513_/A sky130_fd_sc_hd__nand4_2
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2401__C _2401_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1443_ _1443_/A _2562_/B _1443_/C VGND VGND VPWR VPWR _1803_/C sky130_fd_sc_hd__nor3_4
XFILLER_4_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1499__A1 _1486_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1374_ _2377_/B _2377_/C _1437_/A VGND VGND VPWR VPWR _1374_/Y sky130_fd_sc_hd__nand3_1
XFILLER_55_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1314__A _1353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1968__B _2597_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1671__A1 _1645_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2790__D _2790_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2145__A _2235_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2828_ _2847_/CLK _2828_/D VGND VGND VPWR VPWR _2828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2823__CLK _2901_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2759_ _2768_/CLK _2759_/D VGND VGND VPWR VPWR _2759_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1726__A2 _1725_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2439__B1 _2438_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1878__B _2935_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1662__A1 _1635_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1894__A _1900_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input74_A spi_dat_i[0] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2390__A2 _1409_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2142__A2 _1528_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2875__D _2875_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1653__A1 _1620_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1788__B _1788_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1992_ _2896_/Q _1933_/X _1975_/X _1991_/Y VGND VGND VPWR VPWR _2601_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_14_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1405__A1 _1379_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2846__CLK _2881_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2613_ _2613_/A _2617_/B VGND VGND VPWR VPWR _2906_/D sky130_fd_sc_hd__nor2_1
X_2544_ _2856_/Q _2540_/X _1845_/X _2531_/X VGND VGND VPWR VPWR _2856_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1708__A2 _1689_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2475_ _2493_/A VGND VGND VPWR VPWR _2475_/X sky130_fd_sc_hd__clkbuf_2
X_1426_ _1488_/A VGND VGND VPWR VPWR _1426_/X sky130_fd_sc_hd__buf_2
XFILLER_29_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1357_ _1307_/X _1308_/X _2759_/Q VGND VGND VPWR VPWR _2368_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__2785__D _2785_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1288_ _1343_/A VGND VGND VPWR VPWR _1437_/A sky130_fd_sc_hd__buf_2
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1644__A1 _1624_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2603__A _2603_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2322__B _2332_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2041__C _2294_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1580__B1 _1473_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2695__D _2695_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2719__CLK _2745_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1332__B1 _1331_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1889__A _1889_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2869__CLK _2873_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2096__A1_N _2913_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1399__B1 _1398_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2513__A _2513_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1938__A2 _2353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output180_A _2024_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2363__A2 _1785_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2260_ _2260_/A _2260_/B _2265_/C VGND VGND VPWR VPWR _2261_/A sky130_fd_sc_hd__and3_1
XFILLER_38_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2115__A2 _2251_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2191_ _2191_/A VGND VGND VPWR VPWR _2687_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1323__B1 _1300_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2520__C1 _2514_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1799__A _2027_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1975_ _2058_/A VGND VGND VPWR VPWR _1975_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2051__B2 _2511_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1965__C _2265_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2527_ _2527_/A _2527_/B _2653_/C VGND VGND VPWR VPWR _2528_/A sky130_fd_sc_hd__and3_1
X_2458_ _2453_/X _2208_/A _1728_/X VGND VGND VPWR VPWR _2458_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1409_ _1409_/A _1409_/B VGND VGND VPWR VPWR _1411_/A sky130_fd_sc_hd__nand2_1
XFILLER_60_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2389_ _2389_/A VGND VGND VPWR VPWR _2395_/B sky130_fd_sc_hd__buf_2
XFILLER_56_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2333__A _2333_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2578__C1 _2382_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2042__A1 _2834_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2052__B _2612_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1553__B1 _1552_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input37_A cpu_dat_i[11] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2502__C1 _2501_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2691__CLK _2839_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1856__A1 _2858_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2508__A _2508_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1608__A1 _1603_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1760_ _1567_/X _1712_/X _2700_/Q VGND VGND VPWR VPWR _1760_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2243__A _2243_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1691_ _1651_/X _1663_/X _1637_/X _1638_/X input83/X VGND VGND VPWR VPWR _1691_/Y
+ sky130_fd_sc_hd__o2111ai_2
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1544__B1 _2672_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2312_ _2312_/A VGND VGND VPWR VPWR _2332_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_39_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2243_ _2243_/A VGND VGND VPWR VPWR _2362_/A sky130_fd_sc_hd__buf_2
XFILLER_54_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1847__B2 _1846_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2174_ _1619_/Y _1621_/Y _2156_/X VGND VGND VPWR VPWR _2680_/D sky130_fd_sc_hd__a21oi_1
XFILLER_54_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2153__A _2153_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1958_ _2891_/Q _1953_/X _1927_/X _2492_/A VGND VGND VPWR VPWR _2595_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2575__A2 _2493_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1889_ _1889_/A _2940_/Q VGND VGND VPWR VPWR _1890_/A sky130_fd_sc_hd__and2_1
XANTENNA__2600__B _2604_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput106 spi_err_i VGND VGND VPWR VPWR _1534_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1838__B2 _2925_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1838__A1 _1807_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2328__A _2328_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1453__B1_N _2771_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2063__A _2075_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2907__CLK _2915_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2015__A1 _2830_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2566__A2 _2358_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1774__B1 _1709_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2002__S _2013_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1407__A _2876_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1526__B1 _1493_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output143_A _1868_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1829__A1 _1779_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2883__D _2883_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2238__A _2238_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2930_ _2930_/CLK _2930_/D VGND VGND VPWR VPWR _2930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2861_ _2881_/CLK _2861_/D VGND VGND VPWR VPWR _2861_/Q sky130_fd_sc_hd__dfxtp_1
X_1812_ _1779_/X _1781_/X _2630_/B VGND VGND VPWR VPWR _1812_/Y sky130_fd_sc_hd__a21oi_2
X_2792_ _2847_/CLK _2792_/D VGND VGND VPWR VPWR _2792_/Q sky130_fd_sc_hd__dfxtp_1
X_1743_ _1717_/X _1729_/X _1698_/X _1699_/X input91/X VGND VGND VPWR VPWR _2211_/A
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_7_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1765__B1 _2701_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1674_ _2189_/A _2189_/B _1630_/X VGND VGND VPWR VPWR _1674_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1317__A _1354_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ _2537_/A VGND VGND VPWR VPWR _2227_/A sky130_fd_sc_hd__buf_4
XFILLER_54_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2793__D _2793_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2148__A _2148_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2157_ _1537_/Y _1544_/Y _2156_/X VGND VGND VPWR VPWR _2672_/D sky130_fd_sc_hd__a21oi_1
XFILLER_26_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2088_ _2109_/A _2109_/B _2313_/A VGND VGND VPWR VPWR _2088_/X sky130_fd_sc_hd__or3_2
XFILLER_41_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2611__A _2611_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1756__B1 _1702_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2330__B _2330_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2058__A _2058_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1897__A _1897_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2505__B _2508_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1995__A0 _2722_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2521__A _2521_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1836__S _1860_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1747__B1 _1739_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2878__D _2878_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1390_ _1390_/A VGND VGND VPWR VPWR _1428_/A sky130_fd_sc_hd__buf_2
X_2011_ _2011_/A _2604_/A VGND VGND VPWR VPWR _2011_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2913_ _2915_/CLK _2913_/D VGND VGND VPWR VPWR _2913_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1986__B1 _1985_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1450__A2 _1523_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2844_ _2881_/CLK _2844_/D VGND VGND VPWR VPWR _2844_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_9_CLK_A clkbuf_1_1_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1738__B1 _1679_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2775_ _2880_/CLK _2775_/D VGND VGND VPWR VPWR _2775_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2431__A _2451_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1726_ _1724_/Y _1725_/Y _1679_/X VGND VGND VPWR VPWR _1726_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_7_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2788__D _2788_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2150__B _2670_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1657_ _1735_/A VGND VGND VPWR VPWR _1657_/X sky130_fd_sc_hd__clkbuf_4
X_1588_ _1913_/A VGND VGND VPWR VPWR _1588_/X sky130_fd_sc_hd__buf_2
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2209_ _2209_/A VGND VGND VPWR VPWR _2695_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2752__CLK _2873_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2466__A1 _1758_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2218__A1 _1759_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2606__A _2618_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1510__A _1510_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2325__B _2325_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1441__A2 _1477_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2341__A _2374_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2698__D _2698_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2060__B _2072_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2154__B1 _2235_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2457__A1 _1722_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2516__A _2516_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1680__A2 _1678_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1420__A _1447_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1432__A2 _1477_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput207 _2126_/Y VGND VGND VPWR VPWR spi_sel_o[1] sky130_fd_sc_hd__buf_2
XFILLER_5_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2393__B1 _2772_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2251__A _2251_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2560_ _2577_/A _2560_/B VGND VGND VPWR VPWR _2865_/D sky130_fd_sc_hd__nand2_1
X_2491_ _2820_/Q _2475_/X _1949_/X _2488_/X VGND VGND VPWR VPWR _2820_/D sky130_fd_sc_hd__o211a_1
X_1511_ _1511_/A _2573_/B _1511_/C VGND VGND VPWR VPWR _1512_/D sky130_fd_sc_hd__nor3_1
XFILLER_4_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1442_ _1442_/A _1442_/B _1510_/C _1510_/D VGND VGND VPWR VPWR _1443_/C sky130_fd_sc_hd__nand4_2
X_1373_ _1451_/A _1452_/A _2762_/Q VGND VGND VPWR VPWR _2377_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__2775__CLK _2880_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1499__A2 _1487_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1314__B _1354_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1671__A2 _1657_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1330__A _1414_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2827_ _2901_/CLK _2827_/D VGND VGND VPWR VPWR _2827_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2161__A _2161_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2758_ _2776_/CLK _2758_/D VGND VGND VPWR VPWR _2758_/Q sky130_fd_sc_hd__dfxtp_1
X_1709_ _1709_/A VGND VGND VPWR VPWR _1709_/X sky130_fd_sc_hd__buf_2
XFILLER_63_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2689_ _2839_/CLK _2689_/D VGND VGND VPWR VPWR _2689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2439__A1 _2427_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2336__A _2526_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1662__A2 _1617_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1894__B _2942_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input67_A cpu_sel_i[0] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1583__D1 input99/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2390__A3 _1452_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2798__CLK _2840_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2127__A0 _2709_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2891__D _2891_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1653__A2 _1640_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1788__C _1803_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2246__A _2246_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1991_ _2826_/Q _1961_/X _1990_/X VGND VGND VPWR VPWR _1991_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_9_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1405__A2 _1488_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2612_ _2612_/A _2616_/B VGND VGND VPWR VPWR _2905_/D sky130_fd_sc_hd__nand2_1
XFILLER_9_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2543_ _2543_/A VGND VGND VPWR VPWR _2855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2118__A0 _2707_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2474_ _2474_/A VGND VGND VPWR VPWR _2493_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__1325__A _1325_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1425_ _1445_/A VGND VGND VPWR VPWR _1815_/A sky130_fd_sc_hd__buf_2
X_1356_ _1447_/C _1447_/D input8/X _1429_/A VGND VGND VPWR VPWR _2368_/A sky130_fd_sc_hd__nand4_2
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1287_ _1335_/C VGND VGND VPWR VPWR _1287_/X sky130_fd_sc_hd__buf_4
XFILLER_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2156__A _2224_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1644__A2 _1609_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2241__C_N _2227_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2603__B _2605_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2940__CLK _2946_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2322__C _2337_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1580__A1 _1575_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1332__A1 _1329_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1889__B _2940_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1399__A1 _2772_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2513__B _2521_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output173_A _2949_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1844__S _2127_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2886__D _2886_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2016__A2_N _2000_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2190_ _2190_/A _2194_/B VGND VGND VPWR VPWR _2191_/A sky130_fd_sc_hd__or2_1
XANTENNA__1323__A1 _2879_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2520__B1 _2088_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2813__CLK _2925_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1974_ _1980_/A _2598_/A VGND VGND VPWR VPWR _1974_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2526_ _2526_/A VGND VGND VPWR VPWR _2653_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__2796__D _2796_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2457_ _1722_/X _1726_/Y _2456_/X _2451_/X VGND VGND VPWR VPWR _2800_/D sky130_fd_sc_hd__o211a_1
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1408_ _1379_/X _1380_/A _1407_/Y VGND VGND VPWR VPWR _1408_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2388_ _2366_/B _1330_/C _2366_/A _1329_/X _2365_/Y VGND VGND VPWR VPWR _2770_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_21_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1339_ _2382_/B _2382_/C _1343_/A VGND VGND VPWR VPWR _1339_/Y sky130_fd_sc_hd__nand3_4
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2614__A _2614_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2578__B1 _1490_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2042__A2 _2025_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1553__A1 _1551_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2502__B1 _2003_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2836__CLK _2840_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1856__A2 _1841_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2508__B _2508_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1608__A2 _1607_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2569__B1 _2552_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1690_ _1635_/X _1689_/X _2796_/Q VGND VGND VPWR VPWR _1690_/X sky130_fd_sc_hd__o21a_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1544__A1 _2152_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2311_ _2311_/A VGND VGND VPWR VPWR _2736_/D sky130_fd_sc_hd__clkbuf_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2242_ _2242_/A VGND VGND VPWR VPWR _2708_/D sky130_fd_sc_hd__clkbuf_1
X_2173_ _2173_/A VGND VGND VPWR VPWR _2679_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1480__A0 _2327_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1957_ _2821_/Q _2474_/A _1956_/X VGND VGND VPWR VPWR _2492_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__2709__CLK _2776_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1888_ _1888_/A VGND VGND VPWR VPWR _1888_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2080__A1_N _2910_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2859__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2509_ _2834_/Q _2506_/X _2041_/X _2501_/X VGND VGND VPWR VPWR _2834_/D sky130_fd_sc_hd__o211a_1
Xinput107 spi_rty_i VGND VGND VPWR VPWR _1534_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2609__A _2609_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1838__A2 _2542_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2496__C1 _2488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1513__A _1513_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1471__B1 _1470_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2344__A _2344_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2063__B _2614_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1759__D1 input94/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2015__A2 _1961_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1774__A1 _1723_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2566__A3 _2380_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2420__C1 _2405_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1526__A1 _1490_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1526__B2 _1339_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1829__A2 _1824_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output136_A _1602_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2519__A _2540_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1423__A _1423_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2238__B _2260_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2860_ _2929_/CLK _2860_/D VGND VGND VPWR VPWR _2860_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2254__A _2254_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1811_ _1807_/X _2534_/B _1789_/X _2921_/Q VGND VGND VPWR VPWR _2630_/B sky130_fd_sc_hd__o22ai_2
XFILLER_50_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2791_ _2839_/CLK _2791_/D VGND VGND VPWR VPWR _2791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1765__A1 _1744_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2411__C1 _1469_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1742_ _1696_/X _1682_/X _2803_/Q VGND VGND VPWR VPWR _1742_/X sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_1_1_0_CLK_A clkbuf_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1673_ _1672_/X _1612_/X _2687_/Q VGND VGND VPWR VPWR _2189_/B sky130_fd_sc_hd__o21ai_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ _2225_/A VGND VGND VPWR VPWR _2703_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1333__A _1333_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2156_ _2224_/B VGND VGND VPWR VPWR _2156_/X sky130_fd_sc_hd__buf_2
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2087_ _2737_/Q input53/X _2108_/S VGND VGND VPWR VPWR _2313_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2164__A _2164_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2611__B _2617_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1756__A1 _2215_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2681__CLK _2901_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2103__S _2113_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1508__A _1508_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2469__C1 _2451_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2339__A _2344_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2325__C_N _2305_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1995__A1 input37/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input97_A spi_dat_i[30] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2521__B _2521_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1747__A1 _1742_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2013__S _2013_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2894__D _2894_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2249__A _2249_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2010_ _2899_/Q _1953_/X _1994_/X _2503_/A VGND VGND VPWR VPWR _2604_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1683__B1 _2795_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2912_ _2917_/CLK _2912_/D VGND VGND VPWR VPWR _2912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1435__B1 _2870_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1986__A1 _2825_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2843_ _2847_/CLK _2843_/D VGND VGND VPWR VPWR _2843_/Q sky130_fd_sc_hd__dfxtp_1
X_2774_ _2776_/CLK _2774_/D VGND VGND VPWR VPWR _2774_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1738__A1 _1736_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1725_ _1692_/X _1712_/X _2694_/Q VGND VGND VPWR VPWR _1725_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2396__D1 _2395_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2150__C _2401_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1656_ _1624_/X _1609_/X _2791_/Q VGND VGND VPWR VPWR _1656_/X sky130_fd_sc_hd__o21a_1
X_1587_ _1517_/X _1519_/X _2782_/Q VGND VGND VPWR VPWR _1587_/X sky130_fd_sc_hd__o21a_1
XFILLER_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2159__A _2198_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2208_ _2208_/A _2216_/B VGND VGND VPWR VPWR _2209_/A sky130_fd_sc_hd__or2_1
XANTENNA__2348__C_N _2329_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2466__A2 _1761_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2139_ _2580_/A VGND VGND VPWR VPWR _2639_/B sky130_fd_sc_hd__buf_2
XFILLER_26_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1674__B1 _1630_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2218__A2 _1760_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1510__B _1510_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2622__A _2622_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2387__D1 _2382_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2060__C _2301_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2154__A1 _1696_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2457__A2 _1726_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1665__B1 _2686_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input12_A cpu_adr_i[19] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2516__B _2521_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2090__B1 _2039_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2889__D _2889_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput208 _2131_/Y VGND VGND VPWR VPWR spi_sel_o[2] sky130_fd_sc_hd__buf_2
XFILLER_64_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2393__A1 _2395_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2490_ _2490_/A _2495_/B VGND VGND VPWR VPWR _2819_/D sky130_fd_sc_hd__nand2_1
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1510_ _1510_/A _1510_/B _1510_/C _1510_/D VGND VGND VPWR VPWR _1511_/C sky130_fd_sc_hd__nand4_1
X_1441_ _2769_/Q _1477_/A _1440_/Y _1444_/A VGND VGND VPWR VPWR _1510_/D sky130_fd_sc_hd__o211ai_2
XFILLER_4_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1372_ _1372_/A VGND VGND VPWR VPWR _1452_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__1656__B1 _2791_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1330__B _1414_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1408__B1 _1407_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2826_ _2847_/CLK _2826_/D VGND VGND VPWR VPWR _2826_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2799__D _2799_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2757_ _2764_/CLK _2757_/D VGND VGND VPWR VPWR _2757_/Q sky130_fd_sc_hd__dfxtp_1
X_2688_ _2839_/CLK _2688_/D VGND VGND VPWR VPWR _2688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1708_ _1707_/X _1689_/X _2798_/Q VGND VGND VPWR VPWR _1708_/X sky130_fd_sc_hd__o21a_1
X_1639_ _1576_/X _1588_/X _1637_/X _1638_/X input75/X VGND VGND VPWR VPWR _1639_/Y
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input4_A cpu_adr_i[11] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2439__A2 _2428_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2617__A _2617_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1647__B1 _2683_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1521__A _1717_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2352__A _2352_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1583__C1 _1565_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2127__A1 input69/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_8_CLK_A clkbuf_1_1_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1431__A _1431_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2527__A _2527_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1990_ _2014_/A _1990_/B _2274_/A VGND VGND VPWR VPWR _1990_/X sky130_fd_sc_hd__or3_1
XFILLER_60_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1810__A0 _2334_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2262__A _2272_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2611_ _2611_/A _2617_/B VGND VGND VPWR VPWR _2904_/D sky130_fd_sc_hd__nor2_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2542_ _2548_/A _2542_/B _2537_/X VGND VGND VPWR VPWR _2543_/A sky130_fd_sc_hd__or3b_1
XANTENNA__2742__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1574__C1 _1556_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1606__A _1702_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2118__A1 input67/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2473_ _2395_/B _2395_/D _2231_/A _2366_/B _1470_/Y VGND VGND VPWR VPWR _2811_/D
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__2892__CLK _2917_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1424_ _1424_/A VGND VGND VPWR VPWR _1445_/A sky130_fd_sc_hd__buf_2
XANTENNA__1325__B _1390_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1355_ _1355_/A VGND VGND VPWR VPWR _1429_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1629__B1 _2681_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1286_ _1343_/A VGND VGND VPWR VPWR _1335_/C sky130_fd_sc_hd__buf_2
XFILLER_36_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1341__A _1341_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2172__A _2172_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2809_ _2809_/CLK _2809_/D VGND VGND VPWR VPWR _2809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1580__A2 _1579_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1516__A _1696_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1868__B1 _2639_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1332__A2 _1479_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2347__A _2347_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2765__CLK _2768_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1399__A2 _1428_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output166_A _1823_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1426__A _1488_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1323__A2 _1287_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2520__A1 _2842_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1860__S _1860_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2257__A _2352_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1973_ _2893_/Q _1953_/X _1927_/X _2495_/A VGND VGND VPWR VPWR _2598_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__2036__B1 _2035_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2525_ _2525_/A _2525_/B VGND VGND VPWR VPWR _2847_/D sky130_fd_sc_hd__nand2_1
X_2456_ _2558_/A VGND VGND VPWR VPWR _2456_/X sky130_fd_sc_hd__clkbuf_4
X_1407_ _2876_/Q VGND VGND VPWR VPWR _1407_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2387_ _2769_/Q _1785_/S _1440_/Y _2386_/D _2382_/A VGND VGND VPWR VPWR _2769_/D
+ sky130_fd_sc_hd__o2111a_1
X_1338_ _1296_/X _1372_/A _2766_/Q VGND VGND VPWR VPWR _2382_/C sky130_fd_sc_hd__o21ai_2
XFILLER_56_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2167__A _2167_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2788__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2614__B _2616_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2578__A1 _2401_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2630__A _2632_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1553__A2 _1482_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2502__A1 _2828_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2569__A1 _1504_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1777__C1 _1633_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2540__A _2540_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2897__D _2897_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1544__A2 _1543_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2310_ _2320_/A _2310_/B _2305_/X VGND VGND VPWR VPWR _2311_/A sky130_fd_sc_hd__or3b_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2241_ _2540_/A _2241_/B _2227_/A VGND VGND VPWR VPWR _2242_/A sky130_fd_sc_hd__or3b_1
XFILLER_39_926 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2172_ _2172_/A _2172_/B VGND VGND VPWR VPWR _2173_/A sky130_fd_sc_hd__or2_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2930__CLK _2930_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2009__B1 _2008_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1480__A1 _2848_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1956_ _1971_/A _2008_/B _2262_/B VGND VGND VPWR VPWR _1956_/X sky130_fd_sc_hd__or3_2
X_1887_ _1889_/A _2939_/Q VGND VGND VPWR VPWR _1888_/A sky130_fd_sc_hd__and2_1
XANTENNA__2062__A2_N _2018_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2508_ _2508_/A _2508_/B VGND VGND VPWR VPWR _2833_/D sky130_fd_sc_hd__nand2_1
X_2439_ _2427_/X _2428_/X _2438_/Y VGND VGND VPWR VPWR _2791_/D sky130_fd_sc_hd__o21ai_1
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2609__B _2617_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2496__B1 _1977_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2625__A _2625_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1471__A1 _2395_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2344__B _2344_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1759__C1 _1710_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2420__B1 _2416_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1774__A2 _1729_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2360__A _2665_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2803__CLK _2809_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1526__A2 _1335_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input42_A cpu_dat_i[16] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1704__A _1739_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1423__B _1508_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2238__C _2386_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output129_A _1762_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2535__A _2535_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2254__B _2260_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1810_ _2334_/B _2851_/Q _2374_/A VGND VGND VPWR VPWR _2534_/B sky130_fd_sc_hd__mux2_1
XFILLER_62_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2790_ _2847_/CLK _2790_/D VGND VGND VPWR VPWR _2790_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2411__B1 _1545_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1741_ _1734_/X _1738_/Y _1739_/X _1740_/X VGND VGND VPWR VPWR _1741_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1765__A2 _1543_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1672_ _1744_/A VGND VGND VPWR VPWR _1672_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_16_CLK clkbuf_1_1_0_CLK/X VGND VGND VPWR VPWR _2745_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2270__A _2270_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ _2224_/A _2224_/B VGND VGND VPWR VPWR _2225_/A sky130_fd_sc_hd__or2_1
XFILLER_39_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2155_ _2198_/A VGND VGND VPWR VPWR _2224_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__1333__B _1390_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2086_ _2102_/A _2619_/A VGND VGND VPWR VPWR _2086_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2164__B _2172_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1453__A1 _2389_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2826__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1939_ _2888_/Q _1933_/X _1916_/X _1938_/Y VGND VGND VPWR VPWR _2591_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__1756__A2 _2215_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2277__C_N _2257_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput90 spi_dat_i[24] VGND VGND VPWR VPWR input90/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1508__B _1508_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2469__B1 _2456_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2339__B _2339_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1677__D1 input81/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2355__A _2355_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1747__A2 _1746_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1434__A _1488_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2249__B _2260_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_CLK clkbuf_1_0_0_CLK/X VGND VGND VPWR VPWR _2930_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1683__A1 _1624_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2265__A _2265_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2911_ _2915_/CLK _2911_/D VGND VGND VPWR VPWR _2911_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2849__CLK _2925_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1435__A1 _1815_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1986__A2 _1969_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2842_ _2881_/CLK _2842_/D VGND VGND VPWR VPWR _2842_/Q sky130_fd_sc_hd__dfxtp_1
X_2773_ _2776_/CLK _2773_/D VGND VGND VPWR VPWR _2773_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1430__A_N _1370_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1724_ _1723_/X _1663_/X _1709_/X _1710_/X input88/X VGND VGND VPWR VPWR _1724_/Y
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA__1738__A2 _1737_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1609__A _1682_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2396__C1 _2386_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1655_ _1650_/X _1654_/Y _1632_/X _1633_/X VGND VGND VPWR VPWR _1655_/X sky130_fd_sc_hd__o211a_1
X_1586_ _1581_/X _1585_/Y _1473_/X _1556_/X VGND VGND VPWR VPWR _1586_/X sky130_fd_sc_hd__o211a_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1344__A _1344_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2207_ _2207_/A _2207_/B VGND VGND VPWR VPWR _2208_/A sky130_fd_sc_hd__nand2_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2138_ _1744_/X _1543_/A _2537_/A VGND VGND VPWR VPWR _2580_/A sky130_fd_sc_hd__o21ai_2
XFILLER_27_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1674__A1 _2189_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2069_ _2908_/Q _2064_/X _2039_/X _2068_/Y VGND VGND VPWR VPWR _2615_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__2175__A _2175_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1510__C _1510_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2622__B _2626_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2387__C1 _2386_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1519__A _1682_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2154__A2 _1616_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1665__A1 _1620_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2090__B2 _2089_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output196_A _1940_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1429__A _1429_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2393__A2 _2395_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput209 _2135_/Y VGND VGND VPWR VPWR spi_sel_o[3] sky130_fd_sc_hd__buf_2
XFILLER_5_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1440_ _1440_/A _1454_/B _1454_/C _1454_/D VGND VGND VPWR VPWR _1440_/Y sky130_fd_sc_hd__nand4_1
X_1371_ _1371_/A VGND VGND VPWR VPWR _1451_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2550__C1 _2510_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2671__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1656__A1 _1624_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1330__C _1330_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1408__A1 _1379_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2825_ _2901_/CLK _2825_/D VGND VGND VPWR VPWR _2825_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1339__A _2382_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2756_ _2880_/CLK _2756_/D VGND VGND VPWR VPWR _2756_/Q sky130_fd_sc_hd__dfxtp_1
X_2687_ _2839_/CLK _2687_/D VGND VGND VPWR VPWR _2687_/Q sky130_fd_sc_hd__dfxtp_1
X_1707_ _1707_/A VGND VGND VPWR VPWR _1707_/X sky130_fd_sc_hd__clkbuf_2
X_1638_ _1710_/A VGND VGND VPWR VPWR _1638_/X sky130_fd_sc_hd__buf_2
XANTENNA__2315__C_N _2305_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1569_ _1712_/A VGND VGND VPWR VPWR _1569_/X sky130_fd_sc_hd__clkbuf_2
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2541__C1 _2531_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1647__A1 _1599_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2617__B _2617_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1948__S _2132_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2633__A _2633_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1583__B1 _1564_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2532__C1 _2531_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2694__CLK _2703_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1712__A _1712_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2527__B _2527_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output209_A _2135_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output111_A _1649_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2543__A _2543_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1810__A1 _2851_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2262__B _2262_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2610_ _2610_/A _2616_/B VGND VGND VPWR VPWR _2903_/D sky130_fd_sc_hd__nand2_1
XANTENNA__1466__B1_N _2705_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2541_ _2854_/Q _2540_/X _1832_/X _2531_/X VGND VGND VPWR VPWR _2854_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1574__B1 _1473_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2472_ _2408_/X _2410_/X _1556_/X VGND VGND VPWR VPWR _2810_/D sky130_fd_sc_hd__o21a_1
XFILLER_5_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1423_ _1423_/A _1508_/B _1423_/C _1508_/D VGND VGND VPWR VPWR _1803_/B sky130_fd_sc_hd__and4_2
XANTENNA__1326__B1 _2768_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1354_ _1354_/A VGND VGND VPWR VPWR _1447_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1285_ _1350_/A VGND VGND VPWR VPWR _1343_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__1629__A1 _1599_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1341__B _1341_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2453__A _2453_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2172__B _2172_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2808_ _2847_/CLK _2808_/D VGND VGND VPWR VPWR _2808_/Q sky130_fd_sc_hd__dfxtp_1
X_2739_ _2745_/CLK _2739_/D VGND VGND VPWR VPWR _2739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1868__A1 _1859_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2628__A _2632_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1332__A3 _1330_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1532__A _1698_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input107_A spi_rty_i VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input72_A cpu_we_i VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1707__A _1707_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output159_A _1901_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2538__A _2548_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2520__A2 _2519_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1442__A _1442_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2036__A1 _2833_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2273__A _2273_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1972_ _2823_/Q _1969_/X _1971_/X VGND VGND VPWR VPWR _2495_/A sky130_fd_sc_hd__o21ai_1
XFILLER_14_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1547__B1 _1546_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1617__A _1689_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2524_ _2846_/Q _2519_/X _2109_/X _2514_/X VGND VGND VPWR VPWR _2846_/D sky130_fd_sc_hd__o211a_1
X_2455_ _2447_/X _2448_/X _2454_/Y VGND VGND VPWR VPWR _2799_/D sky130_fd_sc_hd__o21ai_1
XFILLER_60_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2386_ _2386_/A _2386_/B _2386_/C _2386_/D VGND VGND VPWR VPWR _2768_/D sky130_fd_sc_hd__nand4_1
X_1406_ _1509_/B _1406_/B _1509_/A VGND VGND VPWR VPWR _1461_/C sky130_fd_sc_hd__nand3_2
XFILLER_60_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1337_ _1337_/A _1390_/A VGND VGND VPWR VPWR _2382_/B sky130_fd_sc_hd__nand2_2
XANTENNA__2448__A _2448_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2167__B _2167_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2183__A _2183_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2578__A2 _2358_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_leaf_7_CLK_A clkbuf_1_0_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2630__B _2630_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1527__A _1527_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2502__A2 _2493_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2358__A _2358_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2732__CLK _2834_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2882__CLK _2920_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2569__A2 _1327_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1777__B1 _1632_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1437__A _1437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ _2251_/A VGND VGND VPWR VPWR _2540_/A sky130_fd_sc_hd__buf_4
XFILLER_39_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1701__B1 _2691_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2171_ _2171_/A _2171_/B VGND VGND VPWR VPWR _2172_/A sky130_fd_sc_hd__nand2_1
XANTENNA__2268__A _2268_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1900__A _1900_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2009__A1 _2829_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1955_ _2716_/Q input62/X _1970_/S VGND VGND VPWR VPWR _2262_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1768__B1 _2808_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1886_ _1886_/A VGND VGND VPWR VPWR _1886_/X sky130_fd_sc_hd__clkbuf_1
X_2507_ _2832_/Q _2506_/X _2029_/X _2501_/X VGND VGND VPWR VPWR _2832_/D sky130_fd_sc_hd__o211a_1
X_2438_ _2433_/X _2186_/A _1656_/X VGND VGND VPWR VPWR _2438_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__2178__A _2178_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2755__CLK _2764_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2369_ _2526_/A VGND VGND VPWR VPWR _2391_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__2496__A1 _2824_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2625__B _2631_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1471__A2 _2366_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2641__A _2647_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1759__B1 _1709_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2420__A1 _1587_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2184__B1 _2179_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1931__B1 _1927_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input35_A cpu_dat_i[0] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2088__A _2109_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1423__C _1423_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1695__C1 _1668_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1998__B1 _1994_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2254__C _2265_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2411__B2 _1467_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2411__A1 _2706_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1740_ _1740_/A VGND VGND VPWR VPWR _1740_/X sky130_fd_sc_hd__clkbuf_2
X_1671_ _1645_/X _1657_/X _1626_/X _1627_/X input80/X VGND VGND VPWR VPWR _2189_/A
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA__2270__B _2284_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2701__D _2701_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2778__CLK _2816_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ _2223_/A _2223_/B VGND VGND VPWR VPWR _2224_/A sky130_fd_sc_hd__nand2_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2154_ _1696_/A _1616_/A _2235_/A VGND VGND VPWR VPWR _2198_/A sky130_fd_sc_hd__o21ai_4
XFILLER_38_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2085_ _2911_/Q _1914_/X _2058_/X _2518_/A VGND VGND VPWR VPWR _2619_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__1630__A _1630_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1989__A0 _2721_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1438__C1 _1500_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1453__A2 _1452_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1938_ _2818_/Q _2353_/A _1937_/X VGND VGND VPWR VPWR _1938_/Y sky130_fd_sc_hd__o21ai_1
X_1869_ _1902_/A VGND VGND VPWR VPWR _1878_/A sky130_fd_sc_hd__clkbuf_1
Xinput91 spi_dat_i[25] VGND VGND VPWR VPWR input91/X sky130_fd_sc_hd__clkbuf_2
Xinput80 spi_dat_i[15] VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1508__C _1508_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2166__B1 _2156_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2469__A1 _1768_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1677__C1 _1638_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2636__A _2638_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1540__A _1744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2355__B _2355_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2371__A _2371_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2920__CLK _2920_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2157__B1 _2156_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output141_A _1791_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2249__C _2265_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2546__A _2546_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1683__A2 _1682_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2265__B _2284_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2910_ _2915_/CLK _2910_/D VGND VGND VPWR VPWR _2910_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1435__A2 _2019_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2841_ _2901_/CLK _2841_/D VGND VGND VPWR VPWR _2841_/Q sky130_fd_sc_hd__dfxtp_1
X_2772_ _2776_/CLK _2772_/D VGND VGND VPWR VPWR _2772_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2281__A _2352_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1723_ _1723_/A VGND VGND VPWR VPWR _1723_/X sky130_fd_sc_hd__buf_4
XANTENNA__2396__B1 _2386_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1654_ _1652_/Y _1653_/Y _1606_/X VGND VGND VPWR VPWR _1654_/Y sky130_fd_sc_hd__a21oi_1
X_1585_ _2163_/A _2163_/B _1572_/X VGND VGND VPWR VPWR _1585_/Y sky130_fd_sc_hd__a21oi_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2206_ _1724_/Y _1725_/Y _2201_/X VGND VGND VPWR VPWR _2694_/D sky130_fd_sc_hd__a21oi_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1674__A2 _2189_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1360__A _1414_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2137_ input1/X VGND VGND VPWR VPWR _2537_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__2456__A _2558_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2175__B _2175_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2068_ _2838_/Q _2025_/X _2067_/X VGND VGND VPWR VPWR _2068_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_35_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1510__D _1510_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2943__CLK _2946_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2191__A _2191_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2387__B1 _1440_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1535__A _1699_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1665__A2 _1640_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2366__A _2366_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2378__B1 _2365_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output189_A _2075_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2393__A3 _2395_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1445__A _1445_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2040__S _2077_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1370_ _1370_/A _1409_/B VGND VGND VPWR VPWR _2377_/B sky130_fd_sc_hd__nand2_1
XANTENNA__2550__B1 _1865_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2816__CLK _2816_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2276__A _2324_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2267__C_N _2257_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1656__A2 _1609_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1330__D _1367_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1408__A2 _1380_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1931__A1_N _2887_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2824_ _2847_/CLK _2824_/D VGND VGND VPWR VPWR _2824_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1339__B _2382_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1577__D1 input96/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2755_ _2764_/CLK _2755_/D VGND VGND VPWR VPWR _2755_/Q sky130_fd_sc_hd__dfxtp_1
X_2686_ _2901_/CLK _2686_/D VGND VGND VPWR VPWR _2686_/Q sky130_fd_sc_hd__dfxtp_1
X_1706_ _1697_/X _1703_/Y _1704_/X _1705_/X VGND VGND VPWR VPWR _1706_/X sky130_fd_sc_hd__o211a_1
X_1637_ _1709_/A VGND VGND VPWR VPWR _1637_/X sky130_fd_sc_hd__buf_2
XANTENNA__1355__A _1355_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1568_ _1568_/A VGND VGND VPWR VPWR _1712_/A sky130_fd_sc_hd__clkbuf_4
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2541__B1 _1832_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1499_ _1486_/Y _1487_/X _1491_/Y _1494_/Y _1498_/Y VGND VGND VPWR VPWR _1512_/A
+ sky130_fd_sc_hd__o2111a_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2186__A _2186_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1647__A2 _1612_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2633__B _2639_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1964__S _2013_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1583__A1 _1561_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2839__CLK _2839_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2532__B1 _1801_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2527__C _2653_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2031__A1_N _2902_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2540_ _2540_/A VGND VGND VPWR VPWR _2540_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2471_ _2447_/A _2448_/A _2470_/Y VGND VGND VPWR VPWR _2809_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__1574__A1 _1560_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1422_ _1422_/A _1454_/D _1454_/C VGND VGND VPWR VPWR _2366_/A sky130_fd_sc_hd__and3_2
XANTENNA__1326__A1 _1296_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1903__A _1911_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1353_ _1353_/A VGND VGND VPWR VPWR _1447_/C sky130_fd_sc_hd__clkbuf_2
X_1284_ _1304_/A _1372_/A _2881_/Q VGND VGND VPWR VPWR _1350_/A sky130_fd_sc_hd__a21oi_4
XFILLER_49_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1629__A2 _1612_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1341__C _1341_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2807_ _2809_/CLK _2807_/D VGND VGND VPWR VPWR _2807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2738_ _2834_/CLK _2738_/D VGND VGND VPWR VPWR _2738_/Q sky130_fd_sc_hd__dfxtp_1
X_2669_ _2946_/CLK _2669_/D VGND VGND VPWR VPWR _2669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1868__A2 _1853_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1813__A _2092_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2628__B _2628_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2644__A _2647_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input65_A cpu_dat_i[8] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1723__A _1723_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2538__B _2538_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1442__B _1442_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2554__A _2558_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2036__A2 _2033_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2704__D _2704_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1971_ _1971_/A _2008_/B _2267_/B VGND VGND VPWR VPWR _1971_/X sky130_fd_sc_hd__or3_1
XFILLER_14_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1547__A1 _1467_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2523_ _2523_/A _2525_/B VGND VGND VPWR VPWR _2845_/D sky130_fd_sc_hd__nand2_1
XFILLER_6_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2454_ _2453_/X _2204_/A _1716_/X VGND VGND VPWR VPWR _2454_/Y sky130_fd_sc_hd__a21oi_1
X_2385_ _2385_/A VGND VGND VPWR VPWR _2767_/D sky130_fd_sc_hd__clkbuf_1
X_1405_ _1379_/X _1488_/A _2877_/Q VGND VGND VPWR VPWR _1509_/A sky130_fd_sc_hd__o21ai_1
XFILLER_60_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1336_ _2880_/Q _1324_/X _1335_/Y VGND VGND VPWR VPWR _1341_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__1633__A _1633_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput1 RST_N VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__buf_2
XFILLER_64_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1483__B1 _1482_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2578__A3 _2399_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2432__C1 _2431_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2684__CLK _2901_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1808__A _2113_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1538__A1 input73/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1527__B _1527_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2639__A _2639_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2499__C1 _2488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1543__A _1543_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2374__A _2374_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1777__A1 _1773_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2423__C1 _2405_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output171_A _1852_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2549__A _2549_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2170_ _1604_/Y _1605_/Y _2156_/X VGND VGND VPWR VPWR _2678_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__1701__A1 _1672_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1900__B _2945_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2284__A _2284_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2009__A2 _1969_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1954_ _2065_/A VGND VGND VPWR VPWR _2008_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1768__A1 _1558_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1885_ _1889_/A _2938_/Q VGND VGND VPWR VPWR _1886_/A sky130_fd_sc_hd__and2_1
X_2506_ _2540_/A VGND VGND VPWR VPWR _2506_/X sky130_fd_sc_hd__clkbuf_2
X_2437_ _1650_/X _1654_/Y _2436_/X _2431_/X VGND VGND VPWR VPWR _2790_/D sky130_fd_sc_hd__o211a_1
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2368_ _2368_/A _2368_/B VGND VGND VPWR VPWR _2370_/A sky130_fd_sc_hd__nand2_1
XANTENNA__2496__A2 _2493_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2299_ _2299_/A VGND VGND VPWR VPWR _2731_/D sky130_fd_sc_hd__clkbuf_1
X_1319_ _2756_/Q _1409_/B _1318_/Y VGND VGND VPWR VPWR _1319_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2194__A _2194_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1456__B1 _1455_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1759__A1 _1723_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2641__B _2932_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2420__A2 _1591_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2133__S _2243_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2184__A1 _1652_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1931__B2 _2487_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1392__C1 _1431_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput190 _2081_/Y VGND VGND VPWR VPWR spi_dat_o[24] sky130_fd_sc_hd__buf_2
XFILLER_43_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2369__A _2526_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2088__B _2109_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input28_A cpu_adr_i[4] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1423__D _1508_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1695__B1 _1667_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1998__B2 _2500_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2411__A2 _1913_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2270__C _2289_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1670_ _1624_/X _1609_/X _2793_/Q VGND VGND VPWR VPWR _1670_/X sky130_fd_sc_hd__o21a_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2279__A _2279_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _1769_/Y _1770_/Y _2172_/B VGND VGND VPWR VPWR _2702_/D sky130_fd_sc_hd__a21oi_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2153_ _2153_/A VGND VGND VPWR VPWR _2671_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1686__B1 _2689_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1911__A _1911_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_6_CLK_A clkbuf_1_0_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2084_ _2841_/Q _2033_/X _2083_/X VGND VGND VPWR VPWR _2518_/A sky130_fd_sc_hd__o21ai_1
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1989__A1 input36/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1438__B1 _1436_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1358__A _1362_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1937_ _2364_/A _1990_/B _2254_/A VGND VGND VPWR VPWR _1937_/X sky130_fd_sc_hd__or3_1
X_1868_ _1859_/X _1853_/X _2639_/A VGND VGND VPWR VPWR _1868_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__1610__B1 _2785_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput81 spi_dat_i[16] VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput70 cpu_sel_i[3] VGND VGND VPWR VPWR input70/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1508__D _1508_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput92 spi_dat_i[26] VGND VGND VPWR VPWR input92/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2166__A1 _1589_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1799_ _2027_/A VGND VGND VPWR VPWR _1970_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__2722__CLK _2745_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2189__A _2189_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2872__CLK _2880_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2469__A2 _1771_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1677__B1 _1637_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2636__B _2636_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2355__C _2370_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2652__A _2652_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2802__D _2802_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1601__B1 _1572_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2157__A1 _1537_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2099__A _2109_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output134_A _1586_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2265__C _2265_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2093__A0 _2738_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2840_ _2840_/CLK _2840_/D VGND VGND VPWR VPWR _2840_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2562__A _2573_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2396__A1 _2773_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2771_ _2880_/CLK _2771_/D VGND VGND VPWR VPWR _2771_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2745__CLK _2745_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2712__D _2712_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1722_ _1707_/X _1689_/X _2800_/Q VGND VGND VPWR VPWR _1722_/X sky130_fd_sc_hd__o21a_1
X_1653_ _1620_/X _1640_/X _2684_/Q VGND VGND VPWR VPWR _1653_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__1906__A _1906_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2895__CLK _2917_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1584_ _1567_/X _1569_/X _2675_/Q VGND VGND VPWR VPWR _2163_/B sky130_fd_sc_hd__o21ai_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1659__B1 _2685_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2205_ _2205_/A VGND VGND VPWR VPWR _2693_/D sky130_fd_sc_hd__clkbuf_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2136_ _2649_/A VGND VGND VPWR VPWR _2136_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1360__B _1414_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2067_ _2078_/A _2109_/B _2303_/A VGND VGND VPWR VPWR _2067_/X sky130_fd_sc_hd__or3_1
XANTENNA__2084__B1 _2083_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1787__S _2374_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1831__A0 _2749_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2387__A1 _2769_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1816__A _2114_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2121__A2_N _1530_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2647__A _2647_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1551__A _2949_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2366__B _2366_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2768__CLK _2768_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2382__A _2382_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1822__B1 _1804_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input95_A spi_dat_i[29] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2378__A1 _1362_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1586__C1 _1556_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2550__A1 _2860_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1461__A _1461_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2557__A _2557_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2707__D _2707_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2066__A0 _2733_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2292__A _2292_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2823_ _2901_/CLK _2823_/D VGND VGND VPWR VPWR _2823_/Q sky130_fd_sc_hd__dfxtp_1
X_2754_ _2929_/CLK _2754_/D VGND VGND VPWR VPWR _2754_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1339__C _1343_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1577__C1 _1536_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1705_ _1740_/A VGND VGND VPWR VPWR _1705_/X sky130_fd_sc_hd__clkbuf_2
X_2685_ _2839_/CLK _2685_/D VGND VGND VPWR VPWR _2685_/Q sky130_fd_sc_hd__dfxtp_1
X_1636_ _1635_/X _1617_/X _2788_/Q VGND VGND VPWR VPWR _1636_/X sky130_fd_sc_hd__o21a_1
X_1567_ _1744_/A VGND VGND VPWR VPWR _1567_/X sky130_fd_sc_hd__buf_4
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2541__A1 _2854_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ _1495_/Y _1497_/Y _1408_/Y _1411_/Y VGND VGND VPWR VPWR _1498_/Y sky130_fd_sc_hd__a22oi_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1371__A _1371_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2186__B _2194_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1501__C1 _1479_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2119_ _2128_/A _2128_/B _2238_/A VGND VGND VPWR VPWR _2119_/X sky130_fd_sc_hd__or3_1
XFILLER_55_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2910__CLK _2915_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1583__A2 _1582_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2532__A1 _2850_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2377__A _2382_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input10_A cpu_adr_i[17] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2048__A0 _2730_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2470_ _2453_/A _2224_/A _1773_/X VGND VGND VPWR VPWR _2470_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__1574__A2 _1573_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1421_ _1447_/C VGND VGND VPWR VPWR _1454_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1326__A2 _1297_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1352_ _2878_/Q _1343_/X _1351_/Y VGND VGND VPWR VPWR _1508_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__1903__B _2946_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2933__CLK _2946_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1283_ _2777_/Q _1289_/A _1291_/A VGND VGND VPWR VPWR _1372_/A sky130_fd_sc_hd__nand3b_4
XANTENNA__2287__A _2287_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1341__D _1341_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2806_ _2809_/CLK _2806_/D VGND VGND VPWR VPWR _2806_/Q sky130_fd_sc_hd__dfxtp_1
X_2737_ _2745_/CLK _2737_/D VGND VGND VPWR VPWR _2737_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1366__A _1366_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2668_ _2670_/CLK _2668_/D VGND VGND VPWR VPWR _2668_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2900__D _2900_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1867__A2_N _1530_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1619_ _1576_/X _1588_/X _1533_/X _1536_/X _1619_/D1 VGND VGND VPWR VPWR _1619_/Y
+ sky130_fd_sc_hd__o2111ai_2
X_2599_ _2599_/A _2605_/B VGND VGND VPWR VPWR _2894_/D sky130_fd_sc_hd__nor2_1
XFILLER_59_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2197__A _2197_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input2_A cpu_adr_i[0] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1805__A2_N _1792_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2644__B _2934_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2106__A1_N _2915_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2450__B1 _2449_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2660__A _2660_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1992__A1_N _2896_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2202__B1 _2201_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2806__CLK _2809_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2810__D _2810_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input58_A cpu_dat_i[30] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1442__C _1510_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1492__A1 _1445_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1970_ _2718_/Q input64/X _1970_/S VGND VGND VPWR VPWR _2267_/B sky130_fd_sc_hd__mux2_1
XFILLER_42_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2441__B1 _1670_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1547__A2 _1545_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2720__D _2720_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2522_ _2844_/Q _2519_/X _2099_/X _2514_/X VGND VGND VPWR VPWR _2844_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1914__A _2233_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2453_ _2453_/A VGND VGND VPWR VPWR _2453_/X sky130_fd_sc_hd__clkbuf_2
X_2384_ _2384_/A _2391_/B _2399_/C VGND VGND VPWR VPWR _2385_/A sky130_fd_sc_hd__and3_1
X_1404_ _1379_/X _2401_/A _1403_/Y VGND VGND VPWR VPWR _1406_/B sky130_fd_sc_hd__o21a_1
XFILLER_60_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1335_ _2398_/A _2398_/B _1335_/C VGND VGND VPWR VPWR _1335_/Y sky130_fd_sc_hd__nand3_2
Xinput2 cpu_adr_i[0] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1483__A1 _1778_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2829__CLK _2901_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2432__B1 _2416_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2480__A _2529_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1538__A2 _1465_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1527__C _1527_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1824__A _1853_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2639__B _2639_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2499__B1 _1990_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2805__D _2805_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2423__B1 _2416_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1777__A2 _1776_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output164_A _1910_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1701__A2 _1685_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2284__B _2284_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2715__D _2715_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1953_ _2233_/A VGND VGND VPWR VPWR _1953_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2414__B1 _2413_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1909__A _1911_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1884_ _1884_/A VGND VGND VPWR VPWR _1884_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1768__A2 _1559_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_19_CLK clkbuf_1_0_0_CLK/X VGND VGND VPWR VPWR _2881_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1822__A1_N _2922_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2505_ _2505_/A _2508_/B VGND VGND VPWR VPWR _2831_/D sky130_fd_sc_hd__nand2_1
X_2436_ _2558_/A VGND VGND VPWR VPWR _2436_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2367_ _2758_/Q _1457_/X _2365_/Y _2366_/X VGND VGND VPWR VPWR _2758_/D sky130_fd_sc_hd__a211o_1
XFILLER_5_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2298_ _2298_/A _2308_/B _2313_/C VGND VGND VPWR VPWR _2299_/A sky130_fd_sc_hd__and3_1
X_1318_ input5/X _1367_/B _1353_/A _1414_/D VGND VGND VPWR VPWR _1318_/Y sky130_fd_sc_hd__nand4b_4
XFILLER_38_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2475__A _2493_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1456__A1 _1407_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2194__B _2194_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1759__A2 _2533_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2641__C _2653_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2184__A2 _1653_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1392__B1 _1391_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput191 _2086_/Y VGND VGND VPWR VPWR spi_dat_o[25] sky130_fd_sc_hd__buf_2
Xoutput180 _2024_/Y VGND VGND VPWR VPWR spi_dat_o[15] sky130_fd_sc_hd__buf_2
XFILLER_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2088__C _2313_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1695__A1 _1690_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2385__A _2385_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1729__A _1735_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1604__D1 _1604_/D1 VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_opt_3_0_CLK clkbuf_1_1_0_CLK/X VGND VGND VPWR VPWR clkbuf_opt_3_0_CLK/X sky130_fd_sc_hd__clkbuf_16
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2221_ _2221_/A VGND VGND VPWR VPWR _2701_/D sky130_fd_sc_hd__clkbuf_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2279__B _2284_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_8_CLK clkbuf_1_1_0_CLK/X VGND VGND VPWR VPWR _2917_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2674__CLK _2920_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2152_ _2949_/A _2152_/B _2401_/B VGND VGND VPWR VPWR _2153_/A sky130_fd_sc_hd__and3_1
XANTENNA__1686__A1 _1672_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1911__B _2670_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2295__A _2295_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2083_ _2094_/A _2114_/B _2310_/B VGND VGND VPWR VPWR _2083_/X sky130_fd_sc_hd__or3_1
XFILLER_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1438__A1 _2765_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1936_ _2713_/Q input57/X _2132_/S VGND VGND VPWR VPWR _2254_/A sky130_fd_sc_hd__mux2_1
XANTENNA__1358__B _2368_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1867_ _2930_/Q _1530_/X _1840_/X _1866_/Y VGND VGND VPWR VPWR _2639_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__1610__A1 _1558_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput82 spi_dat_i[17] VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__clkbuf_2
Xinput60 cpu_dat_i[3] VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__clkbuf_1
Xinput71 cpu_stb_i VGND VGND VPWR VPWR _1289_/A sky130_fd_sc_hd__buf_2
X_1798_ _2047_/A VGND VGND VPWR VPWR _2027_/A sky130_fd_sc_hd__buf_2
Xinput93 spi_dat_i[27] VGND VGND VPWR VPWR input93/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2166__A2 _1590_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1374__A _2377_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2189__B _2189_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2419_ _2408_/X _2410_/X _2418_/Y VGND VGND VPWR VPWR _2781_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__1677__A1 _1651_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1549__A _1702_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1601__A1 _2167_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2157__A2 _1544_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2697__CLK _2703_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input40_A cpu_dat_i[14] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2099__B _2109_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output127_A _1752_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2093__A1 input54/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2562__B _2562_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2770_ _2776_/CLK _2770_/D VGND VGND VPWR VPWR _2770_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2396__A2 _1785_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1721_ _1716_/X _1720_/Y _1704_/X _1705_/X VGND VGND VPWR VPWR _1721_/X sky130_fd_sc_hd__o211a_1
X_1652_ _1651_/X _1588_/X _1637_/X _1638_/X input77/X VGND VGND VPWR VPWR _1652_/Y
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_7_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1583_ _1561_/X _1582_/X _1564_/X _1565_/X input99/X VGND VGND VPWR VPWR _2163_/A
+ sky130_fd_sc_hd__o2111ai_2
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1659__A1 _1599_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2204_ _2204_/A _2216_/B VGND VGND VPWR VPWR _2205_/A sky130_fd_sc_hd__or2_1
XANTENNA__1922__A _2364_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2135_ _1859_/A _2649_/A _2587_/B VGND VGND VPWR VPWR _2135_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2066_ _2733_/Q input49/X _2077_/S VGND VGND VPWR VPWR _2303_/A sky130_fd_sc_hd__mux2_1
XANTENNA__1360__C _1360_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2084__A1 _2841_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1831__A1 input29/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2903__D _2903_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2387__A2 _1785_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1919_ _2019_/A VGND VGND VPWR VPWR _2358_/A sky130_fd_sc_hd__clkbuf_4
X_2899_ _2901_/CLK _2899_/D VGND VGND VPWR VPWR _2899_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2544__C1 _2531_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1347__B1 _1346_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1832__A _2109_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2647__B _2936_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1551__B _1698_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2366__C input7/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2663__A _2663_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1822__B2 _1821_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2813__D _2813_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2382__B _2382_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input88_A spi_dat_i[22] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2378__A2 _1362_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1586__B1 _1473_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_5_CLK_A clkbuf_1_0_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1338__B1 _2766_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2550__A2 _2540_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1461__B _1511_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2066__A1 input49/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2712__CLK _2745_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2573__A _2573_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2723__D _2723_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2822_ _2847_/CLK _2822_/D VGND VGND VPWR VPWR _2822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2753_ _2764_/CLK _2753_/D VGND VGND VPWR VPWR _2753_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2862__CLK _2873_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1577__B1 _1533_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1917__A _2033_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1704_ _1739_/A VGND VGND VPWR VPWR _1704_/X sky130_fd_sc_hd__clkbuf_2
X_2684_ _2901_/CLK _2684_/D VGND VGND VPWR VPWR _2684_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1329__B1 _2770_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1635_ _1707_/A VGND VGND VPWR VPWR _1635_/X sky130_fd_sc_hd__clkbuf_2
X_1566_ _1561_/X _2064_/A _1564_/X _1565_/X input85/X VGND VGND VPWR VPWR _2158_/A
+ sky130_fd_sc_hd__o2111ai_2
XFILLER_59_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2541__A2 _2540_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1497_ _1367_/A _1457_/A _1496_/Y _1287_/X VGND VGND VPWR VPWR _1497_/Y sky130_fd_sc_hd__o211ai_2
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1501__B1 _1329_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2118_ _2707_/Q input67/X _2127_/S VGND VGND VPWR VPWR _2238_/A sky130_fd_sc_hd__mux2_1
XANTENNA__2483__A _2529_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2049_ _2094_/A _2072_/B _2296_/B VGND VGND VPWR VPWR _2049_/X sky130_fd_sc_hd__or3_1
XFILLER_54_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2517__C1 _2514_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2532__A2 _2519_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1562__A _1562_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2377__B _2377_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2735__CLK _2834_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2808__D _2808_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2048__A1 input45/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2885__CLK _2925_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output194_A _2102_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1420_ _1447_/D VGND VGND VPWR VPWR _1454_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_1351_ _1348_/Y _1306_/A _1349_/Y _1362_/A VGND VGND VPWR VPWR _1351_/Y sky130_fd_sc_hd__o211ai_4
XANTENNA__1731__B1 _2695_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1472__A _2451_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2529__C_N _2352_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1282_ _2776_/Q VGND VGND VPWR VPWR _1304_/A sky130_fd_sc_hd__inv_2
XFILLER_49_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2718__D _2718_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2805_ _2809_/CLK _2805_/D VGND VGND VPWR VPWR _2805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2736_ _2834_/CLK _2736_/D VGND VGND VPWR VPWR _2736_/Q sky130_fd_sc_hd__dfxtp_1
X_2667_ _2946_/CLK _2667_/D VGND VGND VPWR VPWR _2667_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1970__A0 _2718_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1618_ _1517_/X _1617_/X _2786_/Q VGND VGND VPWR VPWR _1618_/X sky130_fd_sc_hd__o21a_1
X_2598_ _2598_/A _2604_/B VGND VGND VPWR VPWR _2893_/D sky130_fd_sc_hd__nand2_1
XFILLER_8_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1549_ _1702_/A VGND VGND VPWR VPWR _1549_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__2478__A _2510_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2758__CLK _2776_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1722__B1 _2800_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2197__B _2197_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2644__C _2653_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2450__A1 _2447_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2202__A1 _1711_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1713__B1 _2692_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1292__A _2777_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1442__D _1510_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output207_A _2126_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1492__A2 _1488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2441__A1 _2433_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1467__A _2705_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2521_ _2521_/A _2521_/B VGND VGND VPWR VPWR _2843_/D sky130_fd_sc_hd__nand2_1
XANTENNA__2900__CLK _2915_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2452_ _1708_/X _1714_/Y _2436_/X _2451_/X VGND VGND VPWR VPWR _2798_/D sky130_fd_sc_hd__o211a_1
X_1403_ _2671_/Q _2706_/Q VGND VGND VPWR VPWR _1403_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2298__A _2298_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2383_ _2383_/A _2383_/B VGND VGND VPWR VPWR _2384_/A sky130_fd_sc_hd__nand2_1
X_1334_ _1296_/X _1297_/X _2775_/Q VGND VGND VPWR VPWR _2398_/B sky130_fd_sc_hd__o21ai_1
Xinput3 cpu_adr_i[10] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1483__A2 _1807_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2432__A1 _1636_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2480__B _2480_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2074__A2_N _2018_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2911__D _2911_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2196__B1 _2179_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2719_ _2745_/CLK _2719_/D VGND VGND VPWR VPWR _2719_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1943__B1 _1942_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2499__A1 _2826_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2001__A _2065_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1840__A _2039_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2120__B1 _2119_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1459__C1 _1500_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input105_A spi_dat_i[9] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2423__A1 _1603_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1287__A _1335_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2821__D _2821_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2923__CLK _2925_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input70_A cpu_sel_i[3] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output157_A _1897_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2111__B1 _1804_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2284__C _2289_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1952_ _1980_/A _2593_/A VGND VGND VPWR VPWR _1952_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2581__A _2650_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2414__A1 _2408_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1883_ _1889_/A _2937_/Q VGND VGND VPWR VPWR _1884_/A sky130_fd_sc_hd__and2_1
XANTENNA__1909__B _2669_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2731__D _2731_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1925__A _1945_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2504_ _2830_/Q _2493_/X _2014_/X _2501_/X VGND VGND VPWR VPWR _2830_/D sky130_fd_sc_hd__o211a_1
X_2435_ _2427_/X _2428_/X _2434_/Y VGND VGND VPWR VPWR _2789_/D sky130_fd_sc_hd__o21ai_1
XFILLER_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2366_ _2366_/A _2366_/B input7/X VGND VGND VPWR VPWR _2366_/X sky130_fd_sc_hd__and3_1
X_1317_ _1354_/A VGND VGND VPWR VPWR _1414_/D sky130_fd_sc_hd__buf_2
X_2297_ _2297_/A VGND VGND VPWR VPWR _2730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2906__D _2906_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1456__A2 _1523_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2247__C_N _2227_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2946__CLK _2946_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1392__A1 _2758_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput170 _1848_/Y VGND VGND VPWR VPWR spi_adr_o[7] sky130_fd_sc_hd__buf_2
XANTENNA__1944__A1_N _2889_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput181 _2032_/Y VGND VGND VPWR VPWR spi_dat_o[16] sky130_fd_sc_hd__buf_2
Xoutput192 _2091_/Y VGND VGND VPWR VPWR spi_dat_o[26] sky130_fd_sc_hd__buf_2
XANTENNA__2666__A _2666_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1695__A2 _1694_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2816__D _2816_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1604__C1 _1536_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _2220_/A _2224_/B VGND VGND VPWR VPWR _2221_/A sky130_fd_sc_hd__or2_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2279__C _2289_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2819__CLK _2920_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2151_ _2151_/A VGND VGND VPWR VPWR _2670_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1686__A2 _1685_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2082_ _2736_/Q input52/X _2093_/S VGND VGND VPWR VPWR _2310_/B sky130_fd_sc_hd__mux2_1
XFILLER_19_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2726__D _2726_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1438__A2 _1477_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1935_ _2114_/B VGND VGND VPWR VPWR _1990_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1358__C _2368_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1866_ _2860_/Q _1841_/X _1865_/X VGND VGND VPWR VPWR _1866_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__1610__A2 _1609_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput72 cpu_we_i VGND VGND VPWR VPWR input72/X sky130_fd_sc_hd__clkbuf_4
Xinput50 cpu_dat_i[23] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_1
Xinput61 cpu_dat_i[4] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__clkbuf_1
X_1797_ _2065_/A VGND VGND VPWR VPWR _2128_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput94 spi_dat_i[28] VGND VGND VPWR VPWR input94/X sky130_fd_sc_hd__clkbuf_2
Xinput83 spi_dat_i[18] VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1374__B _2377_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2571__B1 _2495_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2418_ _2412_/X _2164_/A _1581_/X VGND VGND VPWR VPWR _2418_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__1677__A2 _1663_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2486__A _2510_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2349_ _2349_/A VGND VGND VPWR VPWR _2752_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1390__A _1390_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1598__D1 _1598_/D1 VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1601__A2 _2167_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1565__A _1699_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2099__C _2318_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input33_A cpu_adr_i[9] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2562__C_N _2415_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1589__D1 _1589_/D1 VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1720_ _2203_/A _2203_/B _1702_/X VGND VGND VPWR VPWR _1720_/Y sky130_fd_sc_hd__a21oi_1
X_1651_ _1723_/A VGND VGND VPWR VPWR _1651_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_8_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1475__A _1717_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1582_ _1735_/A VGND VGND VPWR VPWR _1582_/X sky130_fd_sc_hd__buf_4
XFILLER_4_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1659__A2 _1612_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2203_ _2203_/A _2203_/B VGND VGND VPWR VPWR _2204_/A sky130_fd_sc_hd__nand2_1
XANTENNA__1922__B _2358_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2134_ _1853_/A _2483_/B _1789_/A _2885_/Q VGND VGND VPWR VPWR _2587_/B sky130_fd_sc_hd__o22ai_2
XANTENNA__2791__CLK _2839_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1360__D _1367_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2065_ _2065_/A VGND VGND VPWR VPWR _2109_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2084__A2 _2033_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2898_ _2915_/CLK _2898_/D VGND VGND VPWR VPWR _2898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1918_ _2046_/A VGND VGND VPWR VPWR _2364_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1849_ _2752_/Q input32/X _1860_/S VGND VGND VPWR VPWR _2348_/B sky130_fd_sc_hd__mux2_1
XFILLER_8_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2544__B1 _1845_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1347__A1 _2866_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1832__B _1865_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2647__C _2653_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_opt_2_0_CLK clkbuf_1_0_0_CLK/X VGND VGND VPWR VPWR clkbuf_opt_2_1_CLK/A sky130_fd_sc_hd__clkbuf_16
XFILLER_14_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2382__C _2382_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2232__C1 _2577_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1586__A1 _1581_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1295__A _2776_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1338__A1 _1296_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1743__D1 input91/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1461__C _1461_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2573__B _2573_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2821_ _2920_/CLK _2821_/D VGND VGND VPWR VPWR _2821_/Q sky130_fd_sc_hd__dfxtp_1
X_2752_ _2873_/CLK _2752_/D VGND VGND VPWR VPWR _2752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1577__A1 _1576_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1703_ _2197_/A _2197_/B _1702_/X VGND VGND VPWR VPWR _1703_/Y sky130_fd_sc_hd__a21oi_1
X_2683_ _2901_/CLK _2683_/D VGND VGND VPWR VPWR _2683_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1329__A1 _1400_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1634_ _1625_/X _1631_/Y _1632_/X _1633_/X VGND VGND VPWR VPWR _1634_/X sky130_fd_sc_hd__o211a_1
X_1565_ _1699_/A VGND VGND VPWR VPWR _1565_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__1933__A _2064_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1496_ _2389_/A _1452_/X _2764_/Q VGND VGND VPWR VPWR _1496_/Y sky130_fd_sc_hd__o21ai_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1501__A1 _1330_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2117_ _2117_/A _2626_/A VGND VGND VPWR VPWR _2117_/Y sky130_fd_sc_hd__nor2_4
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2483__B _2483_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2048_ _2730_/Q input45/X _2093_/S VGND VGND VPWR VPWR _2296_/B sky130_fd_sc_hd__mux2_1
XANTENNA__2914__D _2914_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2687__CLK _2839_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2517__B1 _2078_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1843__A _2027_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2377__C _2377_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1989__S _2013_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2824__D _2824_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output187_A _2063_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1350_ _1350_/A VGND VGND VPWR VPWR _1362_/A sky130_fd_sc_hd__buf_4
XANTENNA__1731__A1 _1672_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2584__A _2618_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1495__B1 _1365_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2734__D _2734_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2804_ _2809_/CLK _2804_/D VGND VGND VPWR VPWR _2804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2735_ _2834_/CLK _2735_/D VGND VGND VPWR VPWR _2735_/Q sky130_fd_sc_hd__dfxtp_1
X_2666_ _2666_/A VGND VGND VPWR VPWR _2946_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1970__A1 input64/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1617_ _1689_/A VGND VGND VPWR VPWR _1617_/X sky130_fd_sc_hd__clkbuf_2
X_2597_ _2597_/A _2605_/B VGND VGND VPWR VPWR _2892_/D sky130_fd_sc_hd__nor2_1
XANTENNA__1663__A _1913_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1548_ _1548_/A VGND VGND VPWR VPWR _1702_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1722__A1 _1707_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2909__D _2909_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1479_ _1479_/A VGND VGND VPWR VPWR _2243_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_54_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_4_CLK_A clkbuf_1_0_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2450__A2 _2448_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2202__A2 _1713_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1410__B1 _2771_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2702__CLK _2816_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1713__A1 _1692_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1292__B _2776_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2819__D _2819_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2852__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2426__C1 _2405_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2441__A2 _2190_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2520_ _2842_/Q _2519_/X _2088_/X _2514_/X VGND VGND VPWR VPWR _2842_/D sky130_fd_sc_hd__o211a_1
X_2451_ _2451_/A VGND VGND VPWR VPWR _2451_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1402_ _2395_/A _2395_/D _1422_/A VGND VGND VPWR VPWR _2401_/A sky130_fd_sc_hd__o21ai_2
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2298__B _2308_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2382_ _2382_/A _2382_/B _2382_/C _2382_/D VGND VGND VPWR VPWR _2766_/D sky130_fd_sc_hd__nand4_1
XFILLER_57_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1333_ _1333_/A _1390_/A VGND VGND VPWR VPWR _2398_/A sky130_fd_sc_hd__nand2_4
XANTENNA__2729__D _2729_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1468__B1 _1467_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput4 cpu_adr_i[11] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2417__C1 _2405_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2432__A2 _1642_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2196__A1 _1691_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2725__CLK _2745_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2718_ _2745_/CLK _2718_/D VGND VGND VPWR VPWR _2718_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1943__A1 _2819_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2649_ _2649_/A VGND VGND VPWR VPWR _2649_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2875__CLK _2881_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2499__A2 _2493_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_opt_1_0_CLK_A clkbuf_1_0_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2120__A1 _2812_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1459__B1 _1458_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1568__A _1568_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2423__A2 _1607_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1631__B1 _1630_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input63_A cpu_dat_i[6] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2399__A _2399_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2111__B2 _2110_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1951_ _2890_/Q _1933_/X _1916_/X _1950_/Y VGND VGND VPWR VPWR _2593_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__2414__A2 _2410_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2748__CLK _2873_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1882_ _1882_/A VGND VGND VPWR VPWR _1882_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1622__B1 _1606_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1925__B _2588_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2898__CLK _2915_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2503_ _2503_/A _2508_/B VGND VGND VPWR VPWR _2829_/D sky130_fd_sc_hd__nand2_1
XFILLER_6_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2102__A _2102_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2434_ _2433_/X _2182_/A _1644_/X VGND VGND VPWR VPWR _2434_/Y sky130_fd_sc_hd__a21oi_1
X_2365_ _2401_/C _2358_/A _2227_/A VGND VGND VPWR VPWR _2365_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_5_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1316_ _1390_/A VGND VGND VPWR VPWR _1409_/B sky130_fd_sc_hd__buf_2
X_2296_ _2296_/A _2296_/B _2281_/X VGND VGND VPWR VPWR _2297_/A sky130_fd_sc_hd__or3b_1
XANTENNA__1973__A2_N _1953_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1861__A0 _2353_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2922__D _2922_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1388__A _1388_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1613__B1 _2679_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput160 _1904_/X VGND VGND VPWR VPWR spi_adr_o[27] sky130_fd_sc_hd__buf_2
XANTENNA__2012__A _2076_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1392__A2 _1428_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput182 _2038_/Y VGND VGND VPWR VPWR spi_dat_o[17] sky130_fd_sc_hd__buf_2
Xoutput193 _2097_/Y VGND VGND VPWR VPWR spi_dat_o[27] sky130_fd_sc_hd__buf_2
Xoutput171 _1852_/Y VGND VGND VPWR VPWR spi_adr_o[8] sky130_fd_sc_hd__buf_2
XFILLER_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1852__B1 _2636_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1604__B1 _1533_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2832__D _2832_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1368__C1 _1335_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2150_ _2647_/A _2670_/Q _2401_/B VGND VGND VPWR VPWR _2151_/A sky130_fd_sc_hd__and3_1
X_2081_ _2102_/A _2617_/A VGND VGND VPWR VPWR _2081_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2096__B1 _2058_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2592__A _2592_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2742__D _2742_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1934_ _2019_/A VGND VGND VPWR VPWR _2114_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput40 cpu_dat_i[14] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_1
X_1865_ _2128_/A _1865_/B _2355_/A VGND VGND VPWR VPWR _1865_/X sky130_fd_sc_hd__or3_1
Xinput73 spi_ack_i VGND VGND VPWR VPWR input73/X sky130_fd_sc_hd__clkbuf_4
Xinput51 cpu_dat_i[24] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_1
Xinput62 cpu_dat_i[5] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__clkbuf_1
X_1796_ _2019_/A VGND VGND VPWR VPWR _2065_/A sky130_fd_sc_hd__buf_2
Xinput95 spi_dat_i[29] VGND VGND VPWR VPWR input95/X sky130_fd_sc_hd__clkbuf_2
Xinput84 spi_dat_i[19] VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2020__A0 _2726_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1374__C _1437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2571__A1 _1500_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2417_ _1575_/X _1579_/Y _2416_/X _2405_/X VGND VGND VPWR VPWR _2780_/D sky130_fd_sc_hd__o211a_1
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2348_ _2353_/A _2348_/B _2329_/X VGND VGND VPWR VPWR _2349_/A sky130_fd_sc_hd__or3b_1
XFILLER_45_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2917__D _2917_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2279_ _2279_/A _2284_/B _2289_/C VGND VGND VPWR VPWR _2280_/A sky130_fd_sc_hd__and3_1
XANTENNA__2913__CLK _2915_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2087__A0 _2737_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1834__B1 _1804_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1598__C1 _1565_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2827__D _2827_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input26_A cpu_adr_i[31] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1825__A0 _2748_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1589__C1 _1536_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1650_ _1635_/X _1617_/X _2790_/Q VGND VGND VPWR VPWR _1650_/X sky130_fd_sc_hd__o21a_1
X_1581_ _1558_/X _1559_/X _2781_/Q VGND VGND VPWR VPWR _1581_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2002__A0 _2723_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2936__CLK _2946_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2587__A _2632_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2202_ _1711_/Y _1713_/Y _2201_/X VGND VGND VPWR VPWR _2692_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__1922__C _2249_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1398__A_N input22/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2737__D _2737_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2133_ _2247_/B _2815_/Q _2243_/A VGND VGND VPWR VPWR _2483_/B sky130_fd_sc_hd__mux2_1
XANTENNA__2069__B1 _2039_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2064_ _2064_/A VGND VGND VPWR VPWR _2064_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2897_ _2901_/CLK _2897_/D VGND VGND VPWR VPWR _2897_/Q sky130_fd_sc_hd__dfxtp_1
X_1917_ _2033_/A VGND VGND VPWR VPWR _2353_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1958__A1_N _2891_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1848_ _1830_/X _1824_/X _2635_/A VGND VGND VPWR VPWR _1848_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1779_ _1859_/A VGND VGND VPWR VPWR _1779_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2544__A1 _2856_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1347__A2 _1343_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1752__C1 _1740_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2497__A _2510_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1832__C _2342_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2382__D _2382_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1576__A _1723_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2232__B1 _1545_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2809__CLK _2809_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1586__A2 _1585_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2090__A1_N _2912_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1338__A2 _1372_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1743__C1 _1699_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2200__A _2200_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output132_A _1772_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2043__A1_N _2904_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2471__B1 _2470_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2820_ _2847_/CLK _2820_/D VGND VGND VPWR VPWR _2820_/Q sky130_fd_sc_hd__dfxtp_1
X_2751_ _2764_/CLK _2751_/D VGND VGND VPWR VPWR _2751_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1577__A2 _1530_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2682_ _2901_/CLK _2682_/D VGND VGND VPWR VPWR _2682_/Q sky130_fd_sc_hd__dfxtp_1
X_1702_ _1702_/A VGND VGND VPWR VPWR _1702_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1486__A _2870_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1633_ _1633_/A VGND VGND VPWR VPWR _1633_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1329__A2 _1371_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1564_ _1698_/A VGND VGND VPWR VPWR _1564_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_59_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1495_ _1445_/X _1426_/X _1365_/Y VGND VGND VPWR VPWR _1495_/Y sky130_fd_sc_hd__o21ai_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1501__A2 _1477_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2116_ _2917_/Q _1914_/X _1916_/X _2525_/A VGND VGND VPWR VPWR _2626_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2047_ _2047_/A VGND VGND VPWR VPWR _2093_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2462__B1 _2461_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2949_ _2949_/A VGND VGND VPWR VPWR _2949_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2214__B1 _2201_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2930__D _2930_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1396__A _2372_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2517__A1 _2840_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2377__D _2382_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1538__B1_N _2705_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input93_A spi_dat_i[27] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2781__CLK _2816_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2840__D _2840_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1731__A2 _1685_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1495__A1 _1445_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2444__B1 _1683_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1652__D1 input77/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2803_ _2809_/CLK _2803_/D VGND VGND VPWR VPWR _2803_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2750__D _2750_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2734_ _2834_/CLK _2734_/D VGND VGND VPWR VPWR _2734_/Q sky130_fd_sc_hd__dfxtp_1
X_2665_ _2665_/A _2946_/Q _2665_/C VGND VGND VPWR VPWR _2666_/A sky130_fd_sc_hd__and3_1
X_2596_ _2650_/A VGND VGND VPWR VPWR _2605_/B sky130_fd_sc_hd__clkbuf_2
X_1616_ _1616_/A VGND VGND VPWR VPWR _1689_/A sky130_fd_sc_hd__clkbuf_4
Xclkbuf_opt_1_0_CLK clkbuf_1_0_0_CLK/X VGND VGND VPWR VPWR clkbuf_leaf_0_CLK/A sky130_fd_sc_hd__clkbuf_16
X_1547_ _1467_/X _1545_/Y _1546_/Y VGND VGND VPWR VPWR _1548_/A sky130_fd_sc_hd__o21ai_2
XFILLER_8_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1722__A2 _1689_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1478_ _2743_/Q input72/X _2047_/A VGND VGND VPWR VPWR _2327_/A sky130_fd_sc_hd__mux2_2
XFILLER_28_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2925__D _2925_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2435__B1 _2434_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1410__A1 _1451_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1713__A2 _1712_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2835__D _2835_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2426__B1 _2416_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2450_ _2447_/X _2448_/X _2449_/Y VGND VGND VPWR VPWR _2797_/D sky130_fd_sc_hd__o21ai_1
XFILLER_5_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1401_ _1401_/A VGND VGND VPWR VPWR _2395_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__2298__C _2313_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2381_ _2381_/A VGND VGND VPWR VPWR _2765_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2677__CLK _2816_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1332_ _1329_/X _1479_/A _1330_/X _1331_/Y VGND VGND VPWR VPWR _1341_/B sky130_fd_sc_hd__o31ai_4
XANTENNA__2595__A _2595_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1468__A1 _2949_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput5 cpu_adr_i[12] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2745__D _2745_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2417__B1 _2416_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2196__A2 _1693_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2717_ _2745_/CLK _2717_/D VGND VGND VPWR VPWR _2717_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1943__A2 _2474_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2648_ _2648_/A VGND VGND VPWR VPWR _2936_/D sky130_fd_sc_hd__clkbuf_1
X_2579_ _2357_/X _2401_/A _2554_/X _2527_/A VGND VGND VPWR VPWR _2881_/D sky130_fd_sc_hd__o211a_1
XFILLER_19_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1459__A1 _1414_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2120__A2 _1841_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1631__A1 _2175_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1395__B1 _2760_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2399__B _2401_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input56_A cpu_dat_i[29] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1950_ _2820_/Q _2353_/A _1949_/X VGND VGND VPWR VPWR _1950_/Y sky130_fd_sc_hd__o21ai_1
X_1881_ _1889_/A _2936_/Q VGND VGND VPWR VPWR _1882_/A sky130_fd_sc_hd__and2_1
XANTENNA__1622__A1 _1619_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1386__B1 _1385_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2502_ _2828_/Q _2493_/X _2003_/X _2501_/X VGND VGND VPWR VPWR _2828_/D sky130_fd_sc_hd__o211a_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2102__B _2623_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_leaf_3_CLK_A clkbuf_1_0_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2433_ _2453_/A VGND VGND VPWR VPWR _2433_/X sky130_fd_sc_hd__clkbuf_2
X_2364_ _2364_/A VGND VGND VPWR VPWR _2401_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_29_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1315_ _1400_/A _1371_/A _1401_/A VGND VGND VPWR VPWR _1390_/A sky130_fd_sc_hd__nor3_4
XFILLER_57_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2295_ _2295_/A VGND VGND VPWR VPWR _2729_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1861__A1 _2859_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1388__B _1388_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1613__A1 _1599_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2842__CLK _2881_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1377__B1 _2765_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput161 _1906_/X VGND VGND VPWR VPWR spi_adr_o[28] sky130_fd_sc_hd__buf_2
Xoutput150 _1884_/X VGND VGND VPWR VPWR spi_adr_o[18] sky130_fd_sc_hd__buf_2
Xoutput194 _2102_/Y VGND VGND VPWR VPWR spi_dat_o[28] sky130_fd_sc_hd__buf_2
Xoutput183 _2044_/Y VGND VGND VPWR VPWR spi_dat_o[18] sky130_fd_sc_hd__buf_2
Xoutput172 _1858_/Y VGND VGND VPWR VPWR spi_adr_o[9] sky130_fd_sc_hd__buf_2
XFILLER_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1852__A1 _1830_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1604__A1 _1576_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1368__B1 _1367_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2203__A _2203_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output162_A _1908_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2080_ _2910_/Q _2064_/X _2039_/X _2079_/Y VGND VGND VPWR VPWR _2617_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2096__B2 _2521_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2715__CLK _2745_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2592__B _2638_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1933_ _2064_/A VGND VGND VPWR VPWR _1933_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2865__CLK _2873_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1864_ _2755_/Q input4/X _2127_/S VGND VGND VPWR VPWR _2355_/A sky130_fd_sc_hd__mux2_1
Xinput30 cpu_adr_i[6] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_1
Xinput52 cpu_dat_i[25] VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput41 cpu_dat_i[15] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_1
Xinput63 cpu_dat_i[6] VGND VGND VPWR VPWR input63/X sky130_fd_sc_hd__clkbuf_1
X_1795_ _2046_/A VGND VGND VPWR VPWR _1971_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1359__B1 _1358_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput96 spi_dat_i[2] VGND VGND VPWR VPWR input96/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput85 spi_dat_i[1] VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__clkbuf_2
Xinput74 spi_dat_i[0] VGND VGND VPWR VPWR input74/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2020__A1 input41/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2571__A2 _1501_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1952__A _1980_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2416_ _2558_/A VGND VGND VPWR VPWR _2416_/X sky130_fd_sc_hd__clkbuf_2
X_2347_ _2347_/A VGND VGND VPWR VPWR _2751_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2278_ _2278_/A VGND VGND VPWR VPWR _2722_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2087__A1 input53/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2933__D _2933_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1834__B2 _1833_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1598__B1 _1564_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2547__C1 _2531_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1770__B1 _2702_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2738__CLK _2834_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input19_A cpu_adr_i[25] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2888__CLK _2917_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2843__D _2843_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1825__A1 input28/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1589__B1 _1533_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2002__A1 input38/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1580_ _1575_/X _1579_/Y _1473_/X _1556_/X VGND VGND VPWR VPWR _1580_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1761__B1 _1630_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2587__B _2587_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1987__A2_N _1953_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2201_ _2224_/B VGND VGND VPWR VPWR _2201_/X sky130_fd_sc_hd__clkbuf_2
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2132_ _2710_/Q input70/X _2132_/S VGND VGND VPWR VPWR _2247_/B sky130_fd_sc_hd__mux2_1
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2063_ _2075_/A _2614_/A VGND VGND VPWR VPWR _2063_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2069__B2 _2068_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2753__D _2753_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1947__A _2117_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2896_ _2917_/CLK _2896_/D VGND VGND VPWR VPWR _2896_/Q sky130_fd_sc_hd__dfxtp_1
X_1916_ _2058_/A VGND VGND VPWR VPWR _1916_/X sky130_fd_sc_hd__clkbuf_2
X_1847_ _2926_/Q _1792_/X _1840_/X _1846_/Y VGND VGND VPWR VPWR _2635_/A sky130_fd_sc_hd__a2bb2o_1
X_1778_ _1778_/A VGND VGND VPWR VPWR _1859_/A sky130_fd_sc_hd__buf_2
XANTENNA__2544__A2 _2540_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1682__A _1682_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1752__B1 _1739_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2928__D _2928_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2018__A _2233_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2232__B2 _1467_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2232__A1 _2811_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1991__B1 _1990_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1743__B1 _1698_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1592__A _1739_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2838__D _2838_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2010__A2_N _1953_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output125_A _1741_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2471__A1 _2447_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2750_ _2873_/CLK _2750_/D VGND VGND VPWR VPWR _2750_/Q sky130_fd_sc_hd__dfxtp_1
X_1701_ _1672_/X _1685_/X _2691_/Q VGND VGND VPWR VPWR _2197_/B sky130_fd_sc_hd__o21ai_1
X_2681_ _2901_/CLK _2681_/D VGND VGND VPWR VPWR _2681_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1486__B _1523_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2903__CLK _2915_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1632_ _1632_/A VGND VGND VPWR VPWR _1632_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1329__A3 _1401_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2598__A _2598_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1563_ _1735_/A VGND VGND VPWR VPWR _2064_/A sky130_fd_sc_hd__buf_2
XANTENNA__1734__B1 _2802_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1494_ _1492_/Y _1346_/Y _1493_/Y _1339_/Y VGND VGND VPWR VPWR _1494_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2748__D _2748_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2115_ _2847_/Q _2251_/A _2114_/X VGND VGND VPWR VPWR _2525_/A sky130_fd_sc_hd__o21ai_2
X_2046_ _2046_/A VGND VGND VPWR VPWR _2094_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2462__A1 _2447_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2214__A1 _1749_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1396__B _2372_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1973__B1 _1927_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2879_ _2881_/CLK _2879_/D VGND VGND VPWR VPWR _2879_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__2517__A2 _2506_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1725__B1 _2694_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2301__A _2320_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1661__C1 _1633_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2926__CLK _2930_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input86_A spi_dat_i[20] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1964__A0 _2717_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1716__B1 _2799_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2211__A _2211_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2141__B1 _2140_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1495__A2 _1426_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2444__A1 _2433_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1652__C1 _1638_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2802_ _2809_/CLK _2802_/D VGND VGND VPWR VPWR _2802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2733_ _2834_/CLK _2733_/D VGND VGND VPWR VPWR _2733_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1955__A0 _2716_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2664_ _2945_/Q _2649_/X _2650_/X VGND VGND VPWR VPWR _2945_/D sky130_fd_sc_hd__a21o_1
XFILLER_8_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2595_ _2595_/A _2604_/B VGND VGND VPWR VPWR _2891_/D sky130_fd_sc_hd__nand2_1
X_1615_ _1610_/X _1614_/Y _1593_/X _1595_/X VGND VGND VPWR VPWR _1615_/X sky130_fd_sc_hd__o211a_1
X_1546_ _1463_/Y _2527_/A _2811_/Q VGND VGND VPWR VPWR _1546_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1477_ _1477_/A VGND VGND VPWR VPWR _2047_/A sky130_fd_sc_hd__buf_2
XANTENNA__1960__A _2092_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2132__A0 _2710_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2435__A1 _2427_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2029_ _2078_/A _2054_/B _2289_/A VGND VGND VPWR VPWR _2029_/X sky130_fd_sc_hd__or3_1
XFILLER_23_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1643__C1 _1633_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2941__D _2941_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1410__A2 _1452_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1870__A _1878_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2123__A0 _2708_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2426__A1 _1618_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1634__C1 _1633_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2851__D _2851_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output192_A _2091_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1400_ _1400_/A VGND VGND VPWR VPWR _2395_/A sky130_fd_sc_hd__buf_2
X_2380_ _2380_/A _2391_/B _2399_/C VGND VGND VPWR VPWR _2381_/A sky130_fd_sc_hd__and3_1
XANTENNA__1780__A _1807_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1331_ _1424_/A _1380_/A _2875_/Q VGND VGND VPWR VPWR _1331_/Y sky130_fd_sc_hd__o21bai_1
XANTENNA__2595__B _2604_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1468__A2 _1531_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput6 cpu_adr_i[13] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2087__S _2108_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2542__C_N _2537_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2417__A1 _1575_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2761__D _2761_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1834__A1_N _2924_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1928__A0 _2712_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2716_ _2745_/CLK _2716_/D VGND VGND VPWR VPWR _2716_/Q sky130_fd_sc_hd__dfxtp_1
X_2647_ _2647_/A _2936_/Q _2653_/C VGND VGND VPWR VPWR _2648_/A sky130_fd_sc_hd__and3_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2578_ _2401_/C _2358_/A _2399_/A _1490_/Y _2382_/D VGND VGND VPWR VPWR _2880_/D
+ sky130_fd_sc_hd__o311a_1
X_1529_ _1562_/A VGND VGND VPWR VPWR _1913_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__2936__D _2936_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2105__B1 _2104_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2771__CLK _2880_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1459__A2 _1457_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2671__D _2671_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2026__A _2114_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1631__A2 _2175_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1865__A _2128_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1395__A1 _1451_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2399__C _2399_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input49_A cpu_dat_i[22] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2846__D _2846_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output205_A _1988_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1880_ _1902_/A VGND VGND VPWR VPWR _1889_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1622__A2 _1621_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2583__B1 _2312_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1386__A1 _2874_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2501_ _2531_/A VGND VGND VPWR VPWR _2501_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2432_ _1636_/X _1642_/Y _2416_/X _2431_/X VGND VGND VPWR VPWR _2788_/D sky130_fd_sc_hd__o211a_1
X_2363_ _2757_/Q _1785_/S _1414_/Y _2386_/D _2382_/A VGND VGND VPWR VPWR _2757_/D
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__2794__CLK _2839_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1314_ _1353_/A _1354_/A VGND VGND VPWR VPWR _1401_/A sky130_fd_sc_hd__nand2_2
XFILLER_38_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2294_ _2294_/A _2308_/B _2313_/C VGND VGND VPWR VPWR _2295_/A sky130_fd_sc_hd__and3_1
XANTENNA__2756__D _2756_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1613__A2 _1612_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1685__A _1712_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1377__A1 _1307_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput151 _1886_/X VGND VGND VPWR VPWR spi_adr_o[19] sky130_fd_sc_hd__buf_2
Xoutput140 _1634_/X VGND VGND VPWR VPWR cpu_dat_o[9] sky130_fd_sc_hd__buf_2
Xoutput195 _2107_/Y VGND VGND VPWR VPWR spi_dat_o[29] sky130_fd_sc_hd__buf_2
Xoutput184 _2052_/Y VGND VGND VPWR VPWR spi_dat_o[19] sky130_fd_sc_hd__buf_2
Xoutput162 _1908_/X VGND VGND VPWR VPWR spi_adr_o[29] sky130_fd_sc_hd__buf_2
Xoutput173 _2949_/A VGND VGND VPWR VPWR spi_cyc_o sky130_fd_sc_hd__buf_2
XFILLER_0_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input103_A spi_dat_i[7] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1852__A2 _1824_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1604__A2 _1588_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2667__CLK _2946_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1595__A _1633_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1368__A1 _2764_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2565__B1 _2552_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2203__B _2203_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output155_A _1893_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1932_ _1945_/A _2590_/A VGND VGND VPWR VPWR _1932_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1863_ _1859_/X _1853_/X _2638_/B VGND VGND VPWR VPWR _1863_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_30_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput31 cpu_adr_i[7] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_1
Xinput20 cpu_adr_i[26] VGND VGND VPWR VPWR _1330_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_0_CLK_A CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput53 cpu_dat_i[26] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__buf_2
Xinput42 cpu_dat_i[16] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_1
Xinput64 cpu_dat_i[7] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1359__A1 _2864_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1794_ _1815_/A VGND VGND VPWR VPWR _2046_/A sky130_fd_sc_hd__clkbuf_2
Xinput97 spi_dat_i[30] VGND VGND VPWR VPWR input97/X sky130_fd_sc_hd__buf_4
Xinput86 spi_dat_i[20] VGND VGND VPWR VPWR input86/X sky130_fd_sc_hd__clkbuf_2
Xinput75 spi_dat_i[10] VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1764__D1 input95/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1952__B _2593_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2415_ _2415_/A VGND VGND VPWR VPWR _2558_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1525__A2_N _1327_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2346_ _2346_/A _2355_/B _2370_/C VGND VGND VPWR VPWR _2347_/A sky130_fd_sc_hd__and3_1
X_2277_ _2296_/A _2277_/B _2257_/X VGND VGND VPWR VPWR _2278_/A sky130_fd_sc_hd__or3b_1
XFILLER_38_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1598__A1 _1561_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2547__B1 _1855_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2304__A _2304_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1770__A1 _1567_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_2_CLK_A clkbuf_1_0_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1589__A1 _1576_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1761__A1 _1759_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _2200_/A VGND VGND VPWR VPWR _2691_/D sky130_fd_sc_hd__clkbuf_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2131_ _1859_/X _2649_/A _2586_/A VGND VGND VPWR VPWR _2131_/Y sky130_fd_sc_hd__a21oi_2
X_2062_ _2907_/Q _2018_/X _2058_/X _2513_/A VGND VGND VPWR VPWR _2614_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__2832__CLK _2834_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1915_ _2039_/A VGND VGND VPWR VPWR _2058_/A sky130_fd_sc_hd__buf_2
X_2895_ _2917_/CLK _2895_/D VGND VGND VPWR VPWR _2895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1846_ _2856_/Q _1841_/X _1845_/X VGND VGND VPWR VPWR _1846_/Y sky130_fd_sc_hd__o21ai_1
X_1777_ _1773_/X _1776_/Y _1632_/A _1633_/A VGND VGND VPWR VPWR _1777_/X sky130_fd_sc_hd__o211a_2
XANTENNA__1963__A _2027_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1752__A1 _1748_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1504__A1 _1445_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2329_ _2352_/A VGND VGND VPWR VPWR _2329_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_58_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2944__D _2944_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2232__A2 _1464_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1991__A1 _2826_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1873__A _1873_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2705__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1743__A1 _1717_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2855__CLK _2925_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input31_A cpu_adr_i[7] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2854__D _2854_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2209__A _2209_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output118_A _1695_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2471__A2 _2448_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1700_ _1645_/X _1657_/X _1698_/X _1699_/X input84/X VGND VGND VPWR VPWR _2197_/A
+ sky130_fd_sc_hd__o2111ai_4
X_2680_ _2901_/CLK _2680_/D VGND VGND VPWR VPWR _2680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1631_ _2175_/A _2175_/B _1630_/X VGND VGND VPWR VPWR _1631_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1783__A _2047_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2598__B _2604_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1562_ _1562_/A VGND VGND VPWR VPWR _1735_/A sky130_fd_sc_hd__buf_4
XANTENNA__1734__A1 _1707_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1493_ _1445_/X _1488_/X _2871_/Q VGND VGND VPWR VPWR _1493_/Y sky130_fd_sc_hd__o21bai_2
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1498__B1 _1408_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2114_ _2114_/A _2114_/B _2325_/B VGND VGND VPWR VPWR _2114_/X sky130_fd_sc_hd__or3_1
XFILLER_55_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2764__D _2764_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2045_ _2076_/A VGND VGND VPWR VPWR _2075_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2119__A _2128_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2462__A2 _2448_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1670__B1 _2793_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2214__A2 _1750_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2728__CLK _2834_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1396__C _1437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1973__B2 _2495_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2878_ _2881_/CLK _2878_/D VGND VGND VPWR VPWR _2878_/Q sky130_fd_sc_hd__dfxtp_1
X_1829_ _1779_/X _1824_/X _2632_/B VGND VGND VPWR VPWR _1829_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__1725__A1 _1692_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2878__CLK _2881_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2939__D _2939_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2301__B _2301_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2674__D _2674_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2029__A _2078_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1661__B1 _1632_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1964__A1 input63/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input79_A spi_dat_i[14] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1716__A1 _1696_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2211__B _2211_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2849__D _2849_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1924__A2_N _1914_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2141__A1 _2667_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1939__A2_N _1933_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1778__A _1778_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2444__A2 _2194_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1652__B1 _1637_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2801_ _2809_/CLK _2801_/D VGND VGND VPWR VPWR _2801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2732_ _2834_/CLK _2732_/D VGND VGND VPWR VPWR _2732_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1404__B1 _1403_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1955__A1 input62/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2663_ _2663_/A VGND VGND VPWR VPWR _2944_/D sky130_fd_sc_hd__clkbuf_1
X_2594_ _2618_/A VGND VGND VPWR VPWR _2604_/B sky130_fd_sc_hd__clkbuf_2
X_1614_ _2171_/A _2171_/B _1572_/X VGND VGND VPWR VPWR _1614_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__2402__A _2402_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1545_ _1778_/A _1513_/A _1539_/A VGND VGND VPWR VPWR _1545_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__2759__D _2759_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1476_ _1803_/A _1803_/B _1803_/C _1803_/D VGND VGND VPWR VPWR _1807_/A sky130_fd_sc_hd__nand4_4
XANTENNA__2132__A1 input70/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2028_ _2727_/Q input42/X _2077_/S VGND VGND VPWR VPWR _2289_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2435__A2 _2428_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1643__B1 _1632_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2312__A _2312_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2669__D _2669_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1870__B _2931_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2123__A1 input68/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2426__A2 _1622_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2344__C_N _2329_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1634__B1 _1632_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output185_A _1932_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1330_ _1414_/C _1414_/D _1330_/C _1367_/B VGND VGND VPWR VPWR _1330_/X sky130_fd_sc_hd__and4_1
XFILLER_2_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput7 cpu_adr_i[14] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2417__A2 _1579_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1625__B1 _2787_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1301__A _1301_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1928__A1 input46/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2050__B1 _2049_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2715_ _2745_/CLK _2715_/D VGND VGND VPWR VPWR _2715_/Q sky130_fd_sc_hd__dfxtp_1
X_2646_ _2935_/Q _2136_/X _2140_/X VGND VGND VPWR VPWR _2935_/D sky130_fd_sc_hd__a21o_1
XANTENNA__1971__A _1971_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2577_ _2577_/A _2577_/B VGND VGND VPWR VPWR _2879_/D sky130_fd_sc_hd__nand2_1
X_1528_ _1528_/A _1528_/B VGND VGND VPWR VPWR _1562_/A sky130_fd_sc_hd__nor2_1
XANTENNA__2916__CLK _2920_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1459_ _1414_/A _1457_/X _1458_/Y _1500_/B VGND VGND VPWR VPWR _1459_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2105__A1 _2845_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1864__A0 _2755_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2307__A _2307_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1865__B _1865_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1395__A2 _1452_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1881__A _1889_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1607__B1 _1606_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2217__A _2217_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2862__D _2862_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2500_ _2500_/A _2508_/B VGND VGND VPWR VPWR _2827_/D sky130_fd_sc_hd__nand2_1
XANTENNA__2583__A1 _1567_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1386__A2 _1343_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2431_ _2451_/A VGND VGND VPWR VPWR _2431_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2939__CLK _2946_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2362_ _2362_/A VGND VGND VPWR VPWR _2382_/A sky130_fd_sc_hd__buf_2
XFILLER_57_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2293_ _2362_/A VGND VGND VPWR VPWR _2313_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__2098__S _2108_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1313_ _1422_/A _1297_/X _1424_/A VGND VGND VPWR VPWR _1479_/A sky130_fd_sc_hd__a21o_2
XFILLER_38_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1846__B1 _1845_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2772__D _2772_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2023__B1 _1994_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2056__A1_N _2906_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1377__A2 _1308_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput141 _1791_/Y VGND VGND VPWR VPWR spi_adr_o[0] sky130_fd_sc_hd__buf_2
Xoutput152 _1806_/Y VGND VGND VPWR VPWR spi_adr_o[1] sky130_fd_sc_hd__buf_2
X_2629_ _2629_/A _2631_/B VGND VGND VPWR VPWR _2920_/D sky130_fd_sc_hd__nor2_1
Xoutput130 _1767_/X VGND VGND VPWR VPWR cpu_dat_o[29] sky130_fd_sc_hd__buf_2
Xoutput163 _1812_/Y VGND VGND VPWR VPWR spi_adr_o[2] sky130_fd_sc_hd__buf_2
Xoutput185 _1932_/Y VGND VGND VPWR VPWR spi_dat_o[1] sky130_fd_sc_hd__buf_2
Xoutput174 _1925_/Y VGND VGND VPWR VPWR spi_dat_o[0] sky130_fd_sc_hd__buf_2
Xoutput196 _1940_/Y VGND VGND VPWR VPWR spi_dat_o[2] sky130_fd_sc_hd__buf_2
XFILLER_43_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1837__A0 _2344_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2682__D _2682_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1876__A _1878_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1368__A2 _1409_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2565__A1 _1495_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input61_A cpu_dat_i[4] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2500__A _2500_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2857__D _2857_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output148_A _1879_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1828__B1 _1789_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1931_ _2887_/Q _2573_/A _1927_/X _2487_/A VGND VGND VPWR VPWR _2590_/A sky130_fd_sc_hd__a2bb2o_2
XANTENNA__1786__A _2243_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1862_ _1807_/X _2548_/B _1789_/A _2929_/Q VGND VGND VPWR VPWR _2638_/B sky130_fd_sc_hd__o22ai_2
XANTENNA__2005__B1 _1975_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput10 cpu_adr_i[17] VGND VGND VPWR VPWR _1344_/A sky130_fd_sc_hd__clkbuf_1
Xinput21 cpu_adr_i[27] VGND VGND VPWR VPWR _1409_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2761__CLK _2768_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput54 cpu_dat_i[27] VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 cpu_dat_i[17] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_1
Xinput32 cpu_adr_i[8] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1359__A2 _1343_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1793_ _2092_/A VGND VGND VPWR VPWR _2474_/A sky130_fd_sc_hd__buf_2
Xinput98 spi_dat_i[31] VGND VGND VPWR VPWR input98/X sky130_fd_sc_hd__buf_2
Xinput87 spi_dat_i[21] VGND VGND VPWR VPWR input87/X sky130_fd_sc_hd__clkbuf_2
Xinput76 spi_dat_i[11] VGND VGND VPWR VPWR input76/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1764__C1 _1710_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput65 cpu_dat_i[8] VGND VGND VPWR VPWR input65/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2414_ _2408_/X _2410_/X _2413_/Y VGND VGND VPWR VPWR _2779_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__2410__A _2448_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2767__D _2767_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2345_ _2345_/A VGND VGND VPWR VPWR _2750_/D sky130_fd_sc_hd__clkbuf_1
X_2276_ _2324_/A VGND VGND VPWR VPWR _2296_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__1819__A0 _2747_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1598__A2 _1582_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1696__A _1696_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2547__A1 _2858_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1770__A2 _1569_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_21_CLK clkbuf_1_0_0_CLK/X VGND VGND VPWR VPWR _2764_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2320__A _2320_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2677__D _2677_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1691__D1 input83/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1589__A2 _1588_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2784__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1761__A2 _1760_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2230__A _2415_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_12_CLK clkbuf_1_1_0_CLK/X VGND VGND VPWR VPWR _2703_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2130_ _2884_/Q _1530_/X _1840_/X _2129_/Y VGND VGND VPWR VPWR _2586_/A sky130_fd_sc_hd__a2bb2o_2
X_2061_ _2837_/Q _2033_/X _2060_/X VGND VGND VPWR VPWR _2513_/A sky130_fd_sc_hd__o21ai_1
XFILLER_19_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_1_0_0_CLK_A clkbuf_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1914_ _2233_/A VGND VGND VPWR VPWR _1914_/X sky130_fd_sc_hd__buf_2
XANTENNA__2405__A _2451_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2894_ _2917_/CLK _2894_/D VGND VGND VPWR VPWR _2894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1845_ _2128_/A _1865_/B _2346_/A VGND VGND VPWR VPWR _1845_/X sky130_fd_sc_hd__or3_1
X_1776_ _2223_/A _2223_/B _1549_/X VGND VGND VPWR VPWR _1776_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__2140__A _2639_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1752__A2 _1751_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2328_ _2328_/A VGND VGND VPWR VPWR _2743_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1504__A2 _1426_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2259_ _2259_/A VGND VGND VPWR VPWR _2714_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2465__B1 _2464_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2315__A _2320_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1991__A2 _1961_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1743__A2 _1729_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input24_A cpu_adr_i[2] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1664__D1 input79/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_1_CLK clkbuf_1_0_0_CLK/X VGND VGND VPWR VPWR _2873_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2870__D _2870_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2225__A _2225_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1630_ _1630_/A VGND VGND VPWR VPWR _1630_/X sky130_fd_sc_hd__clkbuf_2
X_1561_ _1717_/A VGND VGND VPWR VPWR _1561_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__1734__A2 _1689_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1492_ _1445_/A _1488_/X _2866_/Q VGND VGND VPWR VPWR _1492_/Y sky130_fd_sc_hd__o21bai_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1498__B2 _1411_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1498__A1 _1495_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2113_ _2742_/Q input59/X _2113_/S VGND VGND VPWR VPWR _2325_/B sky130_fd_sc_hd__mux2_1
XFILLER_48_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1304__A _1304_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2044_ _2044_/A _2611_/A VGND VGND VPWR VPWR _2044_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2119__B _2128_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1670__A1 _1624_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2780__D _2780_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2946_ _2946_/CLK _2946_/D VGND VGND VPWR VPWR _2946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2877_ _2881_/CLK _2877_/D VGND VGND VPWR VPWR _2877_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1974__A _1980_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1828_ _1807_/X _2538_/B _1789_/X _2923_/Q VGND VGND VPWR VPWR _2632_/B sky130_fd_sc_hd__o22ai_2
X_1759_ _1723_/X _2533_/A _1709_/X _1710_/X input94/X VGND VGND VPWR VPWR _1759_/Y
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA__1725__A2 _1712_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_1_CLK_A clkbuf_1_0_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1489__A1 _1445_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2438__B1 _1656_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2029__B _2054_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1646__D1 input76/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2690__D _2690_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1661__A1 _1656_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2045__A _2076_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1884__A _1884_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2822__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1716__A2 _1682_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2141__A2 _2136_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2865__D _2865_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output130_A _1767_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2429__B1 _1625_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1652__A1 _1651_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2800_ _2809_/CLK _2800_/D VGND VGND VPWR VPWR _2800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2731_ _2834_/CLK _2731_/D VGND VGND VPWR VPWR _2731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1404__A1 _1379_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1794__A _1815_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2662_ _2665_/A _2944_/Q _2665_/C VGND VGND VPWR VPWR _2663_/A sky130_fd_sc_hd__and3_1
XFILLER_8_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2593_ _2593_/A _2593_/B VGND VGND VPWR VPWR _2890_/D sky130_fd_sc_hd__nor2_1
X_1613_ _1599_/X _1612_/X _2679_/Q VGND VGND VPWR VPWR _2171_/B sky130_fd_sc_hd__o21ai_1
X_1544_ _2152_/B _1543_/X _2672_/Q VGND VGND VPWR VPWR _1544_/Y sky130_fd_sc_hd__o21ai_1
X_1475_ _1717_/A VGND VGND VPWR VPWR _1778_/A sky130_fd_sc_hd__inv_2
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2775__D _2775_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1416__A2_N _1411_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1340__B1 _1339_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1628__D1 _1628_/D1 VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1969__A _2033_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2027_ _2027_/A VGND VGND VPWR VPWR _2077_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_63_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1643__A1 _1636_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2929_ _2929_/CLK _2929_/D VGND VGND VPWR VPWR _2929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2845__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2296__C_N _2281_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2685__D _2685_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1879__A _1879_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1619__D1 _1619_/D1 VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1634__A1 _1625_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input91_A spi_dat_i[25] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2503__A _2503_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output178_A _2011_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1570__B1 _2673_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput8 cpu_adr_i[15] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2718__CLK _2745_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1322__B1 _1321_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1789__A _1789_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2868__CLK _2873_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1625__A1 _1624_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2050__A1 _2835_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2714_ _2745_/CLK _2714_/D VGND VGND VPWR VPWR _2714_/Q sky130_fd_sc_hd__dfxtp_1
X_2645_ _2645_/A VGND VGND VPWR VPWR _2934_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1971__B _2008_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2576_ _2879_/Q _2493_/A _1311_/Y VGND VGND VPWR VPWR _2577_/B sky130_fd_sc_hd__o21ai_1
X_1527_ _1527_/A _1527_/B _1527_/C VGND VGND VPWR VPWR _1528_/A sky130_fd_sc_hd__nand3_2
X_1458_ _2389_/A _1452_/X _2757_/Q VGND VGND VPWR VPWR _1458_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2105__A2 _2251_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1864__A1 input4/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1313__B1 _1424_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1389_ _2863_/Q VGND VGND VPWR VPWR _1389_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1699__A _1699_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2323__A _2323_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1865__C _2355_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1881__B _2936_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1607__A1 _1604_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2568__C1 _2558_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2233__A _2233_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2583__A2 _1569_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1791__B1 _2628_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2430_ _2427_/X _2428_/X _2429_/Y VGND VGND VPWR VPWR _2787_/D sky130_fd_sc_hd__o21ai_1
XFILLER_29_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2361_ _2357_/X _2358_/X _1319_/Y _2382_/D VGND VGND VPWR VPWR _2756_/D sky130_fd_sc_hd__o211ai_1
X_2292_ _2292_/A VGND VGND VPWR VPWR _2728_/D sky130_fd_sc_hd__clkbuf_1
X_1312_ _2881_/Q VGND VGND VPWR VPWR _1424_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2085__A2_N _1914_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2690__CLK _2839_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1846__A1 _2856_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2408__A _2447_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1312__A _2881_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2023__A2_N _2018_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2143__A _2652_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2023__B2 _2505_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2559__C1 _2558_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1982__A _2046_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput142 _1863_/Y VGND VGND VPWR VPWR spi_adr_o[10] sky130_fd_sc_hd__buf_2
X_2628_ _2632_/A _2628_/B VGND VGND VPWR VPWR _2919_/D sky130_fd_sc_hd__nand2_1
Xoutput120 _1574_/X VGND VGND VPWR VPWR cpu_dat_o[1] sky130_fd_sc_hd__buf_2
Xoutput131 _1580_/X VGND VGND VPWR VPWR cpu_dat_o[2] sky130_fd_sc_hd__buf_2
XANTENNA__2334__C_N _2329_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput186 _2057_/Y VGND VGND VPWR VPWR spi_dat_o[20] sky130_fd_sc_hd__buf_2
Xoutput175 _1993_/Y VGND VGND VPWR VPWR spi_dat_o[10] sky130_fd_sc_hd__buf_2
Xoutput164 _1910_/X VGND VGND VPWR VPWR spi_adr_o[30] sky130_fd_sc_hd__buf_2
Xoutput153 _1888_/X VGND VGND VPWR VPWR spi_adr_o[20] sky130_fd_sc_hd__buf_2
X_2559_ _2357_/X _2358_/X _2370_/A _1489_/Y _2558_/X VGND VGND VPWR VPWR _2864_/D
+ sky130_fd_sc_hd__o311a_1
Xoutput197 _2112_/Y VGND VGND VPWR VPWR spi_dat_o[30] sky130_fd_sc_hd__buf_2
XFILLER_29_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1921__S _2132_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1837__A1 _2855_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2318__A _2318_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1876__B _2934_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2565__A2 _1497_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1892__A _1900_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1773__B1 _2809_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2500__B _2508_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input54_A cpu_dat_i[27] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1525__B1 _1500_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2101__A1_N _2914_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1831__S _2108_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1828__B2 _2923_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1828__A1 _1807_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output210_A _2949_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2873__D _2873_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2116__A1_N _2917_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1930_ _2817_/Q _2474_/A _1929_/X VGND VGND VPWR VPWR _2487_/A sky130_fd_sc_hd__o21ai_1
XFILLER_30_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1861_ _2353_/B _2859_/Q _2124_/S VGND VGND VPWR VPWR _2548_/B sky130_fd_sc_hd__mux2_1
XFILLER_14_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2906__CLK _2915_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2005__B2 _2004_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput11 cpu_adr_i[18] VGND VGND VPWR VPWR _1370_/A sky130_fd_sc_hd__clkbuf_1
Xinput22 cpu_adr_i[28] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1792_ _2064_/A VGND VGND VPWR VPWR _1792_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput55 cpu_dat_i[28] VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__buf_2
Xinput44 cpu_dat_i[18] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_1
Xinput33 cpu_adr_i[9] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_1
Xinput88 spi_dat_i[22] VGND VGND VPWR VPWR input88/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput77 spi_dat_i[12] VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1764__B1 _1709_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput66 cpu_dat_i[9] VGND VGND VPWR VPWR input66/X sky130_fd_sc_hd__clkbuf_1
Xinput99 spi_dat_i[3] VGND VGND VPWR VPWR input99/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2413_ _2412_/X _2160_/A _1560_/X VGND VGND VPWR VPWR _2413_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__1307__A _1371_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2344_ _2344_/A _2344_/B _2329_/X VGND VGND VPWR VPWR _2345_/A sky130_fd_sc_hd__or3b_1
XFILLER_57_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2275_ _2275_/A VGND VGND VPWR VPWR _2721_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1819__A1 input27/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2783__D _2783_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1977__A _2014_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2547__A2 _2540_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1755__B1 _2699_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2601__A _2601_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2320__B _2320_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1507__B1 _1392_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2180__B1 _2179_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2693__D _2693_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1887__A _1889_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1691__C1 _1638_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2929__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1746__B1 _1702_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2511__A _2511_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output160_A _1904_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2868__D _2868_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2060_ _2094_/A _2072_/B _2301_/B VGND VGND VPWR VPWR _2060_/X sky130_fd_sc_hd__or3_1
XFILLER_47_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1797__A _2065_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1913_ _1913_/A VGND VGND VPWR VPWR _2233_/A sky130_fd_sc_hd__buf_2
X_2893_ _2917_/CLK _2893_/D VGND VGND VPWR VPWR _2893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1844_ _2751_/Q input31/X _2127_/S VGND VGND VPWR VPWR _2346_/A sky130_fd_sc_hd__mux2_1
XANTENNA__1737__B1 _2696_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1775_ _1744_/X _1543_/A _2703_/Q VGND VGND VPWR VPWR _2223_/B sky130_fd_sc_hd__o21ai_1
XFILLER_7_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2778__D _2778_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2162__B1 _2156_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2327_ _2327_/A _2332_/B _2337_/C VGND VGND VPWR VPWR _2328_/A sky130_fd_sc_hd__and3_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2258_ _2272_/A _2258_/B _2257_/X VGND VGND VPWR VPWR _2259_/A sky130_fd_sc_hd__or3b_1
XFILLER_38_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2189_ _2189_/A _2189_/B VGND VGND VPWR VPWR _2190_/A sky130_fd_sc_hd__nand2_1
XFILLER_25_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2465__A1 _2447_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1500__A _2875_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1976__A0 _2719_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2315__B _2315_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1728__B1 _2801_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2331__A _2331_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2688__D _2688_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1847__A1_N _2926_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input17_A cpu_adr_i[23] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2751__CLK _2764_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1664__C1 _1638_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2506__A _2540_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1967__B1 _1916_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1719__B1 _2693_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1560_ _1558_/X _1559_/X _2779_/Q VGND VGND VPWR VPWR _1560_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2241__A _2540_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1491_ _1489_/Y _1358_/Y _1490_/Y _1335_/Y VGND VGND VPWR VPWR _1491_/Y sky130_fd_sc_hd__a22oi_2
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1498__A2 _1497_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2112_ _2117_/A _2625_/A VGND VGND VPWR VPWR _2112_/Y sky130_fd_sc_hd__nor2_4
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2545__C_N _2537_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2043_ _2904_/Q _2000_/X _2039_/X _2042_/Y VGND VGND VPWR VPWR _2611_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__2119__C _2238_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1655__C1 _1633_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2416__A _2558_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1670__A2 _1609_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2945_ _2946_/CLK _2945_/D VGND VGND VPWR VPWR _2945_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1958__B1 _1927_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2876_ _2880_/CLK _2876_/D VGND VGND VPWR VPWR _2876_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1974__B _2598_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1827_ _2339_/B _2853_/Q _2124_/S VGND VGND VPWR VPWR _2538_/B sky130_fd_sc_hd__mux2_1
XANTENNA__2151__A _2151_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1758_ _1707_/X _1559_/X _2806_/Q VGND VGND VPWR VPWR _1758_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1990__A _2014_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1689_ _1689_/A VGND VGND VPWR VPWR _1689_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2135__B1 _2587_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input9_A cpu_adr_i[16] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1489__A2 _1488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2774__CLK _2776_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2438__A1 _2433_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2029__C _2289_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1646__C1 _1627_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2326__A _2326_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1661__A2 _1660_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2126__B1 _2585_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1489__B1_N _2864_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2429__A1 _2412_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output123_A _1727_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2236__A _2312_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2881__D _2881_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1652__A2 _1588_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2730_ _2834_/CLK _2730_/D VGND VGND VPWR VPWR _2730_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1404__A2 _2401_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2661_ _2943_/Q _2649_/X _2650_/X VGND VGND VPWR VPWR _2943_/D sky130_fd_sc_hd__a21o_1
X_1612_ _1712_/A VGND VGND VPWR VPWR _1612_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2592_ _2592_/A _2638_/A VGND VGND VPWR VPWR _2889_/D sky130_fd_sc_hd__nand2_1
XANTENNA__2365__B1 _2227_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1543_ _1543_/A VGND VGND VPWR VPWR _1543_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2797__CLK _2839_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1474_ _2671_/Q VGND VGND VPWR VPWR _1717_/A sky130_fd_sc_hd__buf_4
XANTENNA__1315__A _1400_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1340__A1 _2871_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1628__C1 _1627_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2026_ _2114_/A VGND VGND VPWR VPWR _2078_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_63_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2791__D _2791_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2146__A _2526_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1643__A2 _1642_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1985__A _2035_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2928_ _2930_/CLK _2928_/D VGND VGND VPWR VPWR _2928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2859_ _2929_/CLK _2859_/D VGND VGND VPWR VPWR _2859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2108__A0 _2741_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1331__A1 _1424_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1619__C1 _1536_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1634__A2 _1631_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1895__A _1895_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input84_A spi_dat_i[19] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2503__B _2508_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1570__A1 _1567_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2876__D _2876_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1322__A1 _1479_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 cpu_adr_i[16] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1625__A2 _1609_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_0_CLK_A clkbuf_leaf_0_CLK/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2050__A2 _2033_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2713_ _2776_/CLK _2713_/D VGND VGND VPWR VPWR _2713_/Q sky130_fd_sc_hd__dfxtp_1
X_2644_ _2647_/A _2934_/Q _2653_/C VGND VGND VPWR VPWR _2645_/A sky130_fd_sc_hd__and3_1
X_2575_ _2878_/Q _2493_/A _2554_/X _1351_/Y VGND VGND VPWR VPWR _2878_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1971__C _2267_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1526_ _1490_/Y _1335_/Y _1493_/Y _1339_/Y VGND VGND VPWR VPWR _1527_/C sky130_fd_sc_hd__a22oi_4
XFILLER_59_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2786__D _2786_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1457_ _1457_/A VGND VGND VPWR VPWR _1457_/X sky130_fd_sc_hd__buf_2
XFILLER_56_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1313__A1 _1422_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1388_ _1388_/A _1388_/B VGND VGND VPWR VPWR _1788_/B sky130_fd_sc_hd__nor2_2
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2812__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2009_ _2829_/Q _1969_/X _2008_/X VGND VGND VPWR VPWR _2503_/A sky130_fd_sc_hd__o21ai_1
XFILLER_51_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2604__A _2604_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1537__D1 input74/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2696__D _2696_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1552__A1 _1744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1607__A2 _1605_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2568__B1 _1503_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2514__A _2531_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output190_A _2081_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1791__A1 _1779_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2360_ _2665_/C VGND VGND VPWR VPWR _2382_/D sky130_fd_sc_hd__buf_2
X_1311_ _1301_/Y _1457_/A _1309_/Y _1431_/A VGND VGND VPWR VPWR _1311_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_2_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2291_ _2296_/A _2291_/B _2281_/X VGND VGND VPWR VPWR _2292_/A sky130_fd_sc_hd__or3b_1
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2835__CLK _2839_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1700__D1 input84/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1846__A2 _1841_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2286__C_N _2281_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2559__B1 _1489_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput110 _1643_/X VGND VGND VPWR VPWR cpu_dat_o[10] sky130_fd_sc_hd__buf_2
Xoutput143 _1868_/Y VGND VGND VPWR VPWR spi_adr_o[11] sky130_fd_sc_hd__buf_2
X_2627_ _1781_/X _2527_/B _1481_/X _2626_/B VGND VGND VPWR VPWR _2918_/D sky130_fd_sc_hd__o211a_1
Xoutput132 _1772_/X VGND VGND VPWR VPWR cpu_dat_o[30] sky130_fd_sc_hd__buf_2
Xoutput121 _1715_/X VGND VGND VPWR VPWR cpu_dat_o[20] sky130_fd_sc_hd__buf_2
Xoutput165 _1912_/X VGND VGND VPWR VPWR spi_adr_o[31] sky130_fd_sc_hd__buf_2
Xoutput154 _1890_/X VGND VGND VPWR VPWR spi_adr_o[21] sky130_fd_sc_hd__buf_2
Xoutput176 _1999_/Y VGND VGND VPWR VPWR spi_dat_o[11] sky130_fd_sc_hd__buf_2
XFILLER_0_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2558_ _2558_/A VGND VGND VPWR VPWR _2558_/X sky130_fd_sc_hd__clkbuf_2
Xoutput187 _2063_/Y VGND VGND VPWR VPWR spi_dat_o[21] sky130_fd_sc_hd__buf_2
Xoutput198 _2117_/Y VGND VGND VPWR VPWR spi_dat_o[31] sky130_fd_sc_hd__buf_2
XFILLER_43_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2489_ _2818_/Q _2475_/X _1937_/X _2488_/X VGND VGND VPWR VPWR _2818_/D sky130_fd_sc_hd__o211a_1
X_1509_ _1509_/A _1509_/B VGND VGND VPWR VPWR _2573_/B sky130_fd_sc_hd__nand2_1
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1298__B1 _2767_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2318__B _2332_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2130__A2_N _1530_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1470__B1 _1469_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2334__A _2344_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2708__CLK _2873_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1892__B _2941_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1773__A1 _1707_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2858__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input47_A cpu_dat_i[20] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1525__B2 _1501_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1828__A2 _2538_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1413__A input6/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output203_A _1974_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1860_ _2754_/Q input3/X _1860_/S VGND VGND VPWR VPWR _2353_/B sky130_fd_sc_hd__mux2_1
XANTENNA__2244__A _2362_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1791_ _1779_/X _1781_/X _2628_/B VGND VGND VPWR VPWR _1791_/Y sky130_fd_sc_hd__a21oi_2
Xinput12 cpu_adr_i[19] VGND VGND VPWR VPWR _1360_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__1749__D1 input92/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput23 cpu_adr_i[29] VGND VGND VPWR VPWR _2395_/C sky130_fd_sc_hd__clkbuf_1
Xinput45 cpu_dat_i[19] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__clkbuf_1
Xinput34 cpu_cyc_i VGND VGND VPWR VPWR _1291_/A sky130_fd_sc_hd__buf_2
Xinput89 spi_dat_i[23] VGND VGND VPWR VPWR input89/X sky130_fd_sc_hd__clkbuf_2
Xinput78 spi_dat_i[13] VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1764__A1 _1717_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput56 cpu_dat_i[29] VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__clkbuf_2
Xinput67 cpu_sel_i[0] VGND VGND VPWR VPWR input67/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2412_ _2453_/A VGND VGND VPWR VPWR _2412_/X sky130_fd_sc_hd__clkbuf_2
X_2343_ _2343_/A VGND VGND VPWR VPWR _2749_/D sky130_fd_sc_hd__clkbuf_1
X_2274_ _2274_/A _2284_/B _2289_/C VGND VGND VPWR VPWR _2275_/A sky130_fd_sc_hd__and3_1
XFILLER_38_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1977__B _1990_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2301__C_N _2281_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1993__A _2011_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1989_ _2721_/Q input36/X _2013_/S VGND VGND VPWR VPWR _2274_/A sky130_fd_sc_hd__mux2_1
XANTENNA__1755__A1 _1744_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2601__B _2605_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1507__A1 _1389_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2180__A1 _1639_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2329__A _2352_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input101_A spi_dat_i[5] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1887__B _2939_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1691__B1 _1637_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2064__A _2064_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2680__CLK _2901_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1746__A1 _2211_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2511__B _2521_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output153_A _1888_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2884__D _2884_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2239__A _2239_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2037__A2_N _2018_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1912_ _1912_/A VGND VGND VPWR VPWR _1912_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2892_ _2917_/CLK _2892_/D VGND VGND VPWR VPWR _2892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1843_ _2027_/A VGND VGND VPWR VPWR _2127_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__1737__A1 _1692_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1774_ _1723_/A _1729_/X _1709_/A _1710_/A input98/X VGND VGND VPWR VPWR _2223_/A
+ sky130_fd_sc_hd__o2111ai_2
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2162__A1 _1577_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2326_ _2326_/A VGND VGND VPWR VPWR _2742_/D sky130_fd_sc_hd__clkbuf_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2257_ _2352_/A VGND VGND VPWR VPWR _2257_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2794__D _2794_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1988__A _2011_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2188_ _1664_/Y _1665_/Y _2179_/X VGND VGND VPWR VPWR _2686_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__2465__A2 _2448_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1673__B1 _2687_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1500__B _1500_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1976__A1 input65/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2612__A _2612_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1728__A1 _1696_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1898__A _1900_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1664__B1 _1637_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1416__B1 _1412_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1967__B2 _1966_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1837__S _2124_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1719__A1 _1672_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2879__D _2879_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2241__B _2241_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1490_ _1445_/X _1488_/X _2880_/Q VGND VGND VPWR VPWR _1490_/Y sky130_fd_sc_hd__o21bai_2
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2111_ _2916_/Q _2064_/X _1804_/X _2110_/Y VGND VGND VPWR VPWR _2625_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_48_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2042_ _2834_/Q _2025_/X _2041_/X VGND VGND VPWR VPWR _2042_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_63_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1655__B1 _1632_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2944_ _2946_/CLK _2944_/D VGND VGND VPWR VPWR _2944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1958__B2 _2492_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2080__B1 _2039_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2875_ _2881_/CLK _2875_/D VGND VGND VPWR VPWR _2875_/Q sky130_fd_sc_hd__dfxtp_1
X_1826_ _2243_/A VGND VGND VPWR VPWR _2124_/S sky130_fd_sc_hd__buf_2
XANTENNA__2789__D _2789_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1757_ _1753_/X _1756_/Y _1739_/X _1740_/X VGND VGND VPWR VPWR _1757_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1990__B _1990_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1688_ _1683_/X _1687_/Y _1667_/X _1668_/X VGND VGND VPWR VPWR _1688_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2919__CLK _2925_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2135__A1 _1859_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _2309_/A VGND VGND VPWR VPWR _2735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2438__A2 _2186_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2607__A _2607_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1646__B1 _1626_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1511__A _1511_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2071__A0 _2734_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2342__A _2342_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2699__D _2699_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2126__A1 _1859_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2069__A1_N _2908_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2429__A2 _2177_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output116_A _1681_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1421__A _1447_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2062__B1 _2058_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2660_ _2660_/A VGND VGND VPWR VPWR _2942_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2252__A _2272_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1611_ _1561_/X _1582_/X _1564_/X _1565_/X _1611_/D1 VGND VGND VPWR VPWR _2171_/A
+ sky130_fd_sc_hd__o2111ai_4
X_2591_ _2591_/A _2593_/B VGND VGND VPWR VPWR _2888_/D sky130_fd_sc_hd__nor2_1
XANTENNA__2365__A1 _2401_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1542_ _1568_/A VGND VGND VPWR VPWR _1543_/A sky130_fd_sc_hd__buf_4
X_1473_ _1739_/A VGND VGND VPWR VPWR _1473_/X sky130_fd_sc_hd__buf_6
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1315__B _1371_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1340__A2 _1324_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1628__B1 _1626_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2427__A _2447_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2025_ _2324_/A VGND VGND VPWR VPWR _2025_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2927_ _2930_/CLK _2927_/D VGND VGND VPWR VPWR _2927_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2053__A0 _2731_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1985__B _2008_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1800__A0 _2745_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2858_ _2929_/CLK _2858_/D VGND VGND VPWR VPWR _2858_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2741__CLK _2745_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1809_ _2746_/Q input24/X _1860_/S VGND VGND VPWR VPWR _2334_/B sky130_fd_sc_hd__mux2_1
X_2789_ _2847_/CLK _2789_/D VGND VGND VPWR VPWR _2789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2108__A1 input58/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2891__CLK _2917_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1867__B1 _1840_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1331__A2 _1380_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1619__B1 _1533_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2337__A _2337_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2072__A _2094_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input77_A spi_dat_i[12] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1570__A2 _1569_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1858__B1 _2637_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1850__S _2124_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1322__A2 _1319_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2892__D _2892_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2247__A _2540_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2764__CLK _2764_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2712_ _2745_/CLK _2712_/D VGND VGND VPWR VPWR _2712_/Q sky130_fd_sc_hd__dfxtp_1
X_2643_ _2933_/Q _2136_/X _2140_/X VGND VGND VPWR VPWR _2933_/D sky130_fd_sc_hd__a21o_1
X_2574_ _2574_/A VGND VGND VPWR VPWR _2877_/D sky130_fd_sc_hd__clkbuf_1
X_1525_ _1504_/Y _1327_/Y _1500_/Y _1501_/Y VGND VGND VPWR VPWR _1527_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_59_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1456_ _1407_/Y _1523_/A _1455_/Y VGND VGND VPWR VPWR _1461_/A sky130_fd_sc_hd__o21ai_1
X_1387_ _1443_/A _1387_/B _1387_/C _1387_/D VGND VGND VPWR VPWR _1388_/B sky130_fd_sc_hd__nand4b_1
XANTENNA__1849__A0 _2752_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1313__A2 _1297_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1996__A _2035_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2008_ _2035_/A _2008_/B _2282_/B VGND VGND VPWR VPWR _2008_/X sky130_fd_sc_hd__or3_1
XFILLER_51_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2604__B _2604_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2620__A _2650_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1537__C1 _1536_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1552__A2 _1568_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2067__A _2078_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2787__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2568__A1 _2401_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output183_A _2044_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1791__A2 _1781_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2530__A _2530_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2887__D _2887_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2290_ _2290_/A VGND VGND VPWR VPWR _2727_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1310_ _1350_/A VGND VGND VPWR VPWR _1431_/A sky130_fd_sc_hd__buf_4
XFILLER_38_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1700__C1 _1699_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2559__A1 _2357_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1767__C1 _1633_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2626_ _2626_/A _2626_/B VGND VGND VPWR VPWR _2917_/D sky130_fd_sc_hd__nand2_1
XANTENNA__2797__D _2797_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput133 _1777_/X VGND VGND VPWR VPWR cpu_dat_o[31] sky130_fd_sc_hd__buf_2
Xoutput122 _1721_/X VGND VGND VPWR VPWR cpu_dat_o[21] sky130_fd_sc_hd__buf_2
Xoutput111 _1649_/X VGND VGND VPWR VPWR cpu_dat_o[11] sky130_fd_sc_hd__buf_2
Xoutput177 _2006_/Y VGND VGND VPWR VPWR spi_dat_o[12] sky130_fd_sc_hd__buf_2
Xoutput155 _1893_/X VGND VGND VPWR VPWR spi_adr_o[22] sky130_fd_sc_hd__buf_2
Xoutput144 _1871_/X VGND VGND VPWR VPWR spi_adr_o[12] sky130_fd_sc_hd__buf_2
Xoutput166 _1823_/Y VGND VGND VPWR VPWR spi_adr_o[3] sky130_fd_sc_hd__buf_2
X_2557_ _2557_/A VGND VGND VPWR VPWR _2863_/D sky130_fd_sc_hd__clkbuf_1
Xoutput188 _2070_/Y VGND VGND VPWR VPWR spi_dat_o[22] sky130_fd_sc_hd__buf_2
Xoutput199 _1945_/Y VGND VGND VPWR VPWR spi_dat_o[3] sky130_fd_sc_hd__buf_2
X_1508_ _1508_/A _1508_/B _1508_/C _1508_/D VGND VGND VPWR VPWR _1512_/C sky130_fd_sc_hd__and4_1
X_2488_ _2531_/A VGND VGND VPWR VPWR _2488_/X sky130_fd_sc_hd__clkbuf_2
X_1439_ _1815_/A _1426_/X _2874_/Q VGND VGND VPWR VPWR _1510_/C sky130_fd_sc_hd__o21ai_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1298__A1 _1296_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2318__C _2337_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2615__A _2615_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1391__A_N input7/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2334__B _2334_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1470__A1 _1464_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2350__A _2350_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1773__A2 _1689_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2525__A _2525_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1790_ _2649_/A _2529_/B _1789_/X _2919_/Q VGND VGND VPWR VPWR _2628_/B sky130_fd_sc_hd__o22ai_2
Xinput13 cpu_adr_i[1] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__buf_2
XANTENNA__1749__C1 _1710_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput35 cpu_dat_i[0] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_1
Xinput46 cpu_dat_i[1] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__clkbuf_1
Xinput24 cpu_adr_i[2] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_1
Xinput79 spi_dat_i[14] VGND VGND VPWR VPWR input79/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1764__A2 _1729_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2260__A _2260_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput57 cpu_dat_i[2] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__clkbuf_1
Xinput68 cpu_sel_i[1] VGND VGND VPWR VPWR input68/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_15_CLK clkbuf_1_1_0_CLK/X VGND VGND VPWR VPWR _2834_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2802__CLK _2809_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2411_ _2706_/Q _1913_/A _1545_/Y _1467_/X _1469_/Y VGND VGND VPWR VPWR _2453_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2342_ _2342_/A _2355_/B _2370_/C VGND VGND VPWR VPWR _2343_/A sky130_fd_sc_hd__and3_1
X_2273_ _2273_/A VGND VGND VPWR VPWR _2720_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1977__C _2270_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1988_ _2011_/A _2600_/A VGND VGND VPWR VPWR _1988_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__1993__B _2601_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1755__A2 _1543_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2609_ _2609_/A _2617_/B VGND VGND VPWR VPWR _2902_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1507__A2 _1444_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2180__A2 _1641_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2468__B1 _2467_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1691__A1 _1651_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2345__A _2345_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2640__B1 _2140_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2825__CLK _2901_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1746__A2 _2211_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output146_A _1875_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1424__A _1424_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2459__B1 _2458_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_4_CLK clkbuf_1_0_0_CLK/X VGND VGND VPWR VPWR _2920_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2255__A _2255_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1911_ _1911_/A _2670_/Q VGND VGND VPWR VPWR _1912_/A sky130_fd_sc_hd__and2_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2891_ _2917_/CLK _2891_/D VGND VGND VPWR VPWR _2891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1842_ _2046_/A VGND VGND VPWR VPWR _2128_/A sky130_fd_sc_hd__buf_2
XFILLER_30_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1737__A2 _1712_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1773_ _1707_/A _1689_/A _2809_/Q VGND VGND VPWR VPWR _1773_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1318__B _1367_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2162__A2 _1578_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2325_ _2344_/A _2325_/B _2305_/X VGND VGND VPWR VPWR _2326_/A sky130_fd_sc_hd__or3b_1
XFILLER_57_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2256_ input1/X VGND VGND VPWR VPWR _2352_/A sky130_fd_sc_hd__buf_4
XANTENNA__1658__D1 input78/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1988__B _2600_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2187_ _2187_/A VGND VGND VPWR VPWR _2685_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1673__A1 _1672_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2165__A _2165_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2848__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2612__B _2616_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1509__A _1509_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1728__A2 _1682_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1361__B1 _2763_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1898__B _2944_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1664__A1 _1651_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2075__A _2075_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1998__A2_N _1953_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1416__B2 _1415_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1419__A _1568_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1719__A2 _1685_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2895__D _2895_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1352__B1 _1351_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2110_ _2846_/Q _1814_/X _2109_/X VGND VGND VPWR VPWR _2110_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2041_ _2078_/A _2054_/B _2294_/A VGND VGND VPWR VPWR _2041_/X sky130_fd_sc_hd__or3_1
XFILLER_63_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1655__A1 _1650_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2943_ _2946_/CLK _2943_/D VGND VGND VPWR VPWR _2943_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2080__B2 _2079_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2874_ _2881_/CLK _2874_/D VGND VGND VPWR VPWR _2874_/Q sky130_fd_sc_hd__dfxtp_1
X_1825_ _2748_/Q input28/X _1860_/S VGND VGND VPWR VPWR _2339_/B sky130_fd_sc_hd__mux2_1
X_1756_ _2215_/A _2215_/B _1702_/X VGND VGND VPWR VPWR _1756_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__1591__B1 _1549_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1687_ _2193_/A _2193_/B _1630_/X VGND VGND VPWR VPWR _1687_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__1990__C _2274_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2135__A2 _2649_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _2308_/A _2308_/B _2313_/C VGND VGND VPWR VPWR _2309_/A sky130_fd_sc_hd__and3_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1999__A _2011_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2239_ _2239_/A VGND VGND VPWR VPWR _2707_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2670__CLK _2670_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2607__B _2616_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1646__A1 _1645_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1511__B _2573_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2623__A _2623_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2071__A1 input50/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2342__B _2355_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2126__A2 _1853_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1334__B1 _2775_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input22_A cpu_adr_i[28] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1702__A _1702_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output109_A _1557_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2062__B2 _2513_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2533__A _2533_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2252__B _2252_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1610_ _1558_/X _1609_/X _2785_/Q VGND VGND VPWR VPWR _1610_/X sky130_fd_sc_hd__o21a_1
X_2590_ _2590_/A _2638_/A VGND VGND VPWR VPWR _2887_/D sky130_fd_sc_hd__nand2_1
XANTENNA__2365__A2 _2358_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1541_ _1692_/A VGND VGND VPWR VPWR _2152_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__1573__B1 _1572_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1472_ _2451_/A VGND VGND VPWR VPWR _1739_/A sky130_fd_sc_hd__clkinv_2
XFILLER_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1315__C _1401_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2522__C1 _2514_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2693__CLK _2703_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1612__A _1712_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2024_ _2044_/A _2607_/A VGND VGND VPWR VPWR _2024_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__1628__A1 _1561_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2926_ _2930_/CLK _2926_/D VGND VGND VPWR VPWR _2926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2053__A1 input47/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1985__C _2272_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2857_ _2925_/CLK _2857_/D VGND VGND VPWR VPWR _2857_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1800__A1 input13/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1808_ _2113_/S VGND VGND VPWR VPWR _1860_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_3_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2788_ _2847_/CLK _2788_/D VGND VGND VPWR VPWR _2788_/Q sky130_fd_sc_hd__dfxtp_1
X_1739_ _1739_/A VGND VGND VPWR VPWR _1739_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1867__B2 _1866_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1522__A _1723_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2618__A _2618_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1619__A1 _1576_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2337__B _2355_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2353__A _2353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2072__B _2072_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1555__B1 _1554_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2504__C1 _2501_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1858__A1 _1830_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2528__A _2528_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2247__B _2247_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2909__CLK _2915_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2263__A _2263_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2711_ _2776_/CLK _2711_/D VGND VGND VPWR VPWR _2711_/Q sky130_fd_sc_hd__dfxtp_1
X_2642_ _2642_/A VGND VGND VPWR VPWR _2932_/D sky130_fd_sc_hd__clkbuf_1
X_2573_ _2573_/A _2573_/B _2415_/A VGND VGND VPWR VPWR _2574_/A sky130_fd_sc_hd__or3b_1
XANTENNA__1546__B1 _2811_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1524_ _2879_/Q _2092_/A _1300_/Y _1311_/Y _2552_/A VGND VGND VPWR VPWR _1527_/A
+ sky130_fd_sc_hd__o2111a_1
X_1455_ _1500_/B _1455_/B _1455_/C VGND VGND VPWR VPWR _1455_/Y sky130_fd_sc_hd__nand3_1
XFILLER_56_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1386_ _2874_/Q _1343_/X _1385_/Y VGND VGND VPWR VPWR _1387_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__1849__A1 input32/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1342__A _1342_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2007_ _2724_/Q input39/X _2034_/S VGND VGND VPWR VPWR _2282_/B sky130_fd_sc_hd__mux2_1
XFILLER_24_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1996__B _2008_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2173__A _2173_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2909_ _2915_/CLK _2909_/D VGND VGND VPWR VPWR _2909_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1785__A0 _2744_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1537__B1 _1533_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1517__A _1707_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2348__A _2353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2067__B _2109_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2083__A _2094_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2568__A2 _2358_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1776__B1 _1549_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output176_A _1999_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_0_CLK CLK VGND VGND VPWR VPWR clkbuf_0_CLK/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__1861__S _2124_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2258__A _2272_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1700__B1 _1698_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2731__CLK _2834_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2559__A2 _2358_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2881__CLK _2881_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1767__B1 _1632_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2625_ _2625_/A _2631_/B VGND VGND VPWR VPWR _2916_/D sky130_fd_sc_hd__nor2_1
XANTENNA__1337__A _1337_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput123 _1727_/X VGND VGND VPWR VPWR cpu_dat_o[22] sky130_fd_sc_hd__buf_2
Xoutput112 _1655_/X VGND VGND VPWR VPWR cpu_dat_o[12] sky130_fd_sc_hd__buf_2
Xoutput134 _1586_/X VGND VGND VPWR VPWR cpu_dat_o[3] sky130_fd_sc_hd__buf_2
Xoutput156 _1895_/X VGND VGND VPWR VPWR spi_adr_o[23] sky130_fd_sc_hd__buf_2
Xoutput145 _1873_/X VGND VGND VPWR VPWR spi_adr_o[13] sky130_fd_sc_hd__buf_2
Xoutput167 _1829_/Y VGND VGND VPWR VPWR spi_adr_o[4] sky130_fd_sc_hd__buf_2
XANTENNA__2192__B1 _2179_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2556_ _2573_/A _2556_/B _2537_/X VGND VGND VPWR VPWR _2557_/A sky130_fd_sc_hd__or3b_1
Xoutput189 _2075_/Y VGND VGND VPWR VPWR spi_dat_o[23] sky130_fd_sc_hd__buf_2
Xoutput178 _2011_/Y VGND VGND VPWR VPWR spi_dat_o[13] sky130_fd_sc_hd__buf_2
X_2487_ _2487_/A _2495_/B VGND VGND VPWR VPWR _2817_/D sky130_fd_sc_hd__nand2_1
X_1507_ _1389_/Y _1444_/A _1392_/Y VGND VGND VPWR VPWR _1508_/A sky130_fd_sc_hd__o21a_1
X_1438_ _2765_/Q _1477_/A _1436_/Y _1500_/B VGND VGND VPWR VPWR _1442_/B sky130_fd_sc_hd__o211ai_1
XFILLER_56_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2168__A _2168_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1298__A2 _1297_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1369_ _1365_/Y _1324_/X _1368_/Y VGND VGND VPWR VPWR _1443_/A sky130_fd_sc_hd__o21ai_2
XFILLER_43_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2615__B _2617_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1470__A2 _1616_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2404__D1 _2403_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1758__B1 _2806_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2631__A _2631_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2350__B _2355_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1930__B1 _1929_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2078__A _2078_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2754__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1710__A _1710_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1997__B1 _1996_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2525__B _2525_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1749__B1 _1709_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput14 cpu_adr_i[20] VGND VGND VPWR VPWR _1366_/A sky130_fd_sc_hd__clkbuf_1
Xinput25 cpu_adr_i[30] VGND VGND VPWR VPWR _1301_/A sky130_fd_sc_hd__clkbuf_1
Xinput36 cpu_dat_i[10] VGND VGND VPWR VPWR input36/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2898__D _2898_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput58 cpu_dat_i[30] VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__buf_2
Xinput47 cpu_dat_i[20] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__clkbuf_1
Xinput69 cpu_sel_i[2] VGND VGND VPWR VPWR input69/X sky130_fd_sc_hd__buf_2
XANTENNA__2260__B _2260_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2410_ _2448_/A VGND VGND VPWR VPWR _2410_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2174__B1 _2156_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2341_ _2374_/A VGND VGND VPWR VPWR _2370_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__1921__A0 _2711_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2272_ _2272_/A _2272_/B _2257_/X VGND VGND VPWR VPWR _2273_/A sky130_fd_sc_hd__or3b_1
XANTENNA__2548__C_N _2537_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1620__A _1692_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1987_ _2895_/Q _1953_/X _1927_/X _2498_/A VGND VGND VPWR VPWR _2600_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2451__A _2451_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2608_ _2650_/A VGND VGND VPWR VPWR _2617_/B sky130_fd_sc_hd__clkbuf_2
X_2539_ _2539_/A VGND VGND VPWR VPWR _2853_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2777__CLK _2881_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2468__A1 _2447_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2626__A _2626_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1691__A2 _1663_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1530__A _1913_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1979__B1 _1975_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2640__A1 _2931_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input52_A cpu_dat_i[25] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1705__A _1740_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2459__A1 _2447_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output139_A _1623_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1440__A _1440_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1910_ _1910_/A VGND VGND VPWR VPWR _1910_/X sky130_fd_sc_hd__clkbuf_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2890_ _2917_/CLK _2890_/D VGND VGND VPWR VPWR _2890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1841_ _2033_/A VGND VGND VPWR VPWR _1841_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2271__A _2271_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1772_ _1768_/X _1771_/Y _1632_/A _1633_/A VGND VGND VPWR VPWR _1772_/X sky130_fd_sc_hd__o211a_4
XFILLER_7_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1318__C _1353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _2324_/A VGND VGND VPWR VPWR _2344_/A sky130_fd_sc_hd__buf_4
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2255_ _2255_/A VGND VGND VPWR VPWR _2713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1658__C1 _1627_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2186_ _2186_/A _2194_/B VGND VGND VPWR VPWR _2187_/A sky130_fd_sc_hd__or2_1
XANTENNA__1673__A2 _1612_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1350__A _1350_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2181__A _2181_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1509__B _1509_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2138__B1 _2537_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1361__A1 _1296_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1649__C1 _1633_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1664__A2 _1663_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2356__A _2356_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2075__B _2616_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2091__A _2102_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2942__CLK _2946_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2129__B1 _2128_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1352__A1 _2878_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2040_ _2729_/Q input44/X _2077_/S VGND VGND VPWR VPWR _2294_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2266__A _2266_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1655__A2 _1654_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2942_ _2946_/CLK _2942_/D VGND VGND VPWR VPWR _2942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2873_ _2873_/CLK _2873_/D VGND VGND VPWR VPWR _2873_/Q sky130_fd_sc_hd__dfxtp_1
X_1824_ _1853_/A VGND VGND VPWR VPWR _1824_/X sky130_fd_sc_hd__buf_2
X_1755_ _1744_/X _1543_/A _2699_/Q VGND VGND VPWR VPWR _2215_/B sky130_fd_sc_hd__o21ai_1
XFILLER_8_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1591__A1 _1589_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1686_ _1672_/X _1685_/X _2689_/Q VGND VGND VPWR VPWR _2193_/B sky130_fd_sc_hd__o21ai_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2307_ _2307_/A VGND VGND VPWR VPWR _2734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1999__B _2602_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2238_ _2238_/A _2260_/B _2386_/A VGND VGND VPWR VPWR _2239_/A sky130_fd_sc_hd__and3_1
XFILLER_54_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2815__CLK _2925_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1646__A2 _1582_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2169_ _2169_/A VGND VGND VPWR VPWR _2677_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2176__A _2198_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1511__C _1511_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2623__B _2631_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2342__C _2370_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1334__A1 _1296_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input15_A cpu_adr_i[21] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2086__A _2102_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1540_ _1744_/A VGND VGND VPWR VPWR _1692_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1864__S _2127_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1573__A1 _2158_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1471_ _2395_/A _2366_/A _1470_/Y VGND VGND VPWR VPWR _2451_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__2838__CLK _2840_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2522__B1 _2099_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1730__D1 input89/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2023_ _2901_/Q _2018_/X _1994_/X _2505_/A VGND VGND VPWR VPWR _2607_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__1628__A2 _1582_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2925_ _2925_/CLK _2925_/D VGND VGND VPWR VPWR _2925_/Q sky130_fd_sc_hd__dfxtp_1
X_2856_ _2929_/CLK _2856_/D VGND VGND VPWR VPWR _2856_/Q sky130_fd_sc_hd__dfxtp_1
X_1807_ _1807_/A VGND VGND VPWR VPWR _1807_/X sky130_fd_sc_hd__buf_2
X_2787_ _2847_/CLK _2787_/D VGND VGND VPWR VPWR _2787_/Q sky130_fd_sc_hd__dfxtp_1
X_1738_ _1736_/Y _1737_/Y _1679_/X VGND VGND VPWR VPWR _1738_/Y sky130_fd_sc_hd__a21oi_1
X_1669_ _1662_/X _1666_/Y _1667_/X _1668_/X VGND VGND VPWR VPWR _1669_/X sky130_fd_sc_hd__o211a_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input7_A cpu_adr_i[14] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1803__A _1803_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1619__A2 _1588_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2337__C _2337_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2634__A _2638_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2353__B _2353_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2072__C _2306_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1555__A1 _1548_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2504__B1 _2014_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1858__A2 _1853_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output121_A _1715_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1491__B1 _1490_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2440__C1 _2431_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2710_ _2873_/CLK _2710_/D VGND VGND VPWR VPWR _2710_/Q sky130_fd_sc_hd__dfxtp_1
X_2641_ _2647_/A _2932_/Q _2653_/C VGND VGND VPWR VPWR _2642_/A sky130_fd_sc_hd__and3_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1546__A1 _1463_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2572_ _2401_/C _2358_/A _2391_/A _1408_/Y _2558_/X VGND VGND VPWR VPWR _2876_/D
+ sky130_fd_sc_hd__o311a_1
X_1523_ _1523_/A VGND VGND VPWR VPWR _2092_/A sky130_fd_sc_hd__clkbuf_4
X_1454_ _1409_/A _1454_/B _1454_/C _1454_/D VGND VGND VPWR VPWR _1455_/C sky130_fd_sc_hd__nand4b_1
X_1385_ _1440_/A _1457_/A _1384_/Y _1362_/A VGND VGND VPWR VPWR _1385_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_56_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1342__B _1342_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2006_ _2011_/A _2603_/A VGND VGND VPWR VPWR _2006_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1482__B1 _1481_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1996__C _2277_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2908_ _2915_/CLK _2908_/D VGND VGND VPWR VPWR _2908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1785__A1 input2/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2839_ _2839_/CLK _2839_/D VGND VGND VPWR VPWR _2839_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1537__A1 _1902_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1533__A _1709_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2629__A _2629_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2348__B _2348_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2067__C _2303_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2364__A _2364_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2083__B _2114_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2568__A3 _2384_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input82_A spi_dat_i[17] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1776__A1 _2223_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2683__CLK _2901_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output169_A _1839_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2539__A _2539_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2489__C1 _2488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1443__A _1443_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2258__B _2258_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1700__A1 _1645_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1464__B1 _1463_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2274__A _2274_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2559__A3 _2370_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1767__A1 _1763_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2624_ _2624_/A _2626_/B VGND VGND VPWR VPWR _2915_/D sky130_fd_sc_hd__nand2_1
XANTENNA__1337__B _1390_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput124 _1733_/X VGND VGND VPWR VPWR cpu_dat_o[23] sky130_fd_sc_hd__buf_2
Xoutput113 _1661_/X VGND VGND VPWR VPWR cpu_dat_o[13] sky130_fd_sc_hd__buf_2
Xoutput157 _1897_/X VGND VGND VPWR VPWR spi_adr_o[24] sky130_fd_sc_hd__buf_2
Xoutput146 _1875_/X VGND VGND VPWR VPWR spi_adr_o[14] sky130_fd_sc_hd__buf_2
Xoutput168 _1835_/Y VGND VGND VPWR VPWR spi_adr_o[5] sky130_fd_sc_hd__buf_2
XANTENNA__2192__A1 _1677_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput135 _1596_/X VGND VGND VPWR VPWR cpu_dat_o[4] sky130_fd_sc_hd__buf_2
X_2555_ _1412_/X _1415_/X _2554_/X _2527_/A VGND VGND VPWR VPWR _2862_/D sky130_fd_sc_hd__o211a_1
Xoutput179 _2017_/Y VGND VGND VPWR VPWR spi_dat_o[14] sky130_fd_sc_hd__buf_2
X_2486_ _2510_/A VGND VGND VPWR VPWR _2495_/B sky130_fd_sc_hd__buf_2
X_1506_ _1500_/Y _1501_/Y _1502_/X _2552_/A _1505_/Y VGND VGND VPWR VPWR _1512_/B
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__1353__A _1353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1437_ _1437_/A VGND VGND VPWR VPWR _1500_/B sky130_fd_sc_hd__buf_2
XFILLER_29_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1368_ _2764_/Q _1409_/B _1367_/Y _1335_/C VGND VGND VPWR VPWR _1368_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_56_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1967__A1_N _2892_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2168__B _2172_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1299_ _1335_/C _2383_/A _2383_/B VGND VGND VPWR VPWR _1299_/Y sky130_fd_sc_hd__nand3_2
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2404__C1 _1469_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1758__A1 _1707_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2631__B _2631_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1528__A _1528_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2123__S _2132_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2350__C _2370_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1930__A1 _2817_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2359__A _2526_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2078__B _2109_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1694__B1 _1679_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2094__A _2094_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1446__B1 _2865_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1997__A1 _2827_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1749__A1 _1723_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput15 cpu_adr_i[21] VGND VGND VPWR VPWR _1376_/A sky130_fd_sc_hd__clkbuf_1
Xinput26 cpu_adr_i[31] VGND VGND VPWR VPWR _1333_/A sky130_fd_sc_hd__clkbuf_1
Xinput37 cpu_dat_i[11] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput59 cpu_dat_i[31] VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__buf_2
Xinput48 cpu_dat_i[21] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2260__C _2265_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2174__A1 _1619_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2340_ _2340_/A VGND VGND VPWR VPWR _2748_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2269__A _2362_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2271_ _2271_/A VGND VGND VPWR VPWR _2719_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1921__A1 input35/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1901__A _1901_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1986_ _2825_/Q _1969_/X _1985_/X VGND VGND VPWR VPWR _2498_/A sky130_fd_sc_hd__o21ai_1
XFILLER_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2005__A1_N _2898_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1348__A _2395_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2607_ _2607_/A _2616_/B VGND VGND VPWR VPWR _2901_/D sky130_fd_sc_hd__nand2_1
X_2538_ _2548_/A _2538_/B _2537_/X VGND VGND VPWR VPWR _2539_/A sky130_fd_sc_hd__or3b_1
XANTENNA__2179__A _2224_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2469_ _1768_/X _1771_/Y _2456_/X _2451_/A VGND VGND VPWR VPWR _2808_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2468__A2 _2448_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1676__B1 _2794_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2626__B _2626_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2118__S _2127_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1979__B2 _1978_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_986 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2640__A2 _2136_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2642__A _2642_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1600__B1 _2677_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2721__CLK _2745_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input45_A cpu_dat_i[19] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2459__A2 _2448_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2871__CLK _2873_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output201_A _1959_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2028__S _2077_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1440__B _1454_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1840_ _2039_/A VGND VGND VPWR VPWR _1840_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2552__A _2552_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2702__D _2702_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1771_ _1769_/Y _1770_/Y _1630_/A VGND VGND VPWR VPWR _1771_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__1318__D _1414_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _2323_/A VGND VGND VPWR VPWR _2741_/D sky130_fd_sc_hd__clkbuf_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2254_ _2254_/A _2260_/B _2265_/C VGND VGND VPWR VPWR _2255_/A sky130_fd_sc_hd__and3_1
XFILLER_38_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1658__B1 _1626_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2185_ _2185_/A _2185_/B VGND VGND VPWR VPWR _2186_/A sky130_fd_sc_hd__nand2_1
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2181__B _2181_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1969_ _2033_/A VGND VGND VPWR VPWR _1969_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2744__CLK _2873_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2138__A1 _1744_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2894__CLK _2917_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1346__C1 _1431_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1361__A2 _1297_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2637__A _2637_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1649__B1 _1632_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1541__A _1692_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2074__B1 _2058_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2372__A _2382_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1821__B1 _1820_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2538__C_N _2537_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2091__B _2621_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2129__A1 _2814_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output151_A _1886_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1352__A2 _1343_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1451__A _1451_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2941_ _2946_/CLK _2941_/D VGND VGND VPWR VPWR _2941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1812__B1 _2630_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2282__A _2296_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2767__CLK _2880_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2872_ _2880_/CLK _2872_/D VGND VGND VPWR VPWR _2872_/Q sky130_fd_sc_hd__dfxtp_1
X_1823_ _1779_/X _1781_/X _2631_/A VGND VGND VPWR VPWR _1823_/Y sky130_fd_sc_hd__a21oi_2
X_1754_ _1717_/X _1729_/X _1698_/X _1699_/X input93/X VGND VGND VPWR VPWR _2215_/A
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_8_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1626__A _1698_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1591__A2 _1590_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1685_ _1712_/A VGND VGND VPWR VPWR _1685_/X sky130_fd_sc_hd__clkbuf_2
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ _2320_/A _2306_/B _2305_/X VGND VGND VPWR VPWR _2307_/A sky130_fd_sc_hd__or3b_1
XFILLER_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2237_ _2374_/A VGND VGND VPWR VPWR _2386_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_39_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2168_ _2168_/A _2172_/B VGND VGND VPWR VPWR _2169_/A sky130_fd_sc_hd__or2_1
XFILLER_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2099_ _2109_/A _2109_/B _2318_/A VGND VGND VPWR VPWR _2099_/X sky130_fd_sc_hd__or3_2
XANTENNA__2056__B1 _2039_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1536__A _1710_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1970__S _1970_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1334__A2 _1297_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2086__B _2619_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output199_A _1945_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1573__A2 _2158_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1470_ _1464_/X _1616_/A _1469_/Y VGND VGND VPWR VPWR _1470_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2522__A1 _2844_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1730__C1 _1699_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2277__A _2296_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2022_ _2831_/Q _1969_/X _2021_/X VGND VGND VPWR VPWR _2505_/A sky130_fd_sc_hd__o21ai_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2924_ _2930_/CLK _2924_/D VGND VGND VPWR VPWR _2924_/Q sky130_fd_sc_hd__dfxtp_1
X_2855_ _2925_/CLK _2855_/D VGND VGND VPWR VPWR _2855_/Q sky130_fd_sc_hd__dfxtp_1
X_1806_ _1779_/X _1781_/X _2629_/A VGND VGND VPWR VPWR _1806_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__2210__B1 _2201_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2786_ _2847_/CLK _2786_/D VGND VGND VPWR VPWR _2786_/Q sky130_fd_sc_hd__dfxtp_1
X_1737_ _1692_/X _1712_/X _2696_/Q VGND VGND VPWR VPWR _1737_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__1356__A _1447_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1668_ _1740_/A VGND VGND VPWR VPWR _1668_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1599_ _1692_/A VGND VGND VPWR VPWR _1599_/X sky130_fd_sc_hd__clkbuf_2
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1803__B _1803_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1721__C1 _1705_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2932__CLK _2946_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2187__A _2187_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2634__B _2634_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2650__A _2650_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1555__A2 _1553_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2800__D _2800_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2504__A1 _2830_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2097__A _2102_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output114_A _1669_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1491__A1 _1489_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1491__B2 _1335_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2440__B1 _2436_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2640_ _2931_/Q _2136_/X _2140_/X VGND VGND VPWR VPWR _2931_/D sky130_fd_sc_hd__a21o_1
XANTENNA__2560__A _2577_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2805__CLK _2809_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2571_ _1500_/Y _1501_/Y _2495_/B VGND VGND VPWR VPWR _2875_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__2710__D _2710_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1522_ _1723_/A VGND VGND VPWR VPWR _1902_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1546__A2 _2527_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1453_ _2389_/A _1452_/X _2771_/Q VGND VGND VPWR VPWR _1455_/B sky130_fd_sc_hd__o21bai_1
XANTENNA__1904__A _1904_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1384_ _1451_/A _1452_/A _2769_/Q VGND VGND VPWR VPWR _1384_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_55_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2005_ _2898_/Q _2000_/X _1975_/X _2004_/Y VGND VGND VPWR VPWR _2603_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1482__A1 _1807_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2907_ _2915_/CLK _2907_/D VGND VGND VPWR VPWR _2907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1785__S _1785_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2838_ _2840_/CLK _2838_/D VGND VGND VPWR VPWR _2838_/Q sky130_fd_sc_hd__dfxtp_1
X_2769_ _2776_/CLK _2769_/D VGND VGND VPWR VPWR _2769_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1537__A2 _1530_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1814__A _2033_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2629__B _2631_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2645__A _2645_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2083__C _2310_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2422__B1 _2421_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2828__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1776__A2 _2223_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2380__A _2380_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input75_A spi_dat_i[10] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2489__B1 _1937_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1443__B _2562_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1700__A2 _1657_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2661__B1 _2650_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1464__A1 _1342_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2274__B _2284_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2705__D _2705_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2413__B1 _1560_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1767__A2 _1766_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_18_CLK clkbuf_1_1_0_CLK/X VGND VGND VPWR VPWR _2816_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2290__A _2290_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2623_ _2623_/A _2631_/B VGND VGND VPWR VPWR _2914_/D sky130_fd_sc_hd__nor2_1
Xoutput125 _1741_/X VGND VGND VPWR VPWR cpu_dat_o[24] sky130_fd_sc_hd__buf_2
Xoutput114 _1669_/X VGND VGND VPWR VPWR cpu_dat_o[14] sky130_fd_sc_hd__buf_2
X_2554_ _2558_/A VGND VGND VPWR VPWR _2554_/X sky130_fd_sc_hd__clkbuf_4
Xoutput158 _1899_/X VGND VGND VPWR VPWR spi_adr_o[25] sky130_fd_sc_hd__buf_2
Xoutput147 _1877_/X VGND VGND VPWR VPWR spi_adr_o[15] sky130_fd_sc_hd__buf_2
XANTENNA__2192__A2 _1678_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput136 _1602_/X VGND VGND VPWR VPWR cpu_dat_o[5] sky130_fd_sc_hd__buf_2
X_1505_ _1503_/Y _1299_/Y _1504_/Y _1327_/Y VGND VGND VPWR VPWR _1505_/Y sky130_fd_sc_hd__a22oi_4
Xoutput169 _1839_/Y VGND VGND VPWR VPWR spi_adr_o[6] sky130_fd_sc_hd__buf_2
X_2485_ _2816_/Q _2475_/X _1922_/X _2525_/B VGND VGND VPWR VPWR _2816_/D sky130_fd_sc_hd__o211a_1
X_1436_ _1436_/A _1454_/B _1454_/C _1454_/D VGND VGND VPWR VPWR _1436_/Y sky130_fd_sc_hd__nand4_1
XFILLER_29_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1367_ _1367_/A _1367_/B _1414_/C _1414_/D VGND VGND VPWR VPWR _1367_/Y sky130_fd_sc_hd__nand4_2
XFILLER_56_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1298_ _1296_/X _1297_/X _2767_/Q VGND VGND VPWR VPWR _2383_/B sky130_fd_sc_hd__o21ai_1
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2404__B1 _2231_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1758__A2 _1559_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1528__B _1528_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1930__A2 _2474_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2078__C _2308_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1694__A1 _1691_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_984 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2375__A _2375_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2643__B1 _2140_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2094__B _2114_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1446__A1 _1445_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1997__A2 _1969_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2096__A2_N _1914_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1749__A2 _2533_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput16 cpu_adr_i[22] VGND VGND VPWR VPWR _1337_/A sky130_fd_sc_hd__clkbuf_1
Xinput27 cpu_adr_i[3] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output181_A _2032_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput49 cpu_dat_i[22] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_1
Xinput38 cpu_dat_i[12] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2174__A2 _1621_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1382__B1 _1381_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2270_ _2270_/A _2284_/B _2289_/C VGND VGND VPWR VPWR _2271_/A sky130_fd_sc_hd__and3_1
XFILLER_42_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_CLK clkbuf_1_0_0_CLK/X VGND VGND VPWR VPWR _2670_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2285__A _2285_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1985_ _2035_/A _2008_/B _2272_/B VGND VGND VPWR VPWR _1985_/X sky130_fd_sc_hd__or3_1
XFILLER_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2606_ _2618_/A VGND VGND VPWR VPWR _2616_/B sky130_fd_sc_hd__clkbuf_2
X_2537_ _2537_/A VGND VGND VPWR VPWR _2537_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1373__B1 _2762_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1364__A _1423_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2570__C1 _1385_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2468_ _2447_/A _2448_/A _2467_/Y VGND VGND VPWR VPWR _2807_/D sky130_fd_sc_hd__o21ai_1
X_1419_ _1568_/A VGND VGND VPWR VPWR _2949_/A sky130_fd_sc_hd__inv_4
XFILLER_56_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2399_ _2399_/A _2401_/B _2399_/C VGND VGND VPWR VPWR _2400_/A sky130_fd_sc_hd__and3_1
XFILLER_56_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2673__CLK _2816_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1676__A1 _1635_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2195__A _2195_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1539__A _1539_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1600__A1 _1599_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2561__C1 _2558_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input38_A cpu_dat_i[12] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1440__C _1454_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1951__A1_N _2890_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2552__B _2552_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1770_ _1567_/X _1569_/X _2702_/Q VGND VGND VPWR VPWR _1770_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1449__A _1449_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2322_ _2322_/A _2332_/B _2337_/C VGND VGND VPWR VPWR _2323_/A sky130_fd_sc_hd__and3_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2696__CLK _2703_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1912__A _1912_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2253_ _2253_/A VGND VGND VPWR VPWR _2712_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1658__A1 _1645_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2184_ _1652_/Y _1653_/Y _2179_/X VGND VGND VPWR VPWR _2684_/D sky130_fd_sc_hd__a21oi_1
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1968_ _1980_/A _2597_/A VGND VGND VPWR VPWR _1968_/Y sky130_fd_sc_hd__nor2_1
X_1899_ _1899_/A VGND VGND VPWR VPWR _1899_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2138__A2 _1543_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1346__B1 _1345_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2637__B _2639_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1649__A1 _1644_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2653__A _2665_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2074__B2 _2516_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2051__A1_N _2905_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1821__A1 _2852_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2372__B _2372_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2803__D _2803_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1585__B1 _1572_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2129__A2 _1841_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output144_A _1871_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2940_ _2946_/CLK _2940_/D VGND VGND VPWR VPWR _2940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2563__A _2563_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1812__A1 _1779_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2282__B _2282_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2871_ _2873_/CLK _2871_/D VGND VGND VPWR VPWR _2871_/Q sky130_fd_sc_hd__dfxtp_1
X_1822_ _2922_/Q _1792_/X _1804_/X _1821_/Y VGND VGND VPWR VPWR _2631_/A sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2713__D _2713_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1753_ _1696_/X _1689_/A _2805_/Q VGND VGND VPWR VPWR _1753_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1907__A _1911_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1684_ _1645_/X _1657_/X _1626_/X _1627_/X input82/X VGND VGND VPWR VPWR _2193_/A
+ sky130_fd_sc_hd__o2111ai_4
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1328__B1 _1327_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _2352_/A VGND VGND VPWR VPWR _2305_/X sky130_fd_sc_hd__clkbuf_2
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2236_ _2312_/A VGND VGND VPWR VPWR _2260_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2167_ _2167_/A _2167_/B VGND VGND VPWR VPWR _2168_/A sky130_fd_sc_hd__nand2_1
XFILLER_41_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2098_ _2739_/Q input55/X _2108_/S VGND VGND VPWR VPWR _2318_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2056__B2 _2055_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2711__CLK _2776_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2861__CLK _2881_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1817__A _2065_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1319__B1 _1318_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2648__A _2648_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2383__A _2383_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2507__C1 _2501_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2558__A _2558_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2522__A2 _2519_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1730__B1 _1698_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1462__A _1803_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2277__B _2277_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2021_ _2035_/A _2072_/B _2286_/B VGND VGND VPWR VPWR _2021_/X sky130_fd_sc_hd__or3_1
XANTENNA__2708__D _2708_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2734__CLK _2834_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2293__A _2362_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2884__CLK _2920_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2923_ _2925_/CLK _2923_/D VGND VGND VPWR VPWR _2923_/Q sky130_fd_sc_hd__dfxtp_1
X_2854_ _2929_/CLK _2854_/D VGND VGND VPWR VPWR _2854_/Q sky130_fd_sc_hd__dfxtp_1
X_1805_ _2920_/Q _1792_/X _1802_/Y _1804_/X VGND VGND VPWR VPWR _2629_/A sky130_fd_sc_hd__a2bb2o_2
X_2785_ _2816_/CLK _2785_/D VGND VGND VPWR VPWR _2785_/Q sky130_fd_sc_hd__dfxtp_1
X_1736_ _1723_/X _2533_/A _1709_/X _1710_/X input90/X VGND VGND VPWR VPWR _1736_/Y
+ sky130_fd_sc_hd__o2111ai_2
XANTENNA__1637__A _1709_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2210__A1 _1736_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1356__B _1447_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1667_ _1739_/A VGND VGND VPWR VPWR _1667_/X sky130_fd_sc_hd__clkbuf_2
X_1598_ _1561_/X _1582_/X _1564_/X _1565_/X _1598_/D1 VGND VGND VPWR VPWR _2167_/A
+ sky130_fd_sc_hd__o2111ai_4
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1803__C _1803_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1372__A _1372_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1721__B1 _1704_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2219_ _2219_/A _2219_/B VGND VGND VPWR VPWR _2220_/A sky130_fd_sc_hd__nand2_1
XFILLER_27_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2504__A2 _2493_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2757__CLK _2764_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1282__A _2776_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2097__B _2622_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input20_A cpu_adr_i[26] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1491__A2 _1358_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2440__A1 _1662_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2560__B _2560_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1457__A _1457_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2570_ _2874_/Q _2493_/A _2554_/X _1385_/Y VGND VGND VPWR VPWR _2874_/D sky130_fd_sc_hd__o211a_1
X_1521_ _1717_/A VGND VGND VPWR VPWR _1723_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1951__B1 _1916_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1452_ _1452_/A VGND VGND VPWR VPWR _1452_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2288__A _2312_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1703__B1 _1702_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1383_ _1383_/A VGND VGND VPWR VPWR _1440_/A sky130_fd_sc_hd__inv_2
XFILLER_55_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2004_ _2828_/Q _1961_/X _2003_/X VGND VGND VPWR VPWR _2004_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__1920__A _2113_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1482__A2 _2527_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2906_ _2915_/CLK _2906_/D VGND VGND VPWR VPWR _2906_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2901__D _2901_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2837_ _2839_/CLK _2837_/D VGND VGND VPWR VPWR _2837_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1367__A _1367_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2768_ _2768_/CLK _2768_/D VGND VGND VPWR VPWR _2768_/Q sky130_fd_sc_hd__dfxtp_1
X_2699_ _2703_/CLK _2699_/D VGND VGND VPWR VPWR _2699_/Q sky130_fd_sc_hd__dfxtp_1
X_1719_ _1672_/X _1685_/X _2693_/Q VGND VGND VPWR VPWR _2203_/B sky130_fd_sc_hd__o21ai_1
XFILLER_2_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2198__A _2198_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1830__A _1859_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1976__S _2013_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2422__A1 _2408_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2380__B _2391_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2811__D _2811_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input68_A cpu_sel_i[1] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2489__A1 _2818_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1443__C _1443_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1740__A _1740_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2110__B1 _2109_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2661__A1 _2943_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2274__C _2289_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1464__A2 _1342_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2413__A1 _2412_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2721__D _2721_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2622_ _2622_/A _2626_/B VGND VGND VPWR VPWR _2913_/D sky130_fd_sc_hd__nand2_1
XANTENNA__2922__CLK _2930_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput115 _1675_/X VGND VGND VPWR VPWR cpu_dat_o[15] sky130_fd_sc_hd__buf_2
X_2553_ _2553_/A VGND VGND VPWR VPWR _2861_/D sky130_fd_sc_hd__clkbuf_1
Xoutput159 _1901_/X VGND VGND VPWR VPWR spi_adr_o[26] sky130_fd_sc_hd__buf_2
Xoutput148 _1879_/X VGND VGND VPWR VPWR spi_adr_o[16] sky130_fd_sc_hd__buf_2
XANTENNA__1924__B1 _1916_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1915__A _2039_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput126 _1747_/X VGND VGND VPWR VPWR cpu_dat_o[25] sky130_fd_sc_hd__buf_2
Xoutput137 _1608_/X VGND VGND VPWR VPWR cpu_dat_o[6] sky130_fd_sc_hd__buf_2
X_1504_ _1445_/X _1426_/X _2873_/Q VGND VGND VPWR VPWR _1504_/Y sky130_fd_sc_hd__o21bai_4
X_2484_ _2484_/A VGND VGND VPWR VPWR _2815_/D sky130_fd_sc_hd__clkbuf_1
X_1435_ _1815_/A _2019_/A _2870_/Q VGND VGND VPWR VPWR _1442_/A sky130_fd_sc_hd__o21ai_1
X_1366_ _1366_/A VGND VGND VPWR VPWR _1367_/A sky130_fd_sc_hd__clkinv_2
XANTENNA__1688__C1 _1668_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1297_ _1372_/A VGND VGND VPWR VPWR _1297_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_36_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2101__B1 _1804_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2481__A _2481_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2404__A1 _2395_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2656__A _2665_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1694__A2 _1693_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2375__B _2391_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2643__A1 _2933_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2094__C _2315_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1446__A2 _1426_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2806__D _2806_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2945__CLK _2946_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2391__A _2391_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput28 cpu_adr_i[4] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_1
Xinput17 cpu_adr_i[23] VGND VGND VPWR VPWR _1294_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_7_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput39 cpu_dat_i[13] VGND VGND VPWR VPWR input39/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_output174_A _1925_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1735__A _1735_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1454__B _1454_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1382__A1 _1479_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2716__D _2716_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1984_ _2720_/Q input66/X _2034_/S VGND VGND VPWR VPWR _2272_/B sky130_fd_sc_hd__mux2_1
XFILLER_9_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2605_ _2605_/A _2605_/B VGND VGND VPWR VPWR _2900_/D sky130_fd_sc_hd__nor2_1
XANTENNA__1645__A _1717_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1373__A1 _1451_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2536_ _2852_/Q _2519_/X _1820_/X _2531_/X VGND VGND VPWR VPWR _2852_/D sky130_fd_sc_hd__o211a_1
X_2467_ _2453_/X _2220_/A _1763_/X VGND VGND VPWR VPWR _2467_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__1364__B _1508_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2570__B1 _2554_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1418_ _1803_/A _1788_/B _1803_/D _2671_/Q VGND VGND VPWR VPWR _1568_/A sky130_fd_sc_hd__a31oi_4
XFILLER_56_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2398_ _2398_/A _2398_/B VGND VGND VPWR VPWR _2399_/A sky130_fd_sc_hd__nand2_1
XANTENNA__2818__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1349_ _1307_/X _1308_/X _2773_/Q VGND VGND VPWR VPWR _1349_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__1380__A _1380_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1676__A2 _1617_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1600__A2 _1569_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2561__B1 _1492_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2386__A _2386_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1290__A _1353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1440__D _1454_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1449__B _1449_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1465__A _1534_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2321_ _2321_/A VGND VGND VPWR VPWR _2740_/D sky130_fd_sc_hd__clkbuf_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2252_ _2272_/A _2252_/B _2227_/A VGND VGND VPWR VPWR _2253_/A sky130_fd_sc_hd__or3b_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1658__A2 _1657_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2183_ _2183_/A VGND VGND VPWR VPWR _2683_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2296__A _2296_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1967_ _2892_/Q _1933_/X _1916_/X _1966_/Y VGND VGND VPWR VPWR _2597_/A sky130_fd_sc_hd__a2bb2o_1
X_1898_ _1900_/A _2944_/Q VGND VGND VPWR VPWR _1899_/A sky130_fd_sc_hd__and2_1
XFILLER_49_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2080__A2_N _2064_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1346__A1 _1344_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2519_ _2540_/A VGND VGND VPWR VPWR _2519_/X sky130_fd_sc_hd__buf_2
XFILLER_57_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1649__A2 _1648_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2790__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2653__B _2938_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2372__C _2372_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1821__A2 _1814_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1984__S _2034_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1585__A1 _2163_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1285__A _1350_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input50_A cpu_dat_i[23] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_19_CLK_A clkbuf_1_0_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output137_A _1608_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1812__A2 _1781_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2870_ _2880_/CLK _2870_/D VGND VGND VPWR VPWR _2870_/Q sky130_fd_sc_hd__dfxtp_1
X_1821_ _2852_/Q _1814_/X _1820_/X VGND VGND VPWR VPWR _1821_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1752_ _1748_/X _1751_/Y _1739_/X _1740_/X VGND VGND VPWR VPWR _1752_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1907__B _2668_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1683_ _1624_/X _1682_/X _2795_/Q VGND VGND VPWR VPWR _1683_/X sky130_fd_sc_hd__o21a_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1328__A1 _2873_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ _2304_/A VGND VGND VPWR VPWR _2733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2111__A1_N _2916_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2235_ _2235_/A VGND VGND VPWR VPWR _2312_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_39_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2166_ _1589_/Y _1590_/Y _2156_/X VGND VGND VPWR VPWR _2676_/D sky130_fd_sc_hd__a21oi_1
XFILLER_54_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2097_ _2102_/A _2622_/A VGND VGND VPWR VPWR _2097_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_1044 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2904__D _2904_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1318__A_N input5/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1319__A1 _2756_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1724__D1 input88/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2383__B _2383_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2814__D _2814_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2452__C1 _2451_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2686__CLK _2901_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input98_A spi_dat_i[31] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2507__B1 _2029_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1730__A1 _1717_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1462__B _1803_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2020_ _2726_/Q input41/X _2034_/S VGND VGND VPWR VPWR _2286_/B sky130_fd_sc_hd__mux2_1
XFILLER_35_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1494__B1 _1493_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2574__A _2574_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2922_ _2930_/CLK _2922_/D VGND VGND VPWR VPWR _2922_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2724__D _2724_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2443__C1 _2431_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2853_ _2925_/CLK _2853_/D VGND VGND VPWR VPWR _2853_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1918__A _2046_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1804_ _2039_/A VGND VGND VPWR VPWR _1804_/X sky130_fd_sc_hd__clkbuf_2
X_2784_ _2847_/CLK _2784_/D VGND VGND VPWR VPWR _2784_/Q sky130_fd_sc_hd__dfxtp_1
X_1735_ _1735_/A VGND VGND VPWR VPWR _2533_/A sky130_fd_sc_hd__buf_6
XANTENNA__2210__A2 _1737_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1356__C input8/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1666_ _1664_/Y _1665_/Y _1606_/X VGND VGND VPWR VPWR _1666_/Y sky130_fd_sc_hd__a21oi_2
X_1597_ _1558_/X _1559_/X _2783_/Q VGND VGND VPWR VPWR _1597_/X sky130_fd_sc_hd__o21a_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1721__A1 _1716_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1803__D _1803_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2218_ _1759_/Y _1760_/Y _2201_/X VGND VGND VPWR VPWR _2700_/D sky130_fd_sc_hd__a21oi_1
X_2149_ _2669_/Q _2136_/X _2140_/X VGND VGND VPWR VPWR _2669_/D sky130_fd_sc_hd__a21o_1
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2484__A _2484_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2659__A _2665_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1563__A _1735_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2809__D _2809_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input13_A cpu_adr_i[1] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2440__A2 _1666_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1520_ _1517_/X _1519_/X _2778_/Q VGND VGND VPWR VPWR _1520_/X sky130_fd_sc_hd__o21a_1
XFILLER_45_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1951__B2 _1950_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1857__A1_N _2928_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1451_ _1451_/A VGND VGND VPWR VPWR _2389_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2701__CLK _2703_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1382_ _1479_/A _2380_/A _1381_/Y VGND VGND VPWR VPWR _1387_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__1473__A _1739_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1703__A1 _2197_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2719__D _2719_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2851__CLK _2925_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2003_ _2014_/A _2054_/B _2279_/A VGND VGND VPWR VPWR _2003_/X sky130_fd_sc_hd__or3_1
XFILLER_35_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2905_ _2915_/CLK _2905_/D VGND VGND VPWR VPWR _2905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2836_ _2840_/CLK _2836_/D VGND VGND VPWR VPWR _2836_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1367__B _1367_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2767_ _2880_/CLK _2767_/D VGND VGND VPWR VPWR _2767_/Q sky130_fd_sc_hd__dfxtp_1
X_1718_ _1717_/X _1657_/X _1698_/X _1699_/X input87/X VGND VGND VPWR VPWR _2203_/A
+ sky130_fd_sc_hd__o2111ai_4
X_2698_ _2703_/CLK _2698_/D VGND VGND VPWR VPWR _2698_/Q sky130_fd_sc_hd__dfxtp_1
X_1649_ _1644_/X _1648_/Y _1632_/X _1633_/X VGND VGND VPWR VPWR _1649_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1383__A _1383_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input5_A cpu_adr_i[12] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1458__B1 _2757_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2407__C1 _2537_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2422__A2 _2410_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1558__A _1696_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2380__C _2399_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2724__CLK _2745_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2389__A _2389_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1293__A _1355_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2874__CLK _2881_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2489__A2 _2475_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1697__B1 _2797_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2110__A1 _2846_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2661__A2 _2649_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1464__A3 _1528_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2413__A2 _2160_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1621__B1 _2680_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2621_ _2621_/A _2631_/B VGND VGND VPWR VPWR _2912_/D sky130_fd_sc_hd__nor2_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput116 _1681_/X VGND VGND VPWR VPWR cpu_dat_o[16] sky130_fd_sc_hd__buf_2
X_2552_ _2552_/A _2552_/B VGND VGND VPWR VPWR _2553_/A sky130_fd_sc_hd__or2_1
Xoutput149 _1882_/X VGND VGND VPWR VPWR spi_adr_o[17] sky130_fd_sc_hd__buf_2
XANTENNA__1924__B2 _1923_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2299__A _2299_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xoutput127 _1752_/X VGND VGND VPWR VPWR cpu_dat_o[26] sky130_fd_sc_hd__buf_2
Xoutput138 _1615_/X VGND VGND VPWR VPWR cpu_dat_o[7] sky130_fd_sc_hd__buf_2
XANTENNA__1385__C1 _1362_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1503_ _1445_/A _1488_/X _2872_/Q VGND VGND VPWR VPWR _1503_/Y sky130_fd_sc_hd__o21bai_2
X_2483_ _2529_/A _2483_/B _2352_/X VGND VGND VPWR VPWR _2484_/A sky130_fd_sc_hd__or3b_1
X_1434_ _1488_/A VGND VGND VPWR VPWR _2019_/A sky130_fd_sc_hd__buf_2
X_1365_ _2869_/Q VGND VGND VPWR VPWR _1365_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1688__B1 _1667_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1296_ _1371_/A VGND VGND VPWR VPWR _1296_/X sky130_fd_sc_hd__buf_2
XANTENNA__2101__B2 _2100_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1860__A0 _2754_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2912__D _2912_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2747__CLK _2768_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2404__A2 _2366_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2819_ _2920_/CLK _2819_/D VGND VGND VPWR VPWR _2819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2897__CLK _2901_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1841__A _2033_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2656__B _2940_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2375__C _2399_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2643__A2 _2136_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1851__B1 _1789_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2391__B _2391_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1288__A _1343_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2822__D _2822_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input80_A spi_dat_i[15] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput18 cpu_adr_i[24] VGND VGND VPWR VPWR _1325_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1603__B1 _2784_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput29 cpu_adr_i[5] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output167_A _1829_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1382__A2 _2380_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1454__C _1454_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2095__B1 _2094_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2582__A _2582_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1983_ _2047_/A VGND VGND VPWR VPWR _2034_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__2732__D _2732_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2604_ _2604_/A _2604_/B VGND VGND VPWR VPWR _2899_/D sky130_fd_sc_hd__nand2_1
XANTENNA__1926__A _2233_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2535_ _2535_/A VGND VGND VPWR VPWR _2851_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1373__A2 _1452_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2570__A1 _2874_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1364__C _1423_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2466_ _1758_/X _1761_/Y _2456_/X _2451_/X VGND VGND VPWR VPWR _2806_/D sky130_fd_sc_hd__o211a_1
X_1417_ _2556_/B _2560_/B _1461_/C _1417_/D VGND VGND VPWR VPWR _1803_/D sky130_fd_sc_hd__nor4_4
X_2397_ _1301_/Y _1457_/X _1309_/Y _2231_/A _2386_/A VGND VGND VPWR VPWR _2774_/D
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_3_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2907__D _2907_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1348_ _2395_/C VGND VGND VPWR VPWR _1348_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2492__A _2492_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1833__B1 _1832_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2010__B1 _1994_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2561__A1 _2357_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1571__A _1702_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2386__B _2386_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2912__CLK _2917_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2817__D _2817_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2077__A0 _2735_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1465__B _1534_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2320_ _2320_/A _2320_/B _2305_/X VGND VGND VPWR VPWR _2321_/A sky130_fd_sc_hd__or3b_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2251_ _2251_/A VGND VGND VPWR VPWR _2272_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2577__A _2577_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2182_ _2182_/A _2194_/B VGND VGND VPWR VPWR _2183_/A sky130_fd_sc_hd__or2_1
XANTENNA__2296__B _2296_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2727__D _2727_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2068__B1 _2067_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1966_ _2822_/Q _1961_/X _1965_/X VGND VGND VPWR VPWR _1966_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1897_ _1897_/A VGND VGND VPWR VPWR _1897_/X sky130_fd_sc_hd__clkbuf_1
X_2518_ _2518_/A _2521_/B VGND VGND VPWR VPWR _2841_/D sky130_fd_sc_hd__nand2_1
XFILLER_1_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1346__A2 _1457_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2487__A _2487_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2935__CLK _2946_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2449_ _2433_/X _2199_/A _1697_/X VGND VGND VPWR VPWR _2449_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2059__A0 _2732_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2653__C _2653_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1806__B1 _2629_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2372__D _2382_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1585__A2 _2163_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input43_A cpu_dat_i[17] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2470__B1 _1773_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1820_ _2109_/A _1865_/B _2337_/A VGND VGND VPWR VPWR _1820_/X sky130_fd_sc_hd__or3_1
XFILLER_31_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2808__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1751_ _1749_/Y _1750_/Y _1630_/A VGND VGND VPWR VPWR _1751_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__2222__B1 _2172_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1476__A _1803_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2071__S _2093_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1682_ _1682_/A VGND VGND VPWR VPWR _1682_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_7_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1328__A2 _1324_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ _2303_/A _2308_/B _2313_/C VGND VGND VPWR VPWR _2304_/A sky130_fd_sc_hd__and3_1
XANTENNA__1733__C1 _1705_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ _2706_/Q _2529_/A _1519_/X _2811_/Q _2577_/A VGND VGND VPWR VPWR _2706_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_39_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2165_ _2165_/A VGND VGND VPWR VPWR _2675_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2096_ _2913_/Q _1914_/X _2058_/X _2521_/A VGND VGND VPWR VPWR _2622_/A sky130_fd_sc_hd__a2bb2o_2
XFILLER_62_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2461__B1 _1742_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2920__D _2920_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1949_ _2364_/A _1990_/B _2260_/A VGND VGND VPWR VPWR _1949_/X sky130_fd_sc_hd__or3_1
XANTENNA__1319__A2 _1409_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1724__C1 _1710_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2452__B1 _2436_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1995__S _2034_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1296__A _1371_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2830__D _2830_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2507__A1 _2832_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1715__C1 _1705_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1730__A2 _1729_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1462__C _1462_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1494__B2 _1339_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1494__A1 _1492_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2066__S _2077_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2921_ _2925_/CLK _2921_/D VGND VGND VPWR VPWR _2921_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2443__B1 _2436_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2590__A _2590_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2852_ _2929_/CLK _2852_/D VGND VGND VPWR VPWR _2852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1803_ _1803_/A _1803_/B _1803_/C _1803_/D VGND VGND VPWR VPWR _2039_/A sky130_fd_sc_hd__and4_2
X_2783_ _2816_/CLK _2783_/D VGND VGND VPWR VPWR _2783_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2740__D _2740_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1734_ _1707_/X _1689_/X _2802_/Q VGND VGND VPWR VPWR _1734_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2780__CLK _2816_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1665_ _1620_/X _1640_/X _2686_/Q VGND VGND VPWR VPWR _1665_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__1356__D _1429_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1934__A _2019_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1596_ _1587_/X _1591_/Y _1593_/X _1595_/X VGND VGND VPWR VPWR _1596_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1706__C1 _1705_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1721__A2 _1720_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2217_ _2217_/A VGND VGND VPWR VPWR _2699_/D sky130_fd_sc_hd__clkbuf_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2148_ _2148_/A VGND VGND VPWR VPWR _2668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2915__D _2915_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2079_ _2840_/Q _2025_/X _2078_/X VGND VGND VPWR VPWR _2079_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_41_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2434__B1 _1644_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_leaf_18_CLK_A clkbuf_1_1_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2659__B _2942_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2825__D _2825_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2425__B1 _2424_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output197_A _2112_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1450_ _1389_/Y _1523_/A _1392_/Y _1508_/C VGND VGND VPWR VPWR _1462_/C sky130_fd_sc_hd__o211a_1
X_1381_ _1379_/X _1488_/A _2870_/Q VGND VGND VPWR VPWR _1381_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_45_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1703__A2 _2197_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2361__C1 _2382_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2585__A _2632_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2664__B1 _2650_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2002_ _2723_/Q input38/X _2013_/S VGND VGND VPWR VPWR _2279_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2735__D _2735_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1929__A _1971_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2904_ _2915_/CLK _2904_/D VGND VGND VPWR VPWR _2904_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2835_ _2839_/CLK _2835_/D VGND VGND VPWR VPWR _2835_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1367__C _1414_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2766_ _2768_/CLK _2766_/D VGND VGND VPWR VPWR _2766_/Q sky130_fd_sc_hd__dfxtp_1
X_1717_ _1717_/A VGND VGND VPWR VPWR _1717_/X sky130_fd_sc_hd__buf_4
X_2697_ _2703_/CLK _2697_/D VGND VGND VPWR VPWR _2697_/Q sky130_fd_sc_hd__dfxtp_1
X_1648_ _2181_/A _2181_/B _1630_/X VGND VGND VPWR VPWR _1648_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1979__A1_N _2894_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1579_ _1577_/Y _1578_/Y _1549_/X VGND VGND VPWR VPWR _1579_/Y sky130_fd_sc_hd__a21oi_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2676__CLK _2816_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2495__A _2495_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2655__B1 _2650_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1458__A1 _2389_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2407__B1 _1469_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1697__A1 _1696_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2646__B1 _2140_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2110__A2 _1814_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output112_A _1655_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1621__A1 _1620_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2620_ _2650_/A VGND VGND VPWR VPWR _2631_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__1484__A _2076_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1385__B1 _1384_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2551_ _1528_/A _1528_/B _2415_/A VGND VGND VPWR VPWR _2552_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__2699__CLK _2703_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2482_ _2814_/Q _2475_/X _2128_/X _2525_/B VGND VGND VPWR VPWR _2814_/D sky130_fd_sc_hd__o211a_1
Xoutput128 _1757_/X VGND VGND VPWR VPWR cpu_dat_o[27] sky130_fd_sc_hd__buf_2
Xoutput117 _1688_/X VGND VGND VPWR VPWR cpu_dat_o[17] sky130_fd_sc_hd__buf_2
Xoutput139 _1623_/X VGND VGND VPWR VPWR cpu_dat_o[8] sky130_fd_sc_hd__buf_2
X_1502_ _2879_/Q _1444_/A _1406_/B _1311_/Y VGND VGND VPWR VPWR _1502_/X sky130_fd_sc_hd__o211a_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1433_ _1510_/A _1510_/B VGND VGND VPWR VPWR _2562_/B sky130_fd_sc_hd__nand2_1
X_1364_ _1423_/A _1508_/B _1423_/C _1508_/D VGND VGND VPWR VPWR _1388_/A sky130_fd_sc_hd__nand4_2
XANTENNA__1688__A1 _1683_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1295_ _2776_/Q VGND VGND VPWR VPWR _1371_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2948__213 VGND VGND VPWR VPWR _2948__213/HI cpu_rty_o sky130_fd_sc_hd__conb_1
XFILLER_64_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1860__A1 input3/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2818_ _2847_/CLK _2818_/D VGND VGND VPWR VPWR _2818_/Q sky130_fd_sc_hd__dfxtp_1
X_2749_ _2768_/CLK _2749_/D VGND VGND VPWR VPWR _2749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1394__A input9/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2656__C _2665_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_976 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1300__B1 _1299_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1851__B2 _2927_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1851__A1 _1807_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1569__A _1712_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2391__C _2399_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1603__A1 _1517_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xinput19 cpu_adr_i[25] VGND VGND VPWR VPWR _1383_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_11_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input73_A spi_ack_i VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2841__CLK _2901_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2564__C1 _1362_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1454__D _1454_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2095__A1 _2843_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2582__B _2593_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1479__A _1479_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1982_ _2046_/A VGND VGND VPWR VPWR _2035_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2603_ _2603_/A _2605_/B VGND VGND VPWR VPWR _2898_/D sky130_fd_sc_hd__nor2_1
X_2534_ _2548_/A _2534_/B _2352_/X VGND VGND VPWR VPWR _2535_/A sky130_fd_sc_hd__or3b_1
XANTENNA__2555__C1 _2527_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2465_ _2447_/X _2448_/X _2464_/Y VGND VGND VPWR VPWR _2805_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__2570__A2 _2493_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1942__A _1971_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1364__D _1508_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2396_ _2773_/Q _1785_/S _2386_/D _2386_/A _2395_/X VGND VGND VPWR VPWR _2773_/D
+ sky130_fd_sc_hd__o2111a_1
X_1416_ _1408_/Y _1411_/Y _1412_/X _1415_/X VGND VGND VPWR VPWR _1417_/D sky130_fd_sc_hd__o2bb2ai_2
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1347_ _2866_/Q _1343_/X _1346_/Y VGND VGND VPWR VPWR _1423_/A sky130_fd_sc_hd__o21ai_1
XFILLER_3_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_924 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2714__CLK _2745_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2492__B _2495_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1833__A1 _2854_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2923__D _2923_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1389__A _2863_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2864__CLK _2880_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1597__B1 _2783_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1349__B1 _2773_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2010__B2 _2503_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2561__A2 _2358_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2386__C _2386_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2077__A1 input51/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2833__D _2833_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1299__A _1335_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1760__B1 _2700_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2250_ _2250_/A VGND VGND VPWR VPWR _2711_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2577__B _2577_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2181_ _2181_/A _2181_/B VGND VGND VPWR VPWR _2182_/A sky130_fd_sc_hd__nand2_1
XANTENNA__2737__CLK _2745_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2593__A _2593_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2068__A1 _2838_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2887__CLK _2920_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2743__D _2743_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2473__D1 _1470_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1965_ _2014_/A _1990_/B _2265_/A VGND VGND VPWR VPWR _1965_/X sky130_fd_sc_hd__or3_1
XANTENNA__1579__B1 _1549_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1937__A _2364_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1896_ _1900_/A _2943_/Q VGND VGND VPWR VPWR _1897_/A sky130_fd_sc_hd__and2_1
X_2517_ _2840_/Q _2506_/X _2078_/X _2514_/X VGND VGND VPWR VPWR _2840_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1751__B1 _1630_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1672__A _1744_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2448_ _2448_/A VGND VGND VPWR VPWR _2448_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2487__B _2495_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2918__D _2918_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1391__B _1429_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2379_ _1367_/A _1457_/X _1496_/Y _2231_/A _2386_/A VGND VGND VPWR VPWR _2764_/D
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2059__A1 input48/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1806__A1 _1779_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2008__A _2035_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1582__A _1735_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1742__B1 _2803_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2828__D _2828_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2330__C_N _2329_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input36_A cpu_dat_i[10] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2480__C_N _2352_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2470__A1 _2453_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1750_ _1692_/X _1712_/X _2698_/Q VGND VGND VPWR VPWR _1750_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2222__A1 _1769_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1476__B _1803_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1681_ _1676_/X _1680_/Y _1667_/X _1668_/X VGND VGND VPWR VPWR _1681_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2588__A _2588_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2302_ _2302_/A VGND VGND VPWR VPWR _2732_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1733__B1 _1704_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2738__D _2738_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2233_ _2233_/A VGND VGND VPWR VPWR _2529_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_54_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2164_ _2164_/A _2172_/B VGND VGND VPWR VPWR _2165_/A sky130_fd_sc_hd__or2_1
XANTENNA__1497__C1 _1287_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2095_ _2843_/Q _2251_/A _2094_/X VGND VGND VPWR VPWR _2521_/A sky130_fd_sc_hd__o21ai_2
XFILLER_62_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2461__A1 _2453_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1667__A _1739_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1948_ _2715_/Q input61/X _2132_/S VGND VGND VPWR VPWR _2260_/A sky130_fd_sc_hd__mux2_1
X_1879_ _1879_/A VGND VGND VPWR VPWR _1879_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2902__CLK _2915_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1972__B1 _1971_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2498__A _2498_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2353__C_N _2352_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1724__B1 _1709_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2452__A1 _1708_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2507__A2 _2506_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1715__B1 _1704_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2201__A _2224_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output142_A _1863_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1462__D _1462_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1494__A2 _1346_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2920_ _2920_/CLK _2920_/D VGND VGND VPWR VPWR _2920_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2443__A1 _1676_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2590__B _2638_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2082__S _2093_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2851_ _2925_/CLK _2851_/D VGND VGND VPWR VPWR _2851_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2925__CLK _2925_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2782_ _2847_/CLK _2782_/D VGND VGND VPWR VPWR _2782_/Q sky130_fd_sc_hd__dfxtp_1
X_1802_ _2850_/Q _2474_/A _1801_/X VGND VGND VPWR VPWR _1802_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1387__A_N _1443_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1733_ _1728_/X _1732_/Y _1704_/X _1705_/X VGND VGND VPWR VPWR _1733_/X sky130_fd_sc_hd__o211a_1
X_1664_ _1651_/X _1663_/X _1637_/X _1638_/X input79/X VGND VGND VPWR VPWR _1664_/Y
+ sky130_fd_sc_hd__o2111ai_2
X_1595_ _1633_/A VGND VGND VPWR VPWR _1595_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1706__B1 _1704_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ _2216_/A _2216_/B VGND VGND VPWR VPWR _2217_/A sky130_fd_sc_hd__or2_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2131__B1 _2586_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2147_ _2647_/A _2668_/Q _2401_/B VGND VGND VPWR VPWR _2148_/A sky130_fd_sc_hd__and3_1
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2078_ _2078_/A _2109_/B _2308_/A VGND VGND VPWR VPWR _2078_/X sky130_fd_sc_hd__or3_1
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2434__A1 _2433_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2931__D _2931_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2659__C _2665_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2021__A _2035_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2122__B1 _2582_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2425__A1 _2408_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2841__D _2841_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1936__A0 _2713_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1380_ _1380_/A VGND VGND VPWR VPWR _1488_/A sky130_fd_sc_hd__buf_2
XANTENNA__2361__B1 _1319_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2585__B _2585_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2113__A0 _2742_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2001_ _2065_/A VGND VGND VPWR VPWR _2054_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_64_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2664__A1 _2945_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2077__S _2077_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2903_ _2915_/CLK _2903_/D VGND VGND VPWR VPWR _2903_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2751__D _2751_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1929__B _2128_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1931__A2_N _2573_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2834_ _2834_/CLK _2834_/D VGND VGND VPWR VPWR _2834_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1367__D _1414_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1945__A _1945_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2765_ _2768_/CLK _2765_/D VGND VGND VPWR VPWR _2765_/Q sky130_fd_sc_hd__dfxtp_2
X_2696_ _2703_/CLK _2696_/D VGND VGND VPWR VPWR _2696_/Q sky130_fd_sc_hd__dfxtp_1
X_1716_ _1696_/X _1682_/X _2799_/Q VGND VGND VPWR VPWR _1716_/X sky130_fd_sc_hd__o21a_1
X_1647_ _1599_/X _1612_/X _2683_/Q VGND VGND VPWR VPWR _2181_/B sky130_fd_sc_hd__o21ai_1
XFILLER_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1578_ _2152_/B _1543_/X _2674_/Q VGND VGND VPWR VPWR _1578_/Y sky130_fd_sc_hd__o21ai_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2495__B _2495_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2655__A1 _2939_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2926__D _2926_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1458__A2 _1452_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2407__A1 _1464_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1615__C1 _1595_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1855__A _2128_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1697__A2 _1682_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2646__A1 _2935_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2770__CLK _2776_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2836__D _2836_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2031__A2_N _2000_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1621__A2 _1543_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2550_ _2860_/Q _2540_/X _1865_/X _2510_/A VGND VGND VPWR VPWR _2860_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1385__A1 _1440_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2481_ _2481_/A VGND VGND VPWR VPWR _2813_/D sky130_fd_sc_hd__clkbuf_1
Xoutput129 _1762_/X VGND VGND VPWR VPWR cpu_dat_o[28] sky130_fd_sc_hd__buf_2
Xoutput118 _1695_/X VGND VGND VPWR VPWR cpu_dat_o[18] sky130_fd_sc_hd__buf_2
X_1501_ _1330_/C _1477_/A _1329_/X _1479_/A VGND VGND VPWR VPWR _1501_/Y sky130_fd_sc_hd__a211oi_2
X_1432_ _2762_/Q _1477_/A _1430_/Y _1444_/A VGND VGND VPWR VPWR _1510_/B sky130_fd_sc_hd__o211ai_1
XANTENNA__2596__A _2650_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1363_ _2868_/Q _1324_/X _1362_/Y VGND VGND VPWR VPWR _1508_/D sky130_fd_sc_hd__o21ai_2
XANTENNA__1688__A2 _1687_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1294_ _1414_/C _1354_/A _1294_/C _1367_/B VGND VGND VPWR VPWR _2383_/A sky130_fd_sc_hd__nand4_4
XANTENNA_clkbuf_leaf_17_CLK_A clkbuf_1_1_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2746__D _2746_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2817_ _2920_/CLK _2817_/D VGND VGND VPWR VPWR _2817_/Q sky130_fd_sc_hd__dfxtp_1
X_2748_ _2873_/CLK _2748_/D VGND VGND VPWR VPWR _2748_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1394__B _1409_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2679_ _2816_/CLK _2679_/D VGND VGND VPWR VPWR _2679_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2793__CLK _2839_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1300__A1 _2872_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1851__A2 _2545_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1603__A2 _1519_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input66_A cpu_dat_i[9] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2564__B1 _2554_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1524__D1 _2552_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2095__A2 _2251_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1981_ _2117_/A VGND VGND VPWR VPWR _2011_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2602_ _2602_/A _2604_/B VGND VGND VPWR VPWR _2897_/D sky130_fd_sc_hd__nand2_1
X_2533_ _2533_/A VGND VGND VPWR VPWR _2548_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2555__B1 _2554_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2464_ _2453_/X _2216_/A _1753_/X VGND VGND VPWR VPWR _2464_/Y sky130_fd_sc_hd__a21oi_1
X_1415_ _2757_/Q _1428_/A _1414_/Y _1362_/A VGND VGND VPWR VPWR _1415_/X sky130_fd_sc_hd__o211a_1
X_2395_ _2395_/A _2395_/B _2395_/C _2395_/D VGND VGND VPWR VPWR _2395_/X sky130_fd_sc_hd__or4_1
XANTENNA__1942__B _2128_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1346_ _1344_/Y _1457_/A _1345_/Y _1431_/A VGND VGND VPWR VPWR _1346_/Y sky130_fd_sc_hd__o211ai_4
XFILLER_3_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1833__A2 _1814_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2491__C1 _2488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1597__A1 _1558_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1349__A1 _1307_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1754__D1 input93/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2561__A3 _2375_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1506__D1 _1505_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2386__D _2386_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2482__C1 _2525_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2689__CLK _2839_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1299__B _2383_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2234__C1 _2577_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2204__A _2204_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output172_A _1858_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1760__A1 _1567_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2016__A1_N _2900_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2180_ _1639_/Y _1641_/Y _2179_/X VGND VGND VPWR VPWR _2682_/D sky130_fd_sc_hd__a21oi_1
XFILLER_38_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2593__B _2593_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2068__A2 _2025_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2473__C1 _2366_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1579__A1 _1577_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1964_ _2717_/Q input63/X _2013_/S VGND VGND VPWR VPWR _2265_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1937__B _1990_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1895_ _1895_/A VGND VGND VPWR VPWR _1895_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2114__A _2114_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1953__A _2233_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1736__D1 input90/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2516_ _2516_/A _2521_/B VGND VGND VPWR VPWR _2839_/D sky130_fd_sc_hd__nand2_1
XANTENNA__1751__A1 _1749_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2447_ _2447_/A VGND VGND VPWR VPWR _2447_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1391__C _1447_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2378_ _1362_/B _1362_/C _2365_/Y VGND VGND VPWR VPWR _2763_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__1503__A1 _1445_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1329_ _1400_/A _1371_/A _1401_/A _2770_/Q VGND VGND VPWR VPWR _1329_/X sky130_fd_sc_hd__o31a_2
XANTENNA__2831__CLK _2901_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2934__D _2934_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1806__A2 _1781_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2282__C_N _2281_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2008__B _2008_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2024__A _2044_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1742__A1 _1696_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input29_A cpu_adr_i[5] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2844__D _2844_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2470__A2 _2224_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2222__A2 _1770_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1476__C _1803_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1680_ _1677_/Y _1678_/Y _1679_/X VGND VGND VPWR VPWR _1680_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_7_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2588__B _2593_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1718__D1 input87/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2704__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2301_ _2320_/A _2301_/B _2281_/X VGND VGND VPWR VPWR _2302_/A sky130_fd_sc_hd__or3b_1
XANTENNA__1733__A1 _1728_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2232_ _2811_/Q _1464_/X _1545_/Y _1467_/X _2577_/A VGND VGND VPWR VPWR _2705_/D
+ sky130_fd_sc_hd__o221a_1
XANTENNA__2854__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2163_ _2163_/A _2163_/B VGND VGND VPWR VPWR _2164_/A sky130_fd_sc_hd__nand2_1
XANTENNA__1497__B1 _1496_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2754__D _2754_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2094_ _2094_/A _2114_/B _2315_/B VGND VGND VPWR VPWR _2094_/X sky130_fd_sc_hd__or3_1
XFILLER_62_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2109__A _2109_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2446__C1 _2431_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2461__A2 _2212_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1947_ _2117_/A VGND VGND VPWR VPWR _1980_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1878_ _1878_/A _2935_/Q VGND VGND VPWR VPWR _1879_/A sky130_fd_sc_hd__and2_1
XANTENNA__1972__A1 _2823_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1724__A1 _1723_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2498__B _2508_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2929__D _2929_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2019__A _2019_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2437__C1 _2431_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2452__A2 _1714_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1660__B1 _1630_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2727__CLK _2834_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1412__B1 _2862_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1593__A _1632_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2839__D _2839_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2877__CLK _2881_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1715__A1 _1708_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output135_A _1596_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2443__A2 _1680_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2850_ _2929_/CLK _2850_/D VGND VGND VPWR VPWR _2850_/Q sky130_fd_sc_hd__dfxtp_1
X_1801_ _1971_/A _2128_/B _2332_/A VGND VGND VPWR VPWR _1801_/X sky130_fd_sc_hd__or3_2
X_2781_ _2816_/CLK _2781_/D VGND VGND VPWR VPWR _2781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1732_ _2207_/A _2207_/B _1702_/X VGND VGND VPWR VPWR _1732_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2599__A _2599_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1663_ _1913_/A VGND VGND VPWR VPWR _1663_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__2749__D _2749_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1594_ _1740_/A VGND VGND VPWR VPWR _1633_/A sky130_fd_sc_hd__buf_2
XANTENNA__1706__A1 _1697_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2215_ _2215_/A _2215_/B VGND VGND VPWR VPWR _2216_/A sky130_fd_sc_hd__nand2_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2131__A1 _1859_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2146_ _2526_/A VGND VGND VPWR VPWR _2401_/B sky130_fd_sc_hd__buf_4
XFILLER_54_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2077_ _2735_/Q input51/X _2077_/S VGND VGND VPWR VPWR _2308_/A sky130_fd_sc_hd__mux2_1
XANTENNA__2434__A2 _2182_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1642__B1 _1606_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2320__C_N _2305_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2302__A _2302_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2021__B _2072_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2122__A1 _1859_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1588__A _1913_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2425__A2 _2410_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input96_A spi_dat_i[2] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1936__A1 input57/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2212__A _2212_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2361__A1 _2357_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2000_ _2064_/A VGND VGND VPWR VPWR _2000_/X sky130_fd_sc_hd__buf_2
XANTENNA__2113__A1 input59/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2664__A2 _2649_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2902_ _2915_/CLK _2902_/D VGND VGND VPWR VPWR _2902_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2093__S _2093_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1929__C _2252_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2833_ _2901_/CLK _2833_/D VGND VGND VPWR VPWR _2833_/Q sky130_fd_sc_hd__dfxtp_1
X_2764_ _2764_/CLK _2764_/D VGND VGND VPWR VPWR _2764_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1945__B _2592_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1715_ _1708_/X _1714_/Y _1704_/X _1705_/X VGND VGND VPWR VPWR _1715_/X sky130_fd_sc_hd__o211a_1
X_2695_ _2703_/CLK _2695_/D VGND VGND VPWR VPWR _2695_/Q sky130_fd_sc_hd__dfxtp_1
X_1646_ _1645_/X _1582_/X _1626_/X _1627_/X input76/X VGND VGND VPWR VPWR _2181_/A
+ sky130_fd_sc_hd__o2111ai_4
X_1577_ _1576_/X _1530_/X _1533_/X _1536_/X input96/X VGND VGND VPWR VPWR _1577_/Y
+ sky130_fd_sc_hd__o2111ai_2
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1961__A _2324_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2655__A2 _2649_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1863__B1 _2638_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2129_ _2814_/Q _1841_/X _2128_/X VGND VGND VPWR VPWR _2129_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_15_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2942__D _2942_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2407__A2 _1682_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1615__B1 _1593_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2040__A0 _2729_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1855__B _1865_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2032__A _2044_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1871__A _1871_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2915__CLK _2915_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2646__A2 _2136_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input11_A cpu_adr_i[18] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1854__A0 _2753_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1810__S _2374_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2852__D _2852_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2207__A _2207_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2031__B1 _1975_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1385__A2 _1457_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2480_ _2529_/A _2480_/B _2352_/X VGND VGND VPWR VPWR _2481_/A sky130_fd_sc_hd__or3b_1
Xoutput119 _1706_/X VGND VGND VPWR VPWR cpu_dat_o[19] sky130_fd_sc_hd__buf_2
Xoutput108 _1473_/X VGND VGND VPWR VPWR cpu_ack_o sky130_fd_sc_hd__buf_2
X_1500_ _2875_/Q _1500_/B VGND VGND VPWR VPWR _1500_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1431_ _1431_/A VGND VGND VPWR VPWR _1444_/A sky130_fd_sc_hd__buf_2
XANTENNA__1781__A _1853_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1362_ _1362_/A _1362_/B _1362_/C VGND VGND VPWR VPWR _1362_/Y sky130_fd_sc_hd__nand3_1
X_1293_ _1355_/A VGND VGND VPWR VPWR _1367_/B sky130_fd_sc_hd__buf_2
XFILLER_49_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2098__A0 _2739_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2762__D _2762_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2117__A _2117_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2816_ _2816_/CLK _2816_/D VGND VGND VPWR VPWR _2816_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1956__A _1971_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2022__B1 _2021_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2747_ _2768_/CLK _2747_/D VGND VGND VPWR VPWR _2747_/Q sky130_fd_sc_hd__dfxtp_1
X_2678_ _2901_/CLK _2678_/D VGND VGND VPWR VPWR _2678_/Q sky130_fd_sc_hd__dfxtp_1
X_1629_ _1599_/X _1612_/X _2681_/Q VGND VGND VPWR VPWR _2175_/B sky130_fd_sc_hd__o21ai_1
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2938__CLK _2946_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input3_A cpu_adr_i[10] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2937__D _2937_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2089__B1 _2088_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1836__A0 _2750_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1300__A2 _1437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2672__D _2672_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2106__A2_N _1914_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2027__A _2027_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1992__A2_N _1933_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2013__A0 _2725_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2564__A1 _2868_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input59_A cpu_dat_i[31] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1772__C1 _1633_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1524__C1 _1311_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2847__D _2847_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1827__A0 _2339_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1980_ _1980_/A _2599_/A VGND VGND VPWR VPWR _1980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2601_ _2601_/A _2605_/B VGND VGND VPWR VPWR _2896_/D sky130_fd_sc_hd__nor2_1
XANTENNA__2004__B1 _2003_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2555__A1 _1412_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2532_ _2850_/Q _2519_/X _1801_/X _2531_/X VGND VGND VPWR VPWR _2850_/D sky130_fd_sc_hd__o211a_1
XFILLER_6_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2463_ _1748_/X _1751_/Y _2456_/X _2451_/X VGND VGND VPWR VPWR _2804_/D sky130_fd_sc_hd__o211a_1
X_2394_ input22/X _1785_/S _2393_/X _2365_/Y VGND VGND VPWR VPWR _2772_/D sky130_fd_sc_hd__a211o_1
X_1414_ _1414_/A _1429_/A _1414_/C _1414_/D VGND VGND VPWR VPWR _1414_/Y sky130_fd_sc_hd__nand4_1
XANTENNA__2400__A _2400_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1942__C _2258_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1345_ _1307_/X _1308_/X _2761_/Q VGND VGND VPWR VPWR _1345_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__2757__D _2757_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2491__B1 _1949_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1597__A2 _1559_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1349__A2 _1308_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2760__CLK _2764_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1754__C1 _1699_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_CLK clkbuf_1_0_0_CLK/X VGND VGND VPWR VPWR _2776_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2310__A _2320_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1506__C1 _2552_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2667__D _2667_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1809__A0 _2746_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2482__B1 _2128_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1299__C _2383_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2234__B1 _1519_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2204__B _2216_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_16_CLK_A clkbuf_1_1_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output165_A _1912_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1760__A2 _1712_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2220__A _2220_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_11_CLK clkbuf_1_1_0_CLK/X VGND VGND VPWR VPWR _2839_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_38_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2473__B1 _2231_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1963_ _2027_/A VGND VGND VPWR VPWR _2013_/S sky130_fd_sc_hd__clkbuf_2
X_1894_ _1900_/A _2942_/Q VGND VGND VPWR VPWR _1895_/A sky130_fd_sc_hd__and2_1
XANTENNA__1579__A2 _1578_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1937__C _2254_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2783__CLK _2816_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2114__B _2114_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1822__A2_N _1792_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1736__C1 _1710_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2515_ _2838_/Q _2506_/X _2067_/X _2514_/X VGND VGND VPWR VPWR _2838_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1751__A2 _1750_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2446_ _1690_/X _1694_/Y _2436_/X _2431_/X VGND VGND VPWR VPWR _2796_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1391__D _1447_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1503__A2 _1488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2377_ _2382_/A _2377_/B _2377_/C _2382_/D VGND VGND VPWR VPWR _2762_/D sky130_fd_sc_hd__nand4_1
XFILLER_56_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1328_ _2873_/Q _1324_/X _1327_/Y VGND VGND VPWR VPWR _1341_/A sky130_fd_sc_hd__o21ai_1
XFILLER_37_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2464__B1 _1753_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2008__C _2282_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2305__A _2352_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2024__B _2607_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1727__C1 _1705_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1742__A2 _1682_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2455__B1 _2454_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_CLK clkbuf_leaf_0_CLK/A VGND VGND VPWR VPWR _2880_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2860__D _2860_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2215__A _2215_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1476__D _1803_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1718__C1 _1699_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2300_ _2324_/A VGND VGND VPWR VPWR _2320_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1733__A2 _1732_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2231_ _2231_/A VGND VGND VPWR VPWR _2577_/A sky130_fd_sc_hd__clkbuf_4
X_2162_ _1577_/Y _1578_/Y _2156_/X VGND VGND VPWR VPWR _2674_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__1497__A1 _1367_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2093_ _2738_/Q input54/X _2093_/S VGND VGND VPWR VPWR _2315_/B sky130_fd_sc_hd__mux2_1
XFILLER_53_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2109__B _2109_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2446__B1 _2436_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2770__D _2770_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1946_ _2076_/A VGND VGND VPWR VPWR _2117_/A sky130_fd_sc_hd__clkbuf_4
X_1877_ _1877_/A VGND VGND VPWR VPWR _1877_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1972__A2 _1969_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2062__A1_N _2907_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1724__A2 _1663_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2679__CLK _2816_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2429_ _2412_/X _2177_/A _1625_/X VGND VGND VPWR VPWR _2429_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__2945__D _2945_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2437__B1 _2436_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1660__A1 _2185_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2680__D _2680_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2035__A _2035_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1874__A _1878_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1412__A1 _1379_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1715__A2 _1714_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input41_A cpu_dat_i[15] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2855__D _2855_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output128_A _1757_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1800_ _2745_/Q input13/X _1970_/S VGND VGND VPWR VPWR _2332_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2780_ _2816_/CLK _2780_/D VGND VGND VPWR VPWR _2780_/Q sky130_fd_sc_hd__dfxtp_1
X_1731_ _1672_/X _1685_/X _2695_/Q VGND VGND VPWR VPWR _2207_/B sky130_fd_sc_hd__o21ai_1
XFILLER_11_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1784__A _2113_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2599__B _2605_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1662_ _1635_/X _1617_/X _2792_/Q VGND VGND VPWR VPWR _1662_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2821__CLK _2920_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2272__C_N _2257_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1593_ _1632_/A VGND VGND VPWR VPWR _1593_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1706__A2 _1703_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1283__A_N _2777_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2214_ _1749_/Y _1750_/Y _2201_/X VGND VGND VPWR VPWR _2698_/D sky130_fd_sc_hd__a21oi_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2131__A2 _2649_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2765__D _2765_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2145_ _2235_/A VGND VGND VPWR VPWR _2526_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2076_ _2076_/A VGND VGND VPWR VPWR _2102_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2419__B1 _2418_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1959__A _1980_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_62_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1642__A1 _1639_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1929_ _1971_/A _2128_/B _2252_/B VGND VGND VPWR VPWR _1929_/X sky130_fd_sc_hd__or3_2
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2021__C _2286_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2658__B1 _2650_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2122__A2 _1853_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2675__D _2675_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1869__A _1902_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input89_A spi_dat_i[23] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2844__CLK _2881_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1397__B1 _1396_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2212__B _2216_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_1_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2361__A2 _2358_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1321__B1 _2861_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1779__A _1859_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2901_ _2901_/CLK _2901_/D VGND VGND VPWR VPWR _2901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2832_ _2834_/CLK _2832_/D VGND VGND VPWR VPWR _2832_/Q sky130_fd_sc_hd__dfxtp_1
X_2763_ _2768_/CLK _2763_/D VGND VGND VPWR VPWR _2763_/Q sky130_fd_sc_hd__dfxtp_1
X_1714_ _1711_/Y _1713_/Y _1679_/X VGND VGND VPWR VPWR _1714_/Y sky130_fd_sc_hd__a21oi_1
X_2694_ _2703_/CLK _2694_/D VGND VGND VPWR VPWR _2694_/Q sky130_fd_sc_hd__dfxtp_1
X_1645_ _1717_/A VGND VGND VPWR VPWR _1645_/X sky130_fd_sc_hd__buf_4
X_1576_ _1723_/A VGND VGND VPWR VPWR _1576_/X sky130_fd_sc_hd__buf_2
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1560__B1 _2779_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2717__CLK _2745_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1863__A1 _1859_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2128_ _2128_/A _2128_/B _2245_/A VGND VGND VPWR VPWR _2128_/X sky130_fd_sc_hd__or3_1
XFILLER_54_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2059_ _2732_/Q input48/X _2093_/S VGND VGND VPWR VPWR _2301_/B sky130_fd_sc_hd__mux2_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1689__A _1689_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2867__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1615__A1 _1610_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2040__A1 input44/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2313__A _2313_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1855__C _2350_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2032__B _2609_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1854__A1 input33/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1599__A _1692_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2207__B _2207_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output195_A _2107_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2223__A _2223_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2031__B2 _2030_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput109 _1557_/X VGND VGND VPWR VPWR cpu_dat_o[0] sky130_fd_sc_hd__buf_2
XANTENNA__1790__B1 _1789_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1430_ _1370_/A _1454_/B _1454_/C _1454_/D VGND VGND VPWR VPWR _1430_/Y sky130_fd_sc_hd__nand4b_1
X_1361_ _1296_/X _1297_/X _2763_/Q VGND VGND VPWR VPWR _1362_/C sky130_fd_sc_hd__o21ai_1
X_1292_ _2777_/Q _2776_/Q VGND VGND VPWR VPWR _1355_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2310__C_N _2305_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2098__A1 input55/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1302__A _2777_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2117__B _2626_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1956__B _2008_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2815_ _2925_/CLK _2815_/D VGND VGND VPWR VPWR _2815_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2022__A1 _2831_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2746_ _2925_/CLK _2746_/D VGND VGND VPWR VPWR _2746_/Q sky130_fd_sc_hd__dfxtp_1
X_2677_ _2816_/CLK _2677_/D VGND VGND VPWR VPWR _2677_/Q sky130_fd_sc_hd__dfxtp_1
X_1628_ _1561_/X _1582_/X _1626_/X _1627_/X _1628_/D1 VGND VGND VPWR VPWR _2175_/A
+ sky130_fd_sc_hd__o2111ai_4
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1559_ _1682_/A VGND VGND VPWR VPWR _1559_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2089__A1 _2842_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1836__A1 input30/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2308__A _2308_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2013__A1 input40/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2564__A2 _2540_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1882__A _1882_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1772__B1 _1632_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1524__B1 _1300_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1827__A1 _2853_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2483__C_N _2352_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2863__D _2863_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output208_A _2131_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output110_A _1643_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2600_ _2600_/A _2604_/B VGND VGND VPWR VPWR _2895_/D sky130_fd_sc_hd__nand2_1
XANTENNA__2004__A1 _2828_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2531_ _2531_/A VGND VGND VPWR VPWR _2531_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2555__A2 _1415_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1792__A _2064_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1763__B1 _2807_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2462_ _2447_/X _2448_/X _2461_/Y VGND VGND VPWR VPWR _2803_/D sky130_fd_sc_hd__o21ai_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1413_ input6/X VGND VGND VPWR VPWR _1414_/A sky130_fd_sc_hd__inv_2
X_2393_ _2395_/A _2395_/B _2395_/D _2772_/Q VGND VGND VPWR VPWR _2393_/X sky130_fd_sc_hd__o31a_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1344_ _1344_/A VGND VGND VPWR VPWR _1344_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__2773__D _2773_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2128__A _2128_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2491__A1 _2820_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2228__D1 _1572_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2905__CLK _2915_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2729_ _2834_/CLK _2729_/D VGND VGND VPWR VPWR _2729_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1754__B1 _1698_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2310__B _2310_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1506__B1 _1502_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2683__D _2683_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1809__A1 input24/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2038__A _2044_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2482__A1 _2814_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input106_A spi_err_i VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1877__A _1877_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2234__A1 _2706_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_42_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2234__B2 _2811_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input71_A cpu_stb_i VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1745__B1 _2697_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2501__A _2531_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output158_A _1899_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2220__B _2224_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2858__D _2858_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2170__B1 _2156_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2473__A1 _2395_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1681__C1 _1668_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2928__CLK _2930_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1962_ _2114_/A VGND VGND VPWR VPWR _2014_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1893_ _1893_/A VGND VGND VPWR VPWR _1893_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1984__A0 _2720_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2114__C _2325_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1736__B1 _1709_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2514_ _2531_/A VGND VGND VPWR VPWR _2514_/X sky130_fd_sc_hd__clkbuf_4
X_2445_ _2427_/X _2428_/X _2444_/Y VGND VGND VPWR VPWR _2795_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__2768__D _2768_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2376_ _2376_/A VGND VGND VPWR VPWR _2761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1327_ _2386_/B _2386_/C _1335_/C VGND VGND VPWR VPWR _1327_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__2464__A1 _2453_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1727__B1 _1704_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2321__A _2321_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2678__D _2678_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1944__A2_N _2573_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2455__A1 _2447_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1400__A _1400_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2215__B _2215_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1415__C1 _1362_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1966__B1 _1965_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1718__B1 _1698_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2231__A _2231_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _2415_/A VGND VGND VPWR VPWR _2231_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_39_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2161_ _2161_/A VGND VGND VPWR VPWR _2673_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1497__A2 _1457_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2092_ _2092_/A VGND VGND VPWR VPWR _2251_/A sky130_fd_sc_hd__buf_2
XFILLER_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2446__A1 _1690_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2109__C _2322_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2750__CLK _2873_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1310__A _1350_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1945_ _1945_/A _2592_/A VGND VGND VPWR VPWR _1945_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1957__B1 _1956_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1876_ _1878_/A _2934_/Q VGND VGND VPWR VPWR _1877_/A sky130_fd_sc_hd__and2_1
XFILLER_0_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1980__A _1980_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2134__B1 _1789_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2428_ _2448_/A VGND VGND VPWR VPWR _2428_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2359_ _2526_/A VGND VGND VPWR VPWR _2665_/C sky130_fd_sc_hd__buf_2
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_15_CLK_A clkbuf_1_1_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2437__A1 _1650_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1660__A2 _2185_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2316__A _2316_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2035__B _2072_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1948__A0 _2715_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1874__B _2933_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1412__A2 _1380_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2373__B1 _1345_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1890__A _1890_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2125__B1 _1789_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2773__CLK _2776_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input34_A cpu_cyc_i VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2871__D _2871_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2226__A _2537_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1939__B1 _1916_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1730_ _1717_/X _1729_/X _1698_/X _1699_/X input89/X VGND VGND VPWR VPWR _2207_/A
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1661_ _1656_/X _1660_/Y _1632_/X _1633_/X VGND VGND VPWR VPWR _1661_/X sky130_fd_sc_hd__o211a_1
XFILLER_4_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1592_ _1739_/A VGND VGND VPWR VPWR _1632_/A sky130_fd_sc_hd__buf_2
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2116__B1 _1916_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2213_ _2213_/A VGND VGND VPWR VPWR _2697_/D sky130_fd_sc_hd__clkbuf_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1305__A _2366_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2144_ input1/X VGND VGND VPWR VPWR _2235_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2075_ _2075_/A _2616_/A VGND VGND VPWR VPWR _2075_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2419__A1 _2408_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1959__B _2595_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2136__A _2649_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_50_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1642__A2 _1641_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2781__D _2781_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1975__A _2058_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1928_ _2712_/Q input46/X _1970_/S VGND VGND VPWR VPWR _2252_/B sky130_fd_sc_hd__mux2_1
X_1859_ _1859_/A VGND VGND VPWR VPWR _1859_/X sky130_fd_sc_hd__buf_2
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2796__CLK _2839_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2658__A1 _2941_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2691__D _2691_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2046__A _2046_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1885__A _1889_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1397__A1 _2865_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output140_A _1634_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2866__D _2866_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1321__A1 _1424_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2900_ _2915_/CLK _2900_/D VGND VGND VPWR VPWR _2900_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2669__CLK _2946_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2831_ _2901_/CLK _2831_/D VGND VGND VPWR VPWR _2831_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1795__A _2046_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2762_ _2764_/CLK _2762_/D VGND VGND VPWR VPWR _2762_/Q sky130_fd_sc_hd__dfxtp_1
X_1713_ _1692_/X _1712_/X _2692_/Q VGND VGND VPWR VPWR _1713_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2693_ _2703_/CLK _2693_/D VGND VGND VPWR VPWR _2693_/Q sky130_fd_sc_hd__dfxtp_1
X_1644_ _1624_/X _1609_/X _2789_/Q VGND VGND VPWR VPWR _1644_/X sky130_fd_sc_hd__o21a_1
X_1575_ _1517_/X _1519_/X _2780_/Q VGND VGND VPWR VPWR _1575_/X sky130_fd_sc_hd__o21a_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1560__A1 _1558_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2776__D _2776_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1863__A2 _1853_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2127_ _2709_/Q input69/X _2127_/S VGND VGND VPWR VPWR _2245_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2058_ _2058_/A VGND VGND VPWR VPWR _2058_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1615__A2 _1614_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2576__B1 _1311_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2313__B _2332_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2686__D _2686_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2811__CLK _2881_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2262__C_N _2257_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1819__S _2108_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2567__B1 _2552_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output188_A _2070_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2223__B _2223_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1790__A1 _2649_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1790__B2 _2919_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1360_ _1414_/C _1414_/D _1360_/C _1367_/B VGND VGND VPWR VPWR _1362_/B sky130_fd_sc_hd__nand4_2
XFILLER_49_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1291_ _1291_/A VGND VGND VPWR VPWR _1354_/A sky130_fd_sc_hd__buf_2
XFILLER_64_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2814_ _2929_/CLK _2814_/D VGND VGND VPWR VPWR _2814_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1956__C _2262_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2022__A2 _1969_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2745_ _2745_/CLK _2745_/D VGND VGND VPWR VPWR _2745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2676_ _2816_/CLK _2676_/D VGND VGND VPWR VPWR _2676_/Q sky130_fd_sc_hd__dfxtp_1
X_1627_ _1699_/A VGND VGND VPWR VPWR _1627_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_28_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1558_ _1696_/A VGND VGND VPWR VPWR _1558_/X sky130_fd_sc_hd__clkbuf_2
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1489_ _1445_/A _1488_/X _2864_/Q VGND VGND VPWR VPWR _1489_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_28_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2834__CLK _2834_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2089__A2 _1814_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2494__C1 _2488_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2308__B _2308_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2324__A _2324_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1772__A1 _1768_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1524__A1 _2879_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2485__C1 _2525_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1403__A _2671_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1460__B1 _1459_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2707__CLK _2776_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2004__A2 _1961_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2530_ _2530_/A VGND VGND VPWR VPWR _2849_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2461_ _2453_/X _2212_/A _1742_/X VGND VGND VPWR VPWR _2461_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__1763__A1 _1707_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1412_ _1379_/X _1380_/A _2862_/Q VGND VGND VPWR VPWR _1412_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2857__CLK _2925_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2392_ _2392_/A VGND VGND VPWR VPWR _2771_/D sky130_fd_sc_hd__clkbuf_1
X_1343_ _1343_/A VGND VGND VPWR VPWR _1343_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_58_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2128__B _2128_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2491__A2 _2475_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2228__C1 _2386_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2144__A input1/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1983__A _2047_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2728_ _2834_/CLK _2728_/D VGND VGND VPWR VPWR _2728_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1754__A1 _1717_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2659_ _2665_/A _2942_/Q _2665_/C VGND VGND VPWR VPWR _2660_/A sky130_fd_sc_hd__and3_1
XANTENNA__1506__A1 _1500_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2319__A _2319_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2038__B _2610_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2482__A2 _2475_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1690__B1 _2796_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2234__A2 _2529_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2054__A _2078_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1893__A _1893_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1745__A1 _1744_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input64_A cpu_dat_i[7] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2170__A1 _1604_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2874__D _2874_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2229__A _2235_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2473__A2 _2395_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1681__B1 _1667_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1961_ _2324_/A VGND VGND VPWR VPWR _1961_/X sky130_fd_sc_hd__buf_2
X_1892_ _1900_/A _2941_/Q VGND VGND VPWR VPWR _1893_/A sky130_fd_sc_hd__and2_1
XANTENNA__1984__A1 input66/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1736__A1 _1723_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2513_ _2513_/A _2521_/B VGND VGND VPWR VPWR _2837_/D sky130_fd_sc_hd__nand2_1
XANTENNA__1308__A _1372_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2444_ _2433_/X _2194_/A _1683_/X VGND VGND VPWR VPWR _2444_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_25_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2375_ _2375_/A _2391_/B _2399_/C VGND VGND VPWR VPWR _2376_/A sky130_fd_sc_hd__and3_1
XFILLER_56_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1326_ _1296_/X _1297_/X _2768_/Q VGND VGND VPWR VPWR _2386_/C sky130_fd_sc_hd__o21ai_2
XFILLER_57_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2784__D _2784_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2139__A _2580_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2464__A2 _2216_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2602__A _2602_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1727__A1 _1722_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2694__D _2694_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2049__A _2094_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2455__A2 _2448_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1888__A _1888_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1415__B1 _1414_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1966__A1 _2822_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1827__S _2124_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1718__A1 _1717_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2869__D _2869_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output170_A _1848_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2160_ _2160_/A _2172_/B VGND VGND VPWR VPWR _2161_/A sky130_fd_sc_hd__or2_1
XANTENNA__1351__C1 _1362_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2091_ _2102_/A _2621_/A VGND VGND VPWR VPWR _2091_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1654__B1 _1606_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1798__A _2047_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2446__A2 _1694_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1944_ _2889_/Q _2573_/A _1927_/X _2490_/A VGND VGND VPWR VPWR _2592_/A sky130_fd_sc_hd__a2bb2o_2
XANTENNA__1957__A1 _2821_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1875_ _1875_/A VGND VGND VPWR VPWR _1875_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__2779__D _2779_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1980__B _2599_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2427_ _2447_/A VGND VGND VPWR VPWR _2427_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2134__A1 _1853_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2134__B2 _2885_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2358_ _2358_/A VGND VGND VPWR VPWR _2358_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1309_ _1307_/X _1308_/X _2774_/Q VGND VGND VPWR VPWR _1309_/Y sky130_fd_sc_hd__o21ai_2
X_2289_ _2289_/A _2308_/B _2289_/C VGND VGND VPWR VPWR _2290_/A sky130_fd_sc_hd__and3_1
XFILLER_25_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2437__A2 _1654_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1948__A1 input61/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2035__C _2291_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2332__A _2332_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2689__D _2689_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2373__A1 _1344_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2125__A1 _1853_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2918__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2125__B2 _2883_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input27_A cpu_adr_i[3] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1411__A _1411_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1636__B1 _2788_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1939__B2 _1938_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2061__B1 _2060_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1660_ _2185_/A _2185_/B _1630_/X VGND VGND VPWR VPWR _1660_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__2242__A _2242_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1591_ _1589_/Y _1590_/Y _1549_/X VGND VGND VPWR VPWR _1591_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_7_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2116__B2 _2525_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2212_ _2212_/A _2216_/B VGND VGND VPWR VPWR _2213_/A sky130_fd_sc_hd__or2_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2143_ _2652_/A VGND VGND VPWR VPWR _2647_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__1305__B _1422_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2074_ _2909_/Q _2018_/X _2058_/X _2516_/A VGND VGND VPWR VPWR _2616_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__2419__A2 _2410_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1927_ _2058_/A VGND VGND VPWR VPWR _1927_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1958__A2_N _1953_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1858_ _1830_/X _1853_/X _2637_/A VGND VGND VPWR VPWR _1858_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__2152__A _2949_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1789_ _1789_/A VGND VGND VPWR VPWR _1789_/X sky130_fd_sc_hd__buf_2
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2658__A2 _2649_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1866__B1 _1865_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2327__A _2327_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1618__B1 _2786_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1885__B _2938_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2043__B1 _2039_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2090__A2_N _2064_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1397__A2 _1287_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_5_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2740__CLK _2834_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1406__A _1509_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_945 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2890__CLK _2917_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1857__B1 _1840_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output133_A _1777_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1321__A2 _1380_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2882__D _2882_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2237__A _2374_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2043__A2_N _2000_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2830_ _2847_/CLK _2830_/D VGND VGND VPWR VPWR _2830_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2034__A0 _2728_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2761_ _2768_/CLK _2761_/D VGND VGND VPWR VPWR _2761_/Q sky130_fd_sc_hd__dfxtp_1
X_2692_ _2703_/CLK _2692_/D VGND VGND VPWR VPWR _2692_/Q sky130_fd_sc_hd__dfxtp_1
X_1712_ _1712_/A VGND VGND VPWR VPWR _1712_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2534__C_N _2352_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_14_CLK_A clkbuf_1_1_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1643_ _1636_/X _1642_/Y _1632_/X _1633_/X VGND VGND VPWR VPWR _1643_/X sky130_fd_sc_hd__o211a_1
X_1574_ _1560_/X _1573_/Y _1473_/X _1556_/X VGND VGND VPWR VPWR _1574_/X sky130_fd_sc_hd__o211a_1
XFILLER_59_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1316__A _1390_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1560__A2 _1559_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_39_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1848__B1 _2635_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2126_ _1859_/X _1853_/X _2585_/B VGND VGND VPWR VPWR _2126_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__2147__A _2647_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2057_ _2075_/A _2613_/A VGND VGND VPWR VPWR _2057_/Y sky130_fd_sc_hd__nor2_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2792__D _2792_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2763__CLK _2768_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2576__A1 _2879_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2313__C _2313_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2610__A _2610_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2121__A1_N _2882_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1839__B1 _2634_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2057__A _2075_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1896__A _1900_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input94_A spi_dat_i[28] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2016__B1 _1975_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2567__A1 _1493_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1790__A2 _2529_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2877__D _2877_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1290_ _1353_/A VGND VGND VPWR VPWR _1414_/C sky130_fd_sc_hd__buf_2
XFILLER_49_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2786__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2813_ _2925_/CLK _2813_/D VGND VGND VPWR VPWR _2813_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2007__A0 _2724_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2744_ _2873_/CLK _2744_/D VGND VGND VPWR VPWR _2744_/Q sky130_fd_sc_hd__dfxtp_1
X_2675_ _2816_/CLK _2675_/D VGND VGND VPWR VPWR _2675_/Q sky130_fd_sc_hd__dfxtp_1
X_1626_ _1698_/A VGND VGND VPWR VPWR _1626_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_28_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1557_ _1520_/X _1550_/Y _1473_/X _1556_/X VGND VGND VPWR VPWR _1557_/X sky130_fd_sc_hd__o211a_1
XANTENNA__2787__D _2787_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1488_ _1488_/A VGND VGND VPWR VPWR _1488_/X sky130_fd_sc_hd__clkbuf_2
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1480__S _2243_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2494__B1 _1965_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2109_ _2109_/A _2109_/B _2322_/A VGND VGND VPWR VPWR _2109_/X sky130_fd_sc_hd__or3_2
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2308__C _2313_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2605__A _2605_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1757__C1 _1740_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1772__A2 _1771_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2340__A _2340_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2697__D _2697_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1524__A2 _2092_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2485__B1 _1922_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1403__B _2706_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1460__A1 _2862_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2250__A _2250_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_14_CLK clkbuf_1_1_0_CLK/X VGND VGND VPWR VPWR _2840_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1763__A2 _1689_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2460_ _1734_/X _1738_/Y _2456_/X _2451_/X VGND VGND VPWR VPWR _2802_/D sky130_fd_sc_hd__o211a_1
X_1411_ _1411_/A _1411_/B _1437_/A VGND VGND VPWR VPWR _1411_/Y sky130_fd_sc_hd__nand3_1
X_2391_ _2391_/A _2391_/B _2399_/C VGND VGND VPWR VPWR _2392_/A sky130_fd_sc_hd__and3_1
X_1342_ _1342_/A _1342_/B VGND VGND VPWR VPWR _1803_/A sky130_fd_sc_hd__nor2_4
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2476__B1 _2235_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1684__D1 input82/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2128__C _2245_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2228__B1 _1552_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2727_ _2834_/CLK _2727_/D VGND VGND VPWR VPWR _2727_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1754__A2 _1729_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1867__A1_N _2930_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2160__A _2160_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2658_ _2941_/Q _2649_/X _2650_/X VGND VGND VPWR VPWR _2941_/D sky130_fd_sc_hd__a21o_1
XANTENNA__2801__CLK _2809_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2589_ _2618_/A VGND VGND VPWR VPWR _2638_/A sky130_fd_sc_hd__buf_2
X_1609_ _1682_/A VGND VGND VPWR VPWR _1609_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2252__C_N _2227_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1506__A2 _1501_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input1_A RST_N VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2467__B1 _1763_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1805__A1_N _2920_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1690__A1 _1635_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2335__A _2335_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2054__B _2054_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2070__A _2075_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1745__A2 _1685_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input57_A cpu_dat_i[2] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_2_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2170__A2 _1605_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1414__A _1414_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2458__B1 _1728_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_3_CLK clkbuf_1_0_0_CLK/X VGND VGND VPWR VPWR _2929_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1681__A1 _1676_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2890__D _2890_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_33_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2245__A _2245_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1960_ _2092_/A VGND VGND VPWR VPWR _2324_/A sky130_fd_sc_hd__clkbuf_2
X_1891_ _1902_/A VGND VGND VPWR VPWR _1900_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_30_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2824__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1736__A2 _2533_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2394__C1 _2365_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2512_ _2836_/Q _2506_/X _2054_/X _2501_/X VGND VGND VPWR VPWR _2836_/D sky130_fd_sc_hd__o211a_1
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2443_ _1676_/X _1680_/Y _2436_/X _2431_/X VGND VGND VPWR VPWR _2794_/D sky130_fd_sc_hd__o211a_1
XFILLER_64_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2374_ _2374_/A VGND VGND VPWR VPWR _2399_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_25_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1325_ _1325_/A _1390_/A VGND VGND VPWR VPWR _2386_/B sky130_fd_sc_hd__nand2_4
XANTENNA__1324__A _1343_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2449__B1 _1697_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2155__A _2198_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1994__A _2058_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2602__B _2604_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_clkbuf_opt_3_0_CLK_A clkbuf_1_1_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1727__A2 _1726_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2049__B _2072_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2065__A _2065_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1415__A1 _2757_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2847__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1966__A2 _1961_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1718__A2 _1657_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1409__A _1409_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output163_A _1812_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2885__D _2885_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1351__B1 _1349_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2090_ _2912_/Q _2064_/X _2039_/X _2089_/Y VGND VGND VPWR VPWR _2621_/A sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1639__D1 input75/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_34_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1654__A1 _1652_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1943_ _2819_/Q _2474_/A _1942_/X VGND VGND VPWR VPWR _2490_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__1957__A2 _2474_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1874_ _1878_/A _2933_/Q VGND VGND VPWR VPWR _1875_/A sky130_fd_sc_hd__and2_1
XANTENNA__2367__C1 _2366_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1590__B1 _2676_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_9_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2426_ _1618_/X _1622_/Y _2416_/X _2405_/X VGND VGND VPWR VPWR _2786_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2134__A2 _2483_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2795__D _2795_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2357_ _2364_/A VGND VGND VPWR VPWR _2357_/X sky130_fd_sc_hd__clkbuf_4
X_2288_ _2312_/A VGND VGND VPWR VPWR _2308_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1308_ _1372_/A VGND VGND VPWR VPWR _1308_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2613__A _2613_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1928__S _1970_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2332__B _2332_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2373__A2 _1457_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1581__B1 _2781_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2125__A2 _2480_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1899__A _1899_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1636__A1 _1635_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1411__B _1411_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2061__A1 _2837_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2523__A _2523_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1590_ _2152_/B _1543_/X _2676_/Q VGND VGND VPWR VPWR _1590_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ _2211_/A _2211_/B VGND VGND VPWR VPWR _2212_/A sky130_fd_sc_hd__nand2_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2142_ _1528_/A _1528_/B _1692_/A _1859_/A VGND VGND VPWR VPWR _2652_/A sky130_fd_sc_hd__o22a_1
XANTENNA__1305__C _1354_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2073_ _2839_/Q _2033_/X _2072_/X VGND VGND VPWR VPWR _2516_/A sky130_fd_sc_hd__o21ai_1
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2433__A _2453_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1926_ _2233_/A VGND VGND VPWR VPWR _2573_/A sky130_fd_sc_hd__buf_2
X_1857_ _2928_/Q _1792_/X _1840_/X _1856_/Y VGND VGND VPWR VPWR _2637_/A sky130_fd_sc_hd__a2bb2o_1
XANTENNA__2152__B _2152_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1788_ _1803_/A _1788_/B _1803_/D VGND VGND VPWR VPWR _1789_/A sky130_fd_sc_hd__and3_2
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2409_ _2395_/B _2395_/D _2537_/A _2366_/B VGND VGND VPWR VPWR _2448_/A sky130_fd_sc_hd__o211a_4
XFILLER_57_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2692__CLK _2703_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1866__A1 _2860_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2512__C1 _2501_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2608__A _2650_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1512__A _1512_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2327__B _2332_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1618__A1 _1517_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2579__C1 _2527_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2043__B2 _2042_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2343__A _2343_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1554__B1 _2810_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1406__B _1406_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1857__B2 _1856_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2518__A _2518_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output126_A _1747_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1422__A _1422_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_1_1_0_CLK/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2034__A1 input43/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2760_ _2764_/CLK _2760_/D VGND VGND VPWR VPWR _2760_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2253__A _2253_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1711_ _1651_/X _1663_/X _1709_/X _1710_/X input86/X VGND VGND VPWR VPWR _1711_/Y
+ sky130_fd_sc_hd__o2111ai_2
X_2691_ _2839_/CLK _2691_/D VGND VGND VPWR VPWR _2691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1642_ _1639_/Y _1641_/Y _1606_/X VGND VGND VPWR VPWR _1642_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1545__B1 _1539_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1573_ _2158_/A _2158_/B _1572_/X VGND VGND VPWR VPWR _1573_/Y sky130_fd_sc_hd__a21oi_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1848__A1 _1830_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2125_ _1853_/A _2480_/B _1789_/A _2883_/Q VGND VGND VPWR VPWR _2585_/B sky130_fd_sc_hd__o22ai_2
XFILLER_27_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2428__A _2448_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2147__B _2668_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2056_ _2906_/Q _2000_/X _2039_/X _2055_/Y VGND VGND VPWR VPWR _2613_/A sky130_fd_sc_hd__a2bb2o_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1478__S _2047_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2908__CLK _2915_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2163__A _2163_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1909_ _1911_/A _2669_/Q VGND VGND VPWR VPWR _1910_/A sky130_fd_sc_hd__and2_1
XANTENNA__2576__A2 _2493_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2889_ _2920_/CLK _2889_/D VGND VGND VPWR VPWR _2889_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2610__B _2616_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1839__A1 _1830_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1941__S _1970_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2338__A _2338_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2057__B _2613_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_26_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1896__B _2943_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2016__B2 _2015_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input87_A spi_dat_i[21] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2567__A2 _1339_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1775__B1 _2703_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_12_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1417__A _2556_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2893__D _2893_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2248__A _2248_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2812_ _2929_/CLK _2812_/D VGND VGND VPWR VPWR _2812_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2007__A1 input39/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2743_ _2776_/CLK _2743_/D VGND VGND VPWR VPWR _2743_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1766__B1 _1549_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2674_ _2920_/CLK _2674_/D VGND VGND VPWR VPWR _2674_/Q sky130_fd_sc_hd__dfxtp_1
X_1625_ _1624_/X _1609_/X _2787_/Q VGND VGND VPWR VPWR _1625_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1327__A _2386_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1556_ _1740_/A VGND VGND VPWR VPWR _1556_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1487_ _2389_/A _1436_/A _1452_/X _1377_/Y _1500_/B VGND VGND VPWR VPWR _1487_/X
+ sky130_fd_sc_hd__o311a_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2158__A _2158_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2494__A1 _2822_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2108_ _2741_/Q input58/X _2108_/S VGND VGND VPWR VPWR _2322_/A sky130_fd_sc_hd__mux2_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2039_ _2039_/A VGND VGND VPWR VPWR _2039_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_36_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2730__CLK _2834_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2605__B _2605_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2880__CLK _2880_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1936__S _2132_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1757__B1 _1739_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2621__A _2621_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2485__A1 _2816_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_13_CLK_A clkbuf_opt_3_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2007__S _2034_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1460__A2 _1523_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_14_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output193_A _2097_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1748__B1 _2804_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2531__A _2531_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_10_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2888__D _2888_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1410_ _1451_/A _1452_/A _2771_/Q VGND VGND VPWR VPWR _1411_/B sky130_fd_sc_hd__o21ai_1
X_2390_ _2395_/B _1409_/A _1452_/X _1455_/B VGND VGND VPWR VPWR _2391_/A sky130_fd_sc_hd__o31a_1
X_1341_ _1341_/A _1341_/B _1341_/C _1341_/D VGND VGND VPWR VPWR _1342_/B sky130_fd_sc_hd__nand4_4
XFILLER_64_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2753__CLK _2764_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2476__A1 _1342_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1684__C1 _1627_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2228__A1 _1551_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_17_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1987__B1 _1927_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1834__A2_N _1792_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2726_ _2834_/CLK _2726_/D VGND VGND VPWR VPWR _2726_/Q sky130_fd_sc_hd__dfxtp_1
X_2657_ _2657_/A VGND VGND VPWR VPWR _2940_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__2160__B _2172_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2798__D _2798_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1608_ _1603_/X _1607_/Y _1593_/X _1595_/X VGND VGND VPWR VPWR _1608_/X sky130_fd_sc_hd__o211a_1
X_2588_ _2588_/A _2593_/B VGND VGND VPWR VPWR _2886_/D sky130_fd_sc_hd__nor2_1
XFILLER_59_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1539_ _1539_/A VGND VGND VPWR VPWR _1744_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2467__A1 _2453_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1675__C1 _1668_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2616__A _2616_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_36_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1690__A2 _1689_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1978__B1 _1977_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2054__C _2298_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2351__A _2351_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2070__B _2615_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2776__CLK _2776_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2458__A1 _2453_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1414__B _1429_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output206_A _2122_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1681__A2 _1680_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2526__A _2526_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2245__B _2260_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1890_ _1890_/A VGND VGND VPWR VPWR _1890_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2261__A _2261_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2511_ _2511_/A _2521_/B VGND VGND VPWR VPWR _2835_/D sky130_fd_sc_hd__nand2_1
XANTENNA__2394__B1 _2393_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2442_ _2427_/X _2428_/X _2441_/Y VGND VGND VPWR VPWR _2793_/D sky130_fd_sc_hd__o21ai_1
X_2373_ _1344_/Y _1457_/X _1345_/Y VGND VGND VPWR VPWR _2375_/A sky130_fd_sc_hd__o21ai_1
XFILLER_25_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1324_ _1343_/A VGND VGND VPWR VPWR _1324_/X sky130_fd_sc_hd__buf_2
XANTENNA__2449__A1 _2433_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_25_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2436__A _2558_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_944 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2074__A1_N _2909_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2171__A _2171_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_3_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2709_ _2776_/CLK _2709_/D VGND VGND VPWR VPWR _2709_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2799__CLK _2809_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1515__A _1515_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2049__C _2296_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2346__A _2346_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input104_A spi_dat_i[8] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1415__A2 _1428_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2081__A _2102_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1409__B _1409_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output156_A _1895_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2020__S _2034_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1425__A _1445_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1351__A1 _1348_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1639__C1 _1638_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1654__A2 _1653_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2256__A input1/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1942_ _1971_/A _2128_/B _2258_/B VGND VGND VPWR VPWR _1942_/X sky130_fd_sc_hd__or3_2
X_1873_ _1873_/A VGND VGND VPWR VPWR _1873_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2941__CLK _2946_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2367__B1 _2365_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1590__A1 _2152_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2425_ _2408_/X _2410_/X _2424_/Y VGND VGND VPWR VPWR _2785_/D sky130_fd_sc_hd__o21ai_1
XFILLER_9_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1335__A _2398_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2356_ _2356_/A VGND VGND VPWR VPWR _2755_/D sky130_fd_sc_hd__clkbuf_1
X_1307_ _1371_/A VGND VGND VPWR VPWR _1307_/X sky130_fd_sc_hd__clkbuf_4
X_2287_ _2287_/A VGND VGND VPWR VPWR _2726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2613__B _2617_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2332__C _2337_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1566__D1 input85/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1581__A1 _1558_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2814__CLK _2929_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_56_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2076__A _2076_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1411__C _1437_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1636__A2 _1617_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2061__A2 _2033_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2523__B _2525_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1854__S _2127_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2896__D _2896_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _1736_/Y _1737_/Y _2201_/X VGND VGND VPWR VPWR _2696_/D sky130_fd_sc_hd__a21oi_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2141_ _2667_/Q _2136_/X _2140_/X VGND VGND VPWR VPWR _2667_/D sky130_fd_sc_hd__a21o_1
XANTENNA__1305__D _1353_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2072_ _2094_/A _2072_/B _2306_/B VGND VGND VPWR VPWR _2072_/X sky130_fd_sc_hd__or3_1
XANTENNA__1493__B1_N _2871_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1925_ _1945_/A _2588_/A VGND VGND VPWR VPWR _1925_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2152__C _2401_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1856_ _2858_/Q _1841_/X _1855_/X VGND VGND VPWR VPWR _1856_/Y sky130_fd_sc_hd__o21ai_1
X_1787_ _2330_/B _2849_/Q _2374_/A VGND VGND VPWR VPWR _2529_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2837__CLK _2839_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2408_ _2447_/A VGND VGND VPWR VPWR _2408_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1866__A2 _1841_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2512__B1 _2054_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2339_ _2344_/A _2339_/B _2329_/X VGND VGND VPWR VPWR _2340_/A sky130_fd_sc_hd__or3b_1
XFILLER_29_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1512__B _1512_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2327__C _2337_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1618__A2 _1617_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2624__A _2624_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_41_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2579__B1 _2554_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1554__A1 _1515_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1406__C _1509_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input32_A cpu_adr_i[8] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1711__D1 input86/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2518__B _2521_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1422__B _1454_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output119_A _1706_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_44_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2534__A _2548_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1849__S _1860_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1710_ _1710_/A VGND VGND VPWR VPWR _1710_/X sky130_fd_sc_hd__buf_2
X_2690_ _2839_/CLK _2690_/D VGND VGND VPWR VPWR _2690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1641_ _1620_/X _1640_/X _2682_/Q VGND VGND VPWR VPWR _1641_/Y sky130_fd_sc_hd__o21ai_1
X_1572_ _1630_/A VGND VGND VPWR VPWR _1572_/X sky130_fd_sc_hd__buf_2
XANTENNA__1545__A1 _1778_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1848__A2 _1824_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2124_ _2241_/B _2813_/Q _2124_/S VGND VGND VPWR VPWR _2480_/B sky130_fd_sc_hd__mux2_1
XFILLER_26_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2147__C _2401_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2055_ _2836_/Q _2025_/X _2054_/X VGND VGND VPWR VPWR _2055_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_63_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1481__B1 _2918_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1769__D1 input97/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2163__B _2163_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1908_ _1908_/A VGND VGND VPWR VPWR _1908_/X sky130_fd_sc_hd__clkbuf_1
X_2888_ _2917_/CLK _2888_/D VGND VGND VPWR VPWR _2888_/Q sky130_fd_sc_hd__dfxtp_1
X_1839_ _1830_/X _1824_/X _2634_/B VGND VGND VPWR VPWR _1839_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_2_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2619__A _2619_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1839__A2 _1824_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1523__A _1523_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2354__A _2354_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1775__A1 _1744_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1417__B _2560_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_49_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2529__A _2529_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1433__A _1510_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2264__A _2312_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2811_ _2881_/CLK _2811_/D VGND VGND VPWR VPWR _2811_/Q sky130_fd_sc_hd__dfxtp_1
X_2742_ _2847_/CLK _2742_/D VGND VGND VPWR VPWR _2742_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2682__CLK _2901_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1766__A1 _2219_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2673_ _2816_/CLK _2673_/D VGND VGND VPWR VPWR _2673_/Q sky130_fd_sc_hd__dfxtp_1
X_1624_ _1696_/A VGND VGND VPWR VPWR _1624_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1555_ _1548_/A _1553_/Y _1554_/Y VGND VGND VPWR VPWR _1740_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__1327__B _2386_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_28_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1486_ _2870_/Q _1523_/A VGND VGND VPWR VPWR _1486_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2479__C1 _2525_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1343__A _1343_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2158__B _2158_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2494__A2 _2493_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2107_ _2117_/A _2624_/A VGND VGND VPWR VPWR _2107_/Y sky130_fd_sc_hd__nor2_4
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2038_ _2044_/A _2610_/A VGND VGND VPWR VPWR _2038_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1757__A1 _1753_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2621__B _2631_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1518__A _1616_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2113__S _2113_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_1_0_0_CLK clkbuf_0_CLK/X VGND VGND VPWR VPWR clkbuf_1_0_0_CLK/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2349__A _2349_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2485__A2 _2475_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_46_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1693__B1 _2690_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1748__A1 _1707_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output186_A _2057_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1428__A _1428_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1340_ _2871_/Q _1324_/X _1339_/Y VGND VGND VPWR VPWR _1341_/D sky130_fd_sc_hd__o21ai_1
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2259__A _2259_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2476__A2 _1342_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1684__B1 _1626_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2228__A2 _1482_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1987__B2 _2498_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_32_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2397__D1 _2386_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2725_ _2745_/CLK _2725_/D VGND VGND VPWR VPWR _2725_/Q sky130_fd_sc_hd__dfxtp_1
X_2656_ _2665_/A _2940_/Q _2665_/C VGND VGND VPWR VPWR _2657_/A sky130_fd_sc_hd__and3_1
X_1607_ _1604_/Y _1605_/Y _1606_/X VGND VGND VPWR VPWR _1607_/Y sky130_fd_sc_hd__a21oi_1
X_2587_ _2632_/A _2587_/B VGND VGND VPWR VPWR _2885_/D sky130_fd_sc_hd__nand2_1
X_1538_ input73/X _1465_/X _2705_/Q VGND VGND VPWR VPWR _1539_/A sky130_fd_sc_hd__o21bai_1
XFILLER_41_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2169__A _2169_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1469_ _2811_/Q VGND VGND VPWR VPWR _1469_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2467__A2 _2220_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1675__B1 _1667_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_43_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1801__A _1971_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2616__B _2616_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2108__S _2108_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1427__B1 _2867_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_51_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1978__A1 _2824_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_23_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__2632__A _2632_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1414__C _1414_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_58_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2458__A2 _2208_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1666__B1 _1606_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1418__B1 _2671_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1430__B _1454_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_15_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2245__C _2265_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2542__A _2548_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2379__D1 _2386_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2899__D _2899_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2510_ _2510_/A VGND VGND VPWR VPWR _2521_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__2394__A1 input22/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2441_ _2433_/X _2190_/A _1670_/X VGND VGND VPWR VPWR _2441_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_5_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2720__CLK _2745_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2372_ _2382_/A _2372_/B _2372_/C _2382_/D VGND VGND VPWR VPWR _2760_/D sky130_fd_sc_hd__nand4_1
XFILLER_57_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1323_ _2879_/Q _1287_/X _1300_/Y _1311_/Y _2552_/A VGND VGND VPWR VPWR _1342_/A
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2449__A2 _2199_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2870__CLK _2880_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2082__A0 _2736_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_20_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2171__B _2171_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2056__A2_N _2000_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2708_ _2873_/CLK _2708_/D VGND VGND VPWR VPWR _2708_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_12_CLK_A clkbuf_1_1_0_CLK/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2639_ _2639_/A _2639_/B VGND VGND VPWR VPWR _2930_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1648__B1 _1630_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1531__A _1531_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2346__B _2355_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2073__B1 _2072_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_24_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2362__A _2362_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_11_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2081__B _2617_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_8_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2743__CLK _2776_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_input62_A cpu_dat_i[5] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2893__CLK _2917_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA_output149_A _1882_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1351__A2 _1306_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1639__B1 _1637_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2537__A _2537_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1941_ _2714_/Q input60/X _1970_/S VGND VGND VPWR VPWR _2258_/B sky130_fd_sc_hd__mux2_1
X_1872_ _1878_/A _2932_/Q VGND VGND VPWR VPWR _1873_/A sky130_fd_sc_hd__and2_1
XANTENNA__1811__B1 _1789_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2272__A _2272_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_31_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2367__A1 _2758_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1616__A _1616_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1590__A2 _1543_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2424_ _2412_/X _2172_/A _1610_/X VGND VGND VPWR VPWR _2424_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2355_ _2355_/A _2355_/B _2370_/C VGND VGND VPWR VPWR _2356_/A sky130_fd_sc_hd__and3_1
XFILLER_9_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1335__B _2398_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1306_ _1306_/A VGND VGND VPWR VPWR _1457_/A sky130_fd_sc_hd__buf_4
X_2286_ _2296_/A _2286_/B _2281_/X VGND VGND VPWR VPWR _2287_/A sky130_fd_sc_hd__or3b_1
XFILLER_38_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2447__A _2447_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1973__A1_N _2893_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_52_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2055__B1 _2054_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2182__A _2182_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1802__B1 _1801_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2766__CLK _2768_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1566__C1 _1565_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1581__A2 _1559_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2357__A _2364_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_18_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2092__A _2092_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1557__C1 _1556_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1436__A _1436_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2140_ _2639_/B VGND VGND VPWR VPWR _2140_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2071_ _2734_/Q input50/X _2093_/S VGND VGND VPWR VPWR _2306_/B sky130_fd_sc_hd__mux2_1
XANTENNA__2267__A _2272_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_19_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2789__CLK _2847_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_35_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2037__B1 _1994_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1924_ _2886_/Q _1914_/X _1916_/X _1923_/Y VGND VGND VPWR VPWR _2588_/A sky130_fd_sc_hd__a2bb2o_1
X_1855_ _2128_/A _1865_/B _2350_/A VGND VGND VPWR VPWR _1855_/X sky130_fd_sc_hd__or3_1
X_1786_ _2243_/A VGND VGND VPWR VPWR _2374_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2512__A1 _2836_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2407_ _1464_/X _1682_/A _1469_/Y _2537_/A VGND VGND VPWR VPWR _2447_/A sky130_fd_sc_hd__o211a_4
XFILLER_58_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_2338_ _2338_/A VGND VGND VPWR VPWR _2747_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2177__A _2177_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2269_ _2362_/A VGND VGND VPWR VPWR _2289_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1512__C _1512_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2624__B _2626_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2028__A0 _2727_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_13_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2579__A1 _2357_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1955__S _1970_/S VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_4_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1554__A2 _1616_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1711__C1 _1710_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_29_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input25_A cpu_adr_i[30] VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_63_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__2931__CLK _2946_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1422__C _1454_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_21_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__2534__B _2534_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1490__A1 _1445_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1640_ _1712_/A VGND VGND VPWR VPWR _1640_/X sky130_fd_sc_hd__clkbuf_2
X_1571_ _1702_/A VGND VGND VPWR VPWR _1630_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__2700__D _2700_/D VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1545__A2 _1513_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_6_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2123_ _2708_/Q input68/X _2132_/S VGND VGND VPWR VPWR _2241_/B sky130_fd_sc_hd__mux2_1
XFILLER_48_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2054_ _2078_/A _2054_/B _2298_/A VGND VGND VPWR VPWR _2054_/X sky130_fd_sc_hd__or3_1
XFILLER_50_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1481__A1 _1803_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_22_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1769__C1 _1565_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1907_ _1911_/A _2668_/Q VGND VGND VPWR VPWR _1908_/A sky130_fd_sc_hd__and2_1
X_2887_ _2920_/CLK _2887_/D VGND VGND VPWR VPWR _2887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2430__B1 _2429_/Y VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1838_ _1807_/X _2542_/B _1789_/X _2925_/Q VGND VGND VPWR VPWR _2634_/B sky130_fd_sc_hd__o22ai_2
XANTENNA__2804__CLK _2809_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1769_ _1723_/X _2533_/A _1564_/X _1565_/X input97/X VGND VGND VPWR VPWR _1769_/Y
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_2_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1804__A _2039_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_57_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2619__B _2626_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__2635__A _2635_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_53_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2421__B1 _1597_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1775__A2 _1543_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2370__A _2370_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1492__B1_N _2866_/Q VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__1417__C _1461_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__2529__B _2529_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_0_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1433__B _1510_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output131_A _1580_/X VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_64_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2545__A _2548_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2810_ _2881_/CLK _2810_/D VGND VGND VPWR VPWR _2810_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2827__CLK _2901_/CLK VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_2741_ _2745_/CLK _2741_/D VGND VGND VPWR VPWR _2741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1766__A2 _2219_/B VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XANTENNA__2280__A _2280_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
Xclkbuf_leaf_17_CLK clkbuf_1_1_0_CLK/X VGND VGND VPWR VPWR _2847_/CLK sky130_fd_sc_hd__clkbuf_16
X_2672_ _2920_/CLK _2672_/D VGND VGND VPWR VPWR _2672_/Q sky130_fd_sc_hd__dfxtp_1
X_1623_ _1618_/X _1622_/Y _1593_/X _1595_/X VGND VGND VPWR VPWR _1623_/X sky130_fd_sc_hd__o211a_1
X_1554_ _1515_/A _1616_/A _2810_/Q VGND VGND VPWR VPWR _1554_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__1327__C _1335_/C VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
X_1485_ _1945_/A VGND VGND VPWR VPWR _1485_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_1049 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1624__A _1696_/A VGND VPWR VPWR VGND sky130_ef_sc_hd__fakediode_2
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

