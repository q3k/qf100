VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mkQF100Fabric
  CLASS BLOCK ;
  FOREIGN mkQF100Fabric ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 200.000 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END CLK
  PIN RST_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END RST_N
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 187.920 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 187.920 ;
    END
  END VPWR
  PIN cpu_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END cpu_ack_o
  PIN cpu_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END cpu_adr_i[0]
  PIN cpu_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END cpu_adr_i[10]
  PIN cpu_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END cpu_adr_i[11]
  PIN cpu_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END cpu_adr_i[12]
  PIN cpu_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END cpu_adr_i[13]
  PIN cpu_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END cpu_adr_i[14]
  PIN cpu_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END cpu_adr_i[15]
  PIN cpu_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END cpu_adr_i[16]
  PIN cpu_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END cpu_adr_i[17]
  PIN cpu_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END cpu_adr_i[18]
  PIN cpu_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END cpu_adr_i[19]
  PIN cpu_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END cpu_adr_i[1]
  PIN cpu_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END cpu_adr_i[20]
  PIN cpu_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END cpu_adr_i[21]
  PIN cpu_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END cpu_adr_i[22]
  PIN cpu_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END cpu_adr_i[23]
  PIN cpu_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END cpu_adr_i[24]
  PIN cpu_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END cpu_adr_i[25]
  PIN cpu_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END cpu_adr_i[26]
  PIN cpu_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END cpu_adr_i[27]
  PIN cpu_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END cpu_adr_i[28]
  PIN cpu_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END cpu_adr_i[29]
  PIN cpu_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END cpu_adr_i[2]
  PIN cpu_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END cpu_adr_i[30]
  PIN cpu_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END cpu_adr_i[31]
  PIN cpu_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END cpu_adr_i[3]
  PIN cpu_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END cpu_adr_i[4]
  PIN cpu_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END cpu_adr_i[5]
  PIN cpu_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END cpu_adr_i[6]
  PIN cpu_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END cpu_adr_i[7]
  PIN cpu_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END cpu_adr_i[8]
  PIN cpu_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END cpu_adr_i[9]
  PIN cpu_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END cpu_cyc_i
  PIN cpu_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END cpu_dat_i[0]
  PIN cpu_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END cpu_dat_i[10]
  PIN cpu_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END cpu_dat_i[11]
  PIN cpu_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 0.000 315.470 4.000 ;
    END
  END cpu_dat_i[12]
  PIN cpu_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 0.000 324.670 4.000 ;
    END
  END cpu_dat_i[13]
  PIN cpu_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END cpu_dat_i[14]
  PIN cpu_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END cpu_dat_i[15]
  PIN cpu_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END cpu_dat_i[16]
  PIN cpu_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END cpu_dat_i[17]
  PIN cpu_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END cpu_dat_i[18]
  PIN cpu_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END cpu_dat_i[19]
  PIN cpu_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END cpu_dat_i[1]
  PIN cpu_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 4.000 ;
    END
  END cpu_dat_i[20]
  PIN cpu_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END cpu_dat_i[21]
  PIN cpu_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END cpu_dat_i[22]
  PIN cpu_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END cpu_dat_i[23]
  PIN cpu_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 0.000 427.710 4.000 ;
    END
  END cpu_dat_i[24]
  PIN cpu_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 0.000 436.910 4.000 ;
    END
  END cpu_dat_i[25]
  PIN cpu_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END cpu_dat_i[26]
  PIN cpu_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END cpu_dat_i[27]
  PIN cpu_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 4.000 ;
    END
  END cpu_dat_i[28]
  PIN cpu_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END cpu_dat_i[29]
  PIN cpu_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END cpu_dat_i[2]
  PIN cpu_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 0.000 483.830 4.000 ;
    END
  END cpu_dat_i[30]
  PIN cpu_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END cpu_dat_i[31]
  PIN cpu_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END cpu_dat_i[3]
  PIN cpu_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END cpu_dat_i[4]
  PIN cpu_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END cpu_dat_i[5]
  PIN cpu_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 0.000 259.350 4.000 ;
    END
  END cpu_dat_i[6]
  PIN cpu_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END cpu_dat_i[7]
  PIN cpu_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 0.000 278.210 4.000 ;
    END
  END cpu_dat_i[8]
  PIN cpu_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END cpu_dat_i[9]
  PIN cpu_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END cpu_dat_o[0]
  PIN cpu_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END cpu_dat_o[10]
  PIN cpu_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 4.000 ;
    END
  END cpu_dat_o[11]
  PIN cpu_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END cpu_dat_o[12]
  PIN cpu_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END cpu_dat_o[13]
  PIN cpu_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END cpu_dat_o[14]
  PIN cpu_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END cpu_dat_o[15]
  PIN cpu_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END cpu_dat_o[16]
  PIN cpu_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 4.000 ;
    END
  END cpu_dat_o[17]
  PIN cpu_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.910 0.000 376.190 4.000 ;
    END
  END cpu_dat_o[18]
  PIN cpu_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END cpu_dat_o[19]
  PIN cpu_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END cpu_dat_o[1]
  PIN cpu_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END cpu_dat_o[20]
  PIN cpu_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 0.000 404.250 4.000 ;
    END
  END cpu_dat_o[21]
  PIN cpu_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END cpu_dat_o[22]
  PIN cpu_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 0.000 423.110 4.000 ;
    END
  END cpu_dat_o[23]
  PIN cpu_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 0.000 432.310 4.000 ;
    END
  END cpu_dat_o[24]
  PIN cpu_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END cpu_dat_o[25]
  PIN cpu_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END cpu_dat_o[26]
  PIN cpu_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 0.000 460.370 4.000 ;
    END
  END cpu_dat_o[27]
  PIN cpu_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 0.000 469.570 4.000 ;
    END
  END cpu_dat_o[28]
  PIN cpu_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END cpu_dat_o[29]
  PIN cpu_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END cpu_dat_o[2]
  PIN cpu_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 4.000 ;
    END
  END cpu_dat_o[30]
  PIN cpu_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 4.000 ;
    END
  END cpu_dat_o[31]
  PIN cpu_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END cpu_dat_o[3]
  PIN cpu_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END cpu_dat_o[4]
  PIN cpu_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END cpu_dat_o[5]
  PIN cpu_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END cpu_dat_o[6]
  PIN cpu_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END cpu_dat_o[7]
  PIN cpu_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END cpu_dat_o[8]
  PIN cpu_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END cpu_dat_o[9]
  PIN cpu_err_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END cpu_err_o
  PIN cpu_rty_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END cpu_rty_o
  PIN cpu_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END cpu_sel_i[0]
  PIN cpu_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END cpu_sel_i[1]
  PIN cpu_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END cpu_sel_i[2]
  PIN cpu_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END cpu_sel_i[3]
  PIN cpu_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END cpu_stb_i
  PIN cpu_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END cpu_we_i
  PIN spi_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 196.000 30.730 200.000 ;
    END
  END spi_ack_i
  PIN spi_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 196.000 44.990 200.000 ;
    END
  END spi_adr_o[0]
  PIN spi_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 196.000 91.910 200.000 ;
    END
  END spi_adr_o[10]
  PIN spi_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 196.000 96.970 200.000 ;
    END
  END spi_adr_o[11]
  PIN spi_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 196.000 101.570 200.000 ;
    END
  END spi_adr_o[12]
  PIN spi_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 196.000 106.170 200.000 ;
    END
  END spi_adr_o[13]
  PIN spi_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 196.000 110.770 200.000 ;
    END
  END spi_adr_o[14]
  PIN spi_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 196.000 115.830 200.000 ;
    END
  END spi_adr_o[15]
  PIN spi_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 196.000 120.430 200.000 ;
    END
  END spi_adr_o[16]
  PIN spi_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 196.000 125.030 200.000 ;
    END
  END spi_adr_o[17]
  PIN spi_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 196.000 129.630 200.000 ;
    END
  END spi_adr_o[18]
  PIN spi_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 196.000 134.690 200.000 ;
    END
  END spi_adr_o[19]
  PIN spi_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 196.000 49.590 200.000 ;
    END
  END spi_adr_o[1]
  PIN spi_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 196.000 139.290 200.000 ;
    END
  END spi_adr_o[20]
  PIN spi_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 196.000 143.890 200.000 ;
    END
  END spi_adr_o[21]
  PIN spi_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 196.000 148.490 200.000 ;
    END
  END spi_adr_o[22]
  PIN spi_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 196.000 153.550 200.000 ;
    END
  END spi_adr_o[23]
  PIN spi_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 196.000 158.150 200.000 ;
    END
  END spi_adr_o[24]
  PIN spi_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 196.000 162.750 200.000 ;
    END
  END spi_adr_o[25]
  PIN spi_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 196.000 167.350 200.000 ;
    END
  END spi_adr_o[26]
  PIN spi_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 196.000 172.410 200.000 ;
    END
  END spi_adr_o[27]
  PIN spi_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 196.000 177.010 200.000 ;
    END
  END spi_adr_o[28]
  PIN spi_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 196.000 181.610 200.000 ;
    END
  END spi_adr_o[29]
  PIN spi_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 196.000 54.190 200.000 ;
    END
  END spi_adr_o[2]
  PIN spi_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 196.000 186.210 200.000 ;
    END
  END spi_adr_o[30]
  PIN spi_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 196.000 191.270 200.000 ;
    END
  END spi_adr_o[31]
  PIN spi_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 196.000 59.250 200.000 ;
    END
  END spi_adr_o[3]
  PIN spi_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 196.000 63.850 200.000 ;
    END
  END spi_adr_o[4]
  PIN spi_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 196.000 68.450 200.000 ;
    END
  END spi_adr_o[5]
  PIN spi_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 196.000 73.050 200.000 ;
    END
  END spi_adr_o[6]
  PIN spi_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 196.000 78.110 200.000 ;
    END
  END spi_adr_o[7]
  PIN spi_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 196.000 82.710 200.000 ;
    END
  END spi_adr_o[8]
  PIN spi_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 196.000 87.310 200.000 ;
    END
  END spi_adr_o[9]
  PIN spi_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 196.000 2.670 200.000 ;
    END
  END spi_cyc_o
  PIN spi_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 196.000 195.870 200.000 ;
    END
  END spi_dat_i[0]
  PIN spi_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 196.000 290.170 200.000 ;
    END
  END spi_dat_i[10]
  PIN spi_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 196.000 299.830 200.000 ;
    END
  END spi_dat_i[11]
  PIN spi_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 196.000 309.030 200.000 ;
    END
  END spi_dat_i[12]
  PIN spi_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 196.000 318.690 200.000 ;
    END
  END spi_dat_i[13]
  PIN spi_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 196.000 327.890 200.000 ;
    END
  END spi_dat_i[14]
  PIN spi_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 196.000 337.550 200.000 ;
    END
  END spi_dat_i[15]
  PIN spi_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 196.000 346.750 200.000 ;
    END
  END spi_dat_i[16]
  PIN spi_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 196.000 356.410 200.000 ;
    END
  END spi_dat_i[17]
  PIN spi_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 196.000 365.610 200.000 ;
    END
  END spi_dat_i[18]
  PIN spi_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 196.000 375.270 200.000 ;
    END
  END spi_dat_i[19]
  PIN spi_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 196.000 205.070 200.000 ;
    END
  END spi_dat_i[1]
  PIN spi_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 196.000 384.470 200.000 ;
    END
  END spi_dat_i[20]
  PIN spi_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 196.000 394.130 200.000 ;
    END
  END spi_dat_i[21]
  PIN spi_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 196.000 403.330 200.000 ;
    END
  END spi_dat_i[22]
  PIN spi_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 196.000 412.990 200.000 ;
    END
  END spi_dat_i[23]
  PIN spi_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 196.000 422.190 200.000 ;
    END
  END spi_dat_i[24]
  PIN spi_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 196.000 431.850 200.000 ;
    END
  END spi_dat_i[25]
  PIN spi_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 196.000 441.050 200.000 ;
    END
  END spi_dat_i[26]
  PIN spi_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 196.000 450.710 200.000 ;
    END
  END spi_dat_i[27]
  PIN spi_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 196.000 459.910 200.000 ;
    END
  END spi_dat_i[28]
  PIN spi_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 196.000 469.570 200.000 ;
    END
  END spi_dat_i[29]
  PIN spi_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 196.000 214.730 200.000 ;
    END
  END spi_dat_i[2]
  PIN spi_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 196.000 478.770 200.000 ;
    END
  END spi_dat_i[30]
  PIN spi_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 196.000 488.430 200.000 ;
    END
  END spi_dat_i[31]
  PIN spi_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 196.000 223.930 200.000 ;
    END
  END spi_dat_i[3]
  PIN spi_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 196.000 233.590 200.000 ;
    END
  END spi_dat_i[4]
  PIN spi_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 196.000 242.790 200.000 ;
    END
  END spi_dat_i[5]
  PIN spi_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 196.000 252.450 200.000 ;
    END
  END spi_dat_i[6]
  PIN spi_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 196.000 262.110 200.000 ;
    END
  END spi_dat_i[7]
  PIN spi_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 196.000 271.310 200.000 ;
    END
  END spi_dat_i[8]
  PIN spi_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 196.000 280.970 200.000 ;
    END
  END spi_dat_i[9]
  PIN spi_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 196.000 200.470 200.000 ;
    END
  END spi_dat_o[0]
  PIN spi_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 196.000 294.770 200.000 ;
    END
  END spi_dat_o[10]
  PIN spi_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 196.000 304.430 200.000 ;
    END
  END spi_dat_o[11]
  PIN spi_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 196.000 313.630 200.000 ;
    END
  END spi_dat_o[12]
  PIN spi_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 196.000 323.290 200.000 ;
    END
  END spi_dat_o[13]
  PIN spi_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 196.000 332.490 200.000 ;
    END
  END spi_dat_o[14]
  PIN spi_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 196.000 342.150 200.000 ;
    END
  END spi_dat_o[15]
  PIN spi_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 196.000 351.350 200.000 ;
    END
  END spi_dat_o[16]
  PIN spi_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 196.000 361.010 200.000 ;
    END
  END spi_dat_o[17]
  PIN spi_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 196.000 370.210 200.000 ;
    END
  END spi_dat_o[18]
  PIN spi_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 196.000 379.870 200.000 ;
    END
  END spi_dat_o[19]
  PIN spi_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 196.000 210.130 200.000 ;
    END
  END spi_dat_o[1]
  PIN spi_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 196.000 389.070 200.000 ;
    END
  END spi_dat_o[20]
  PIN spi_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 196.000 398.730 200.000 ;
    END
  END spi_dat_o[21]
  PIN spi_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 196.000 407.930 200.000 ;
    END
  END spi_dat_o[22]
  PIN spi_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 196.000 417.590 200.000 ;
    END
  END spi_dat_o[23]
  PIN spi_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 196.000 426.790 200.000 ;
    END
  END spi_dat_o[24]
  PIN spi_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 196.000 436.450 200.000 ;
    END
  END spi_dat_o[25]
  PIN spi_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 196.000 445.650 200.000 ;
    END
  END spi_dat_o[26]
  PIN spi_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 196.000 455.310 200.000 ;
    END
  END spi_dat_o[27]
  PIN spi_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 196.000 464.510 200.000 ;
    END
  END spi_dat_o[28]
  PIN spi_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 196.000 474.170 200.000 ;
    END
  END spi_dat_o[29]
  PIN spi_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 196.000 219.330 200.000 ;
    END
  END spi_dat_o[2]
  PIN spi_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 196.000 483.370 200.000 ;
    END
  END spi_dat_o[30]
  PIN spi_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 196.000 493.030 200.000 ;
    END
  END spi_dat_o[31]
  PIN spi_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 196.000 228.990 200.000 ;
    END
  END spi_dat_o[3]
  PIN spi_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 196.000 238.190 200.000 ;
    END
  END spi_dat_o[4]
  PIN spi_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 196.000 247.850 200.000 ;
    END
  END spi_dat_o[5]
  PIN spi_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 196.000 257.050 200.000 ;
    END
  END spi_dat_o[6]
  PIN spi_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 196.000 266.710 200.000 ;
    END
  END spi_dat_o[7]
  PIN spi_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 196.000 275.910 200.000 ;
    END
  END spi_dat_o[8]
  PIN spi_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 196.000 285.570 200.000 ;
    END
  END spi_dat_o[9]
  PIN spi_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 196.000 35.330 200.000 ;
    END
  END spi_err_i
  PIN spi_rty_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 196.000 40.390 200.000 ;
    END
  END spi_rty_i
  PIN spi_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 196.000 11.870 200.000 ;
    END
  END spi_sel_o[0]
  PIN spi_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 196.000 16.470 200.000 ;
    END
  END spi_sel_o[1]
  PIN spi_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 196.000 21.530 200.000 ;
    END
  END spi_sel_o[2]
  PIN spi_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 196.000 26.130 200.000 ;
    END
  END spi_sel_o[3]
  PIN spi_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 196.000 7.270 200.000 ;
    END
  END spi_stb_o
  PIN spi_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 196.000 497.630 200.000 ;
    END
  END spi_we_o
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 187.765 ;
      LAYER met1 ;
        RECT 2.370 8.540 497.650 187.920 ;
      LAYER met2 ;
        RECT 0.090 195.720 2.110 196.250 ;
        RECT 2.950 195.720 6.710 196.250 ;
        RECT 7.550 195.720 11.310 196.250 ;
        RECT 12.150 195.720 15.910 196.250 ;
        RECT 16.750 195.720 20.970 196.250 ;
        RECT 21.810 195.720 25.570 196.250 ;
        RECT 26.410 195.720 30.170 196.250 ;
        RECT 31.010 195.720 34.770 196.250 ;
        RECT 35.610 195.720 39.830 196.250 ;
        RECT 40.670 195.720 44.430 196.250 ;
        RECT 45.270 195.720 49.030 196.250 ;
        RECT 49.870 195.720 53.630 196.250 ;
        RECT 54.470 195.720 58.690 196.250 ;
        RECT 59.530 195.720 63.290 196.250 ;
        RECT 64.130 195.720 67.890 196.250 ;
        RECT 68.730 195.720 72.490 196.250 ;
        RECT 73.330 195.720 77.550 196.250 ;
        RECT 78.390 195.720 82.150 196.250 ;
        RECT 82.990 195.720 86.750 196.250 ;
        RECT 87.590 195.720 91.350 196.250 ;
        RECT 92.190 195.720 96.410 196.250 ;
        RECT 97.250 195.720 101.010 196.250 ;
        RECT 101.850 195.720 105.610 196.250 ;
        RECT 106.450 195.720 110.210 196.250 ;
        RECT 111.050 195.720 115.270 196.250 ;
        RECT 116.110 195.720 119.870 196.250 ;
        RECT 120.710 195.720 124.470 196.250 ;
        RECT 125.310 195.720 129.070 196.250 ;
        RECT 129.910 195.720 134.130 196.250 ;
        RECT 134.970 195.720 138.730 196.250 ;
        RECT 139.570 195.720 143.330 196.250 ;
        RECT 144.170 195.720 147.930 196.250 ;
        RECT 148.770 195.720 152.990 196.250 ;
        RECT 153.830 195.720 157.590 196.250 ;
        RECT 158.430 195.720 162.190 196.250 ;
        RECT 163.030 195.720 166.790 196.250 ;
        RECT 167.630 195.720 171.850 196.250 ;
        RECT 172.690 195.720 176.450 196.250 ;
        RECT 177.290 195.720 181.050 196.250 ;
        RECT 181.890 195.720 185.650 196.250 ;
        RECT 186.490 195.720 190.710 196.250 ;
        RECT 191.550 195.720 195.310 196.250 ;
        RECT 196.150 195.720 199.910 196.250 ;
        RECT 200.750 195.720 204.510 196.250 ;
        RECT 205.350 195.720 209.570 196.250 ;
        RECT 210.410 195.720 214.170 196.250 ;
        RECT 215.010 195.720 218.770 196.250 ;
        RECT 219.610 195.720 223.370 196.250 ;
        RECT 224.210 195.720 228.430 196.250 ;
        RECT 229.270 195.720 233.030 196.250 ;
        RECT 233.870 195.720 237.630 196.250 ;
        RECT 238.470 195.720 242.230 196.250 ;
        RECT 243.070 195.720 247.290 196.250 ;
        RECT 248.130 195.720 251.890 196.250 ;
        RECT 252.730 195.720 256.490 196.250 ;
        RECT 257.330 195.720 261.550 196.250 ;
        RECT 262.390 195.720 266.150 196.250 ;
        RECT 266.990 195.720 270.750 196.250 ;
        RECT 271.590 195.720 275.350 196.250 ;
        RECT 276.190 195.720 280.410 196.250 ;
        RECT 281.250 195.720 285.010 196.250 ;
        RECT 285.850 195.720 289.610 196.250 ;
        RECT 290.450 195.720 294.210 196.250 ;
        RECT 295.050 195.720 299.270 196.250 ;
        RECT 300.110 195.720 303.870 196.250 ;
        RECT 304.710 195.720 308.470 196.250 ;
        RECT 309.310 195.720 313.070 196.250 ;
        RECT 313.910 195.720 318.130 196.250 ;
        RECT 318.970 195.720 322.730 196.250 ;
        RECT 323.570 195.720 327.330 196.250 ;
        RECT 328.170 195.720 331.930 196.250 ;
        RECT 332.770 195.720 336.990 196.250 ;
        RECT 337.830 195.720 341.590 196.250 ;
        RECT 342.430 195.720 346.190 196.250 ;
        RECT 347.030 195.720 350.790 196.250 ;
        RECT 351.630 195.720 355.850 196.250 ;
        RECT 356.690 195.720 360.450 196.250 ;
        RECT 361.290 195.720 365.050 196.250 ;
        RECT 365.890 195.720 369.650 196.250 ;
        RECT 370.490 195.720 374.710 196.250 ;
        RECT 375.550 195.720 379.310 196.250 ;
        RECT 380.150 195.720 383.910 196.250 ;
        RECT 384.750 195.720 388.510 196.250 ;
        RECT 389.350 195.720 393.570 196.250 ;
        RECT 394.410 195.720 398.170 196.250 ;
        RECT 399.010 195.720 402.770 196.250 ;
        RECT 403.610 195.720 407.370 196.250 ;
        RECT 408.210 195.720 412.430 196.250 ;
        RECT 413.270 195.720 417.030 196.250 ;
        RECT 417.870 195.720 421.630 196.250 ;
        RECT 422.470 195.720 426.230 196.250 ;
        RECT 427.070 195.720 431.290 196.250 ;
        RECT 432.130 195.720 435.890 196.250 ;
        RECT 436.730 195.720 440.490 196.250 ;
        RECT 441.330 195.720 445.090 196.250 ;
        RECT 445.930 195.720 450.150 196.250 ;
        RECT 450.990 195.720 454.750 196.250 ;
        RECT 455.590 195.720 459.350 196.250 ;
        RECT 460.190 195.720 463.950 196.250 ;
        RECT 464.790 195.720 469.010 196.250 ;
        RECT 469.850 195.720 473.610 196.250 ;
        RECT 474.450 195.720 478.210 196.250 ;
        RECT 479.050 195.720 482.810 196.250 ;
        RECT 483.650 195.720 487.870 196.250 ;
        RECT 488.710 195.720 492.470 196.250 ;
        RECT 493.310 195.720 497.070 196.250 ;
        RECT 0.090 4.280 497.620 195.720 ;
        RECT 0.090 3.670 2.110 4.280 ;
        RECT 2.950 3.670 6.710 4.280 ;
        RECT 7.550 3.670 11.310 4.280 ;
        RECT 12.150 3.670 15.910 4.280 ;
        RECT 16.750 3.670 20.510 4.280 ;
        RECT 21.350 3.670 25.110 4.280 ;
        RECT 25.950 3.670 29.710 4.280 ;
        RECT 30.550 3.670 34.770 4.280 ;
        RECT 35.610 3.670 39.370 4.280 ;
        RECT 40.210 3.670 43.970 4.280 ;
        RECT 44.810 3.670 48.570 4.280 ;
        RECT 49.410 3.670 53.170 4.280 ;
        RECT 54.010 3.670 57.770 4.280 ;
        RECT 58.610 3.670 62.830 4.280 ;
        RECT 63.670 3.670 67.430 4.280 ;
        RECT 68.270 3.670 72.030 4.280 ;
        RECT 72.870 3.670 76.630 4.280 ;
        RECT 77.470 3.670 81.230 4.280 ;
        RECT 82.070 3.670 85.830 4.280 ;
        RECT 86.670 3.670 90.890 4.280 ;
        RECT 91.730 3.670 95.490 4.280 ;
        RECT 96.330 3.670 100.090 4.280 ;
        RECT 100.930 3.670 104.690 4.280 ;
        RECT 105.530 3.670 109.290 4.280 ;
        RECT 110.130 3.670 113.890 4.280 ;
        RECT 114.730 3.670 118.490 4.280 ;
        RECT 119.330 3.670 123.550 4.280 ;
        RECT 124.390 3.670 128.150 4.280 ;
        RECT 128.990 3.670 132.750 4.280 ;
        RECT 133.590 3.670 137.350 4.280 ;
        RECT 138.190 3.670 141.950 4.280 ;
        RECT 142.790 3.670 146.550 4.280 ;
        RECT 147.390 3.670 151.610 4.280 ;
        RECT 152.450 3.670 156.210 4.280 ;
        RECT 157.050 3.670 160.810 4.280 ;
        RECT 161.650 3.670 165.410 4.280 ;
        RECT 166.250 3.670 170.010 4.280 ;
        RECT 170.850 3.670 174.610 4.280 ;
        RECT 175.450 3.670 179.670 4.280 ;
        RECT 180.510 3.670 184.270 4.280 ;
        RECT 185.110 3.670 188.870 4.280 ;
        RECT 189.710 3.670 193.470 4.280 ;
        RECT 194.310 3.670 198.070 4.280 ;
        RECT 198.910 3.670 202.670 4.280 ;
        RECT 203.510 3.670 207.270 4.280 ;
        RECT 208.110 3.670 212.330 4.280 ;
        RECT 213.170 3.670 216.930 4.280 ;
        RECT 217.770 3.670 221.530 4.280 ;
        RECT 222.370 3.670 226.130 4.280 ;
        RECT 226.970 3.670 230.730 4.280 ;
        RECT 231.570 3.670 235.330 4.280 ;
        RECT 236.170 3.670 240.390 4.280 ;
        RECT 241.230 3.670 244.990 4.280 ;
        RECT 245.830 3.670 249.590 4.280 ;
        RECT 250.430 3.670 254.190 4.280 ;
        RECT 255.030 3.670 258.790 4.280 ;
        RECT 259.630 3.670 263.390 4.280 ;
        RECT 264.230 3.670 268.450 4.280 ;
        RECT 269.290 3.670 273.050 4.280 ;
        RECT 273.890 3.670 277.650 4.280 ;
        RECT 278.490 3.670 282.250 4.280 ;
        RECT 283.090 3.670 286.850 4.280 ;
        RECT 287.690 3.670 291.450 4.280 ;
        RECT 292.290 3.670 296.510 4.280 ;
        RECT 297.350 3.670 301.110 4.280 ;
        RECT 301.950 3.670 305.710 4.280 ;
        RECT 306.550 3.670 310.310 4.280 ;
        RECT 311.150 3.670 314.910 4.280 ;
        RECT 315.750 3.670 319.510 4.280 ;
        RECT 320.350 3.670 324.110 4.280 ;
        RECT 324.950 3.670 329.170 4.280 ;
        RECT 330.010 3.670 333.770 4.280 ;
        RECT 334.610 3.670 338.370 4.280 ;
        RECT 339.210 3.670 342.970 4.280 ;
        RECT 343.810 3.670 347.570 4.280 ;
        RECT 348.410 3.670 352.170 4.280 ;
        RECT 353.010 3.670 357.230 4.280 ;
        RECT 358.070 3.670 361.830 4.280 ;
        RECT 362.670 3.670 366.430 4.280 ;
        RECT 367.270 3.670 371.030 4.280 ;
        RECT 371.870 3.670 375.630 4.280 ;
        RECT 376.470 3.670 380.230 4.280 ;
        RECT 381.070 3.670 385.290 4.280 ;
        RECT 386.130 3.670 389.890 4.280 ;
        RECT 390.730 3.670 394.490 4.280 ;
        RECT 395.330 3.670 399.090 4.280 ;
        RECT 399.930 3.670 403.690 4.280 ;
        RECT 404.530 3.670 408.290 4.280 ;
        RECT 409.130 3.670 412.890 4.280 ;
        RECT 413.730 3.670 417.950 4.280 ;
        RECT 418.790 3.670 422.550 4.280 ;
        RECT 423.390 3.670 427.150 4.280 ;
        RECT 427.990 3.670 431.750 4.280 ;
        RECT 432.590 3.670 436.350 4.280 ;
        RECT 437.190 3.670 440.950 4.280 ;
        RECT 441.790 3.670 446.010 4.280 ;
        RECT 446.850 3.670 450.610 4.280 ;
        RECT 451.450 3.670 455.210 4.280 ;
        RECT 456.050 3.670 459.810 4.280 ;
        RECT 460.650 3.670 464.410 4.280 ;
        RECT 465.250 3.670 469.010 4.280 ;
        RECT 469.850 3.670 474.070 4.280 ;
        RECT 474.910 3.670 478.670 4.280 ;
        RECT 479.510 3.670 483.270 4.280 ;
        RECT 484.110 3.670 487.870 4.280 ;
        RECT 488.710 3.670 492.470 4.280 ;
        RECT 493.310 3.670 497.070 4.280 ;
      LAYER met3 ;
        RECT 0.065 101.000 483.440 187.845 ;
        RECT 4.400 99.600 483.440 101.000 ;
        RECT 0.065 8.335 483.440 99.600 ;
      LAYER met4 ;
        RECT 48.135 41.655 97.440 66.465 ;
        RECT 99.840 41.655 174.240 66.465 ;
        RECT 176.640 41.655 192.905 66.465 ;
  END
END mkQF100Fabric
END LIBRARY

