magic
tech sky130A
magscale 1 2
timestamp 1647563318
<< viali >>
rect 10149 28713 10183 28747
rect 23121 28713 23155 28747
rect 8125 28645 8159 28679
rect 13737 28645 13771 28679
rect 20085 28645 20119 28679
rect 21465 28645 21499 28679
rect 13921 28577 13955 28611
rect 19717 28577 19751 28611
rect 8125 28509 8159 28543
rect 8401 28509 8435 28543
rect 9505 28509 9539 28543
rect 10333 28509 10367 28543
rect 10977 28509 11011 28543
rect 11345 28509 11379 28543
rect 12357 28509 12391 28543
rect 13001 28509 13035 28543
rect 13185 28509 13219 28543
rect 13645 28509 13679 28543
rect 14565 28509 14599 28543
rect 15025 28509 15059 28543
rect 16037 28509 16071 28543
rect 16497 28509 16531 28543
rect 17049 28509 17083 28543
rect 17509 28509 17543 28543
rect 18153 28509 18187 28543
rect 18705 28509 18739 28543
rect 18889 28509 18923 28543
rect 20269 28509 20303 28543
rect 20913 28509 20947 28543
rect 21189 28509 21223 28543
rect 21649 28509 21683 28543
rect 22201 28509 22235 28543
rect 22661 28509 22695 28543
rect 23305 28509 23339 28543
rect 23581 28509 23615 28543
rect 27353 28509 27387 28543
rect 8585 28441 8619 28475
rect 8769 28441 8803 28475
rect 9873 28441 9907 28475
rect 8309 28373 8343 28407
rect 10793 28373 10827 28407
rect 11161 28373 11195 28407
rect 11897 28373 11931 28407
rect 12173 28373 12207 28407
rect 13093 28373 13127 28407
rect 13921 28373 13955 28407
rect 14841 28373 14875 28407
rect 15577 28373 15611 28407
rect 15853 28373 15887 28407
rect 16313 28373 16347 28407
rect 17325 28373 17359 28407
rect 17969 28373 18003 28407
rect 19073 28373 19107 28407
rect 20729 28373 20763 28407
rect 22477 28373 22511 28407
rect 27169 28373 27203 28407
rect 4353 28169 4387 28203
rect 7450 28101 7484 28135
rect 2697 28033 2731 28067
rect 3157 28033 3191 28067
rect 4445 28033 4479 28067
rect 4712 28033 4746 28067
rect 9597 28033 9631 28067
rect 9864 28033 9898 28067
rect 12164 28033 12198 28067
rect 14289 28033 14323 28067
rect 14545 28033 14579 28067
rect 16681 28033 16715 28067
rect 16948 28033 16982 28067
rect 18521 28033 18555 28067
rect 18777 28033 18811 28067
rect 20545 28033 20579 28067
rect 21189 28033 21223 28067
rect 22569 28033 22603 28067
rect 23857 28033 23891 28067
rect 26433 28033 26467 28067
rect 26985 28033 27019 28067
rect 27169 28033 27203 28067
rect 7205 27965 7239 27999
rect 11897 27965 11931 27999
rect 26985 27897 27019 27931
rect 2973 27829 3007 27863
rect 5825 27829 5859 27863
rect 8585 27829 8619 27863
rect 10977 27829 11011 27863
rect 13277 27829 13311 27863
rect 15669 27829 15703 27863
rect 18061 27829 18095 27863
rect 19901 27829 19935 27863
rect 20361 27829 20395 27863
rect 21005 27829 21039 27863
rect 22385 27829 22419 27863
rect 23305 27829 23339 27863
rect 23673 27829 23707 27863
rect 26249 27829 26283 27863
rect 13001 27625 13035 27659
rect 18705 27625 18739 27659
rect 21741 27625 21775 27659
rect 1777 27557 1811 27591
rect 13277 27557 13311 27591
rect 15945 27557 15979 27591
rect 23305 27557 23339 27591
rect 4445 27489 4479 27523
rect 13185 27489 13219 27523
rect 18337 27489 18371 27523
rect 21833 27489 21867 27523
rect 1961 27421 1995 27455
rect 2605 27421 2639 27455
rect 3249 27421 3283 27455
rect 4537 27421 4571 27455
rect 4721 27421 4755 27455
rect 5365 27421 5399 27455
rect 5825 27421 5859 27455
rect 6469 27421 6503 27455
rect 8953 27421 8987 27455
rect 9220 27421 9254 27455
rect 11069 27421 11103 27455
rect 11325 27421 11359 27455
rect 12909 27421 12943 27455
rect 13553 27421 13587 27455
rect 13645 27421 13679 27455
rect 13737 27421 13771 27455
rect 13921 27421 13955 27455
rect 15393 27421 15427 27455
rect 15853 27421 15887 27455
rect 16129 27421 16163 27455
rect 17417 27421 17451 27455
rect 18521 27421 18555 27455
rect 19257 27421 19291 27455
rect 21373 27421 21407 27455
rect 21557 27421 21591 27455
rect 22100 27421 22134 27455
rect 23305 27421 23339 27455
rect 23489 27421 23523 27455
rect 23857 27421 23891 27455
rect 24593 27421 24627 27455
rect 25237 27421 25271 27455
rect 25973 27421 26007 27455
rect 26617 27421 26651 27455
rect 27077 27421 27111 27455
rect 6714 27353 6748 27387
rect 16957 27353 16991 27387
rect 19524 27353 19558 27387
rect 2421 27285 2455 27319
rect 3065 27285 3099 27319
rect 3985 27285 4019 27319
rect 4629 27285 4663 27319
rect 5641 27285 5675 27319
rect 7849 27285 7883 27319
rect 10333 27285 10367 27319
rect 12449 27285 12483 27319
rect 13185 27285 13219 27319
rect 14933 27285 14967 27319
rect 15209 27285 15243 27319
rect 15669 27285 15703 27319
rect 16497 27285 16531 27319
rect 17233 27285 17267 27319
rect 20637 27285 20671 27319
rect 23213 27285 23247 27319
rect 23673 27285 23707 27319
rect 24409 27285 24443 27319
rect 25053 27285 25087 27319
rect 25789 27285 25823 27319
rect 26433 27285 26467 27319
rect 27261 27285 27295 27319
rect 5273 27081 5307 27115
rect 6377 27081 6411 27115
rect 8171 27081 8205 27115
rect 11897 27081 11931 27115
rect 12541 27081 12575 27115
rect 19073 27081 19107 27115
rect 27169 27081 27203 27115
rect 3341 27013 3375 27047
rect 16926 27013 16960 27047
rect 18797 27013 18831 27047
rect 21925 27013 21959 27047
rect 1593 26945 1627 26979
rect 2329 26945 2363 26979
rect 3801 26945 3835 26979
rect 4068 26945 4102 26979
rect 5549 26945 5583 26979
rect 5638 26945 5672 26979
rect 5738 26945 5772 26979
rect 5917 26945 5951 26979
rect 6653 26945 6687 26979
rect 6745 26945 6779 26979
rect 6858 26951 6892 26985
rect 7021 26945 7055 26979
rect 9229 26945 9263 26979
rect 10149 26945 10183 26979
rect 11529 26945 11563 26979
rect 11713 26945 11747 26979
rect 12725 26945 12759 26979
rect 12817 26945 12851 26979
rect 13001 26945 13035 26979
rect 13093 26945 13127 26979
rect 13737 26945 13771 26979
rect 13921 26945 13955 26979
rect 14013 26945 14047 26979
rect 14473 26945 14507 26979
rect 14740 26945 14774 26979
rect 16681 26945 16715 26979
rect 18521 26945 18555 26979
rect 18705 26945 18739 26979
rect 18889 26945 18923 26979
rect 19901 26945 19935 26979
rect 20168 26945 20202 26979
rect 21833 26945 21867 26979
rect 22017 26945 22051 26979
rect 22661 26945 22695 26979
rect 23305 26945 23339 26979
rect 23949 26945 23983 26979
rect 24409 26945 24443 26979
rect 24593 26945 24627 26979
rect 25789 26945 25823 26979
rect 26433 26945 26467 26979
rect 27353 26945 27387 26979
rect 7941 26877 7975 26911
rect 9321 26877 9355 26911
rect 10425 26877 10459 26911
rect 2145 26809 2179 26843
rect 22477 26809 22511 26843
rect 24409 26809 24443 26843
rect 1409 26741 1443 26775
rect 2697 26741 2731 26775
rect 2973 26741 3007 26775
rect 5181 26741 5215 26775
rect 9229 26741 9263 26775
rect 9597 26741 9631 26775
rect 13737 26741 13771 26775
rect 15853 26741 15887 26775
rect 18061 26741 18095 26775
rect 21281 26741 21315 26775
rect 23121 26741 23155 26775
rect 23765 26741 23799 26775
rect 25605 26741 25639 26775
rect 26249 26741 26283 26775
rect 4537 26537 4571 26571
rect 5549 26537 5583 26571
rect 9045 26537 9079 26571
rect 9965 26537 9999 26571
rect 14473 26537 14507 26571
rect 14565 26537 14599 26571
rect 16681 26537 16715 26571
rect 19809 26537 19843 26571
rect 21465 26537 21499 26571
rect 26249 26537 26283 26571
rect 1869 26469 1903 26503
rect 7757 26469 7791 26503
rect 15853 26469 15887 26503
rect 18153 26469 18187 26503
rect 20637 26469 20671 26503
rect 26893 26469 26927 26503
rect 3157 26401 3191 26435
rect 4077 26401 4111 26435
rect 4629 26401 4663 26435
rect 7849 26401 7883 26435
rect 11069 26401 11103 26435
rect 11437 26401 11471 26435
rect 12909 26401 12943 26435
rect 20269 26401 20303 26435
rect 21925 26401 21959 26435
rect 2053 26333 2087 26367
rect 3065 26333 3099 26367
rect 3249 26333 3283 26367
rect 3801 26333 3835 26367
rect 3985 26333 4019 26367
rect 4169 26333 4203 26367
rect 4353 26333 4387 26367
rect 4813 26333 4847 26367
rect 5089 26333 5123 26367
rect 5273 26333 5307 26367
rect 5549 26311 5583 26345
rect 6009 26333 6043 26367
rect 6193 26333 6227 26367
rect 7389 26333 7423 26367
rect 7573 26333 7607 26367
rect 7665 26333 7699 26367
rect 7941 26333 7975 26367
rect 9229 26333 9263 26367
rect 9505 26333 9539 26367
rect 10149 26333 10183 26367
rect 10425 26333 10459 26367
rect 10609 26333 10643 26367
rect 11253 26333 11287 26367
rect 11345 26333 11379 26367
rect 11529 26333 11563 26367
rect 12633 26333 12667 26367
rect 14105 26333 14139 26367
rect 14197 26333 14231 26367
rect 14565 26333 14599 26367
rect 15485 26333 15519 26367
rect 15669 26333 15703 26367
rect 16313 26333 16347 26367
rect 16497 26333 16531 26367
rect 17601 26333 17635 26367
rect 17969 26333 18003 26367
rect 19257 26333 19291 26367
rect 19441 26333 19475 26367
rect 19625 26333 19659 26367
rect 20453 26333 20487 26367
rect 21189 26333 21223 26367
rect 21281 26333 21315 26367
rect 24409 26333 24443 26367
rect 26433 26333 26467 26367
rect 27077 26333 27111 26367
rect 2421 26265 2455 26299
rect 5457 26265 5491 26299
rect 6745 26265 6779 26299
rect 17785 26265 17819 26299
rect 17877 26265 17911 26299
rect 19533 26265 19567 26299
rect 22192 26265 22226 26299
rect 24654 26265 24688 26299
rect 4997 26197 5031 26231
rect 6101 26197 6135 26231
rect 6837 26197 6871 26231
rect 9413 26197 9447 26231
rect 14289 26197 14323 26231
rect 23305 26197 23339 26231
rect 25789 26197 25823 26231
rect 8677 25993 8711 26027
rect 11989 25993 12023 26027
rect 13185 25993 13219 26027
rect 14105 25993 14139 26027
rect 15133 25993 15167 26027
rect 18153 25993 18187 26027
rect 19993 25993 20027 26027
rect 22385 25993 22419 26027
rect 24593 25993 24627 26027
rect 25421 25993 25455 26027
rect 2136 25925 2170 25959
rect 4721 25925 4755 25959
rect 8125 25925 8159 25959
rect 9045 25925 9079 25959
rect 10517 25925 10551 25959
rect 10701 25925 10735 25959
rect 13737 25925 13771 25959
rect 14933 25925 14967 25959
rect 17785 25925 17819 25959
rect 19625 25925 19659 25959
rect 22109 25925 22143 25959
rect 23489 25925 23523 25959
rect 3985 25857 4019 25891
rect 4169 25857 4203 25891
rect 4537 25857 4571 25891
rect 5365 25857 5399 25891
rect 5549 25857 5583 25891
rect 5641 25857 5675 25891
rect 6377 25857 6411 25891
rect 7941 25857 7975 25891
rect 8217 25857 8251 25891
rect 8861 25857 8895 25891
rect 9137 25857 9171 25891
rect 9597 25857 9631 25891
rect 9689 25857 9723 25891
rect 12173 25857 12207 25891
rect 12265 25857 12299 25891
rect 12541 25857 12575 25891
rect 13001 25857 13035 25891
rect 13277 25857 13311 25891
rect 13921 25857 13955 25891
rect 15761 25857 15795 25891
rect 16865 25857 16899 25891
rect 17141 25857 17175 25891
rect 17601 25857 17635 25891
rect 17877 25857 17911 25891
rect 17969 25857 18003 25891
rect 18797 25857 18831 25891
rect 18981 25857 19015 25891
rect 19441 25857 19475 25891
rect 19717 25857 19751 25891
rect 19809 25857 19843 25891
rect 20637 25857 20671 25891
rect 21097 25857 21131 25891
rect 21281 25857 21315 25891
rect 21833 25857 21867 25891
rect 22017 25857 22051 25891
rect 22201 25857 22235 25891
rect 23213 25857 23247 25891
rect 23397 25857 23431 25891
rect 23581 25857 23615 25891
rect 24409 25857 24443 25891
rect 25237 25857 25271 25891
rect 26341 25857 26375 25891
rect 27169 25857 27203 25891
rect 1869 25789 1903 25823
rect 4261 25789 4295 25823
rect 4353 25789 4387 25823
rect 6653 25789 6687 25823
rect 24225 25789 24259 25823
rect 25053 25789 25087 25823
rect 5181 25721 5215 25755
rect 7941 25721 7975 25755
rect 9965 25721 9999 25755
rect 13001 25721 13035 25755
rect 15301 25721 15335 25755
rect 16681 25721 16715 25755
rect 21097 25721 21131 25755
rect 23765 25721 23799 25755
rect 3249 25653 3283 25687
rect 6469 25653 6503 25687
rect 6929 25653 6963 25687
rect 9781 25653 9815 25687
rect 12449 25653 12483 25687
rect 15117 25653 15151 25687
rect 15945 25653 15979 25687
rect 18797 25653 18831 25687
rect 20453 25653 20487 25687
rect 26157 25653 26191 25687
rect 26985 25653 27019 25687
rect 1777 25449 1811 25483
rect 4261 25449 4295 25483
rect 9413 25449 9447 25483
rect 9873 25449 9907 25483
rect 12449 25449 12483 25483
rect 14381 25449 14415 25483
rect 15853 25449 15887 25483
rect 19717 25449 19751 25483
rect 22385 25449 22419 25483
rect 24961 25449 24995 25483
rect 2421 25381 2455 25415
rect 7021 25381 7055 25415
rect 7941 25381 7975 25415
rect 14565 25381 14599 25415
rect 16773 25381 16807 25415
rect 4629 25313 4663 25347
rect 4813 25313 4847 25347
rect 6009 25313 6043 25347
rect 12633 25313 12667 25347
rect 12817 25313 12851 25347
rect 15669 25313 15703 25347
rect 18153 25313 18187 25347
rect 20361 25313 20395 25347
rect 23305 25313 23339 25347
rect 25421 25313 25455 25347
rect 1961 25245 1995 25279
rect 2605 25245 2639 25279
rect 3249 25245 3283 25279
rect 4169 25245 4203 25279
rect 4353 25245 4387 25279
rect 5089 25245 5123 25279
rect 5733 25245 5767 25279
rect 5825 25245 5859 25279
rect 6837 25245 6871 25279
rect 9413 25245 9447 25279
rect 9597 25245 9631 25279
rect 9689 25245 9723 25279
rect 10333 25245 10367 25279
rect 12725 25245 12759 25279
rect 12909 25245 12943 25279
rect 15577 25245 15611 25279
rect 17877 25245 17911 25279
rect 21373 25245 21407 25279
rect 21833 25245 21867 25279
rect 22201 25245 22235 25279
rect 23029 25245 23063 25279
rect 24409 25245 24443 25279
rect 24593 25245 24627 25279
rect 24777 25245 24811 25279
rect 25688 25245 25722 25279
rect 3985 25177 4019 25211
rect 6009 25177 6043 25211
rect 7757 25177 7791 25211
rect 10600 25177 10634 25211
rect 14197 25177 14231 25211
rect 16497 25177 16531 25211
rect 20085 25177 20119 25211
rect 22017 25177 22051 25211
rect 22109 25177 22143 25211
rect 24681 25177 24715 25211
rect 3065 25109 3099 25143
rect 11713 25109 11747 25143
rect 14407 25109 14441 25143
rect 16957 25109 16991 25143
rect 20177 25109 20211 25143
rect 21189 25109 21223 25143
rect 26801 25109 26835 25143
rect 3157 24905 3191 24939
rect 5647 24905 5681 24939
rect 6745 24905 6779 24939
rect 9229 24905 9263 24939
rect 10241 24905 10275 24939
rect 10885 24905 10919 24939
rect 11713 24905 11747 24939
rect 18705 24905 18739 24939
rect 19165 24905 19199 24939
rect 19901 24905 19935 24939
rect 22017 24905 22051 24939
rect 4629 24837 4663 24871
rect 7481 24837 7515 24871
rect 12817 24837 12851 24871
rect 16773 24837 16807 24871
rect 20269 24837 20303 24871
rect 22477 24837 22511 24871
rect 13047 24803 13081 24837
rect 1777 24769 1811 24803
rect 2421 24769 2455 24803
rect 3249 24769 3283 24803
rect 3801 24769 3835 24803
rect 4445 24769 4479 24803
rect 5549 24769 5583 24803
rect 5733 24769 5767 24803
rect 5825 24769 5859 24803
rect 6377 24769 6411 24803
rect 7665 24769 7699 24803
rect 7757 24769 7791 24803
rect 8217 24769 8251 24803
rect 9045 24769 9079 24803
rect 9413 24769 9447 24803
rect 9597 24769 9631 24803
rect 10149 24769 10183 24803
rect 10793 24769 10827 24803
rect 10977 24769 11011 24803
rect 11529 24769 11563 24803
rect 11713 24769 11747 24803
rect 12173 24769 12207 24803
rect 12357 24769 12391 24803
rect 13645 24769 13679 24803
rect 14381 24769 14415 24803
rect 15209 24769 15243 24803
rect 16681 24769 16715 24803
rect 16865 24769 16899 24803
rect 17693 24769 17727 24803
rect 19073 24769 19107 24803
rect 21281 24769 21315 24803
rect 22385 24769 22419 24803
rect 23305 24769 23339 24803
rect 23581 24769 23615 24803
rect 24593 24769 24627 24803
rect 24777 24769 24811 24803
rect 24869 24769 24903 24803
rect 24961 24769 24995 24803
rect 25789 24769 25823 24803
rect 26433 24769 26467 24803
rect 27353 24769 27387 24803
rect 3525 24701 3559 24735
rect 6469 24701 6503 24735
rect 8493 24701 8527 24735
rect 15301 24701 15335 24735
rect 17417 24701 17451 24735
rect 19257 24701 19291 24735
rect 20361 24701 20395 24735
rect 20545 24701 20579 24735
rect 22661 24701 22695 24735
rect 2789 24633 2823 24667
rect 3341 24633 3375 24667
rect 7481 24633 7515 24667
rect 8309 24633 8343 24667
rect 8401 24633 8435 24667
rect 12265 24633 12299 24667
rect 13185 24633 13219 24667
rect 14565 24633 14599 24667
rect 1593 24565 1627 24599
rect 2237 24565 2271 24599
rect 3433 24565 3467 24599
rect 3617 24565 3651 24599
rect 4261 24565 4295 24599
rect 4813 24565 4847 24599
rect 6377 24565 6411 24599
rect 9413 24565 9447 24599
rect 13001 24565 13035 24599
rect 13737 24565 13771 24599
rect 15485 24565 15519 24599
rect 21097 24565 21131 24599
rect 25145 24565 25179 24599
rect 25605 24565 25639 24599
rect 26249 24565 26283 24599
rect 27169 24565 27203 24599
rect 3801 24361 3835 24395
rect 4721 24361 4755 24395
rect 5917 24361 5951 24395
rect 7573 24361 7607 24395
rect 9045 24361 9079 24395
rect 9873 24361 9907 24395
rect 12633 24361 12667 24395
rect 14841 24361 14875 24395
rect 17877 24361 17911 24395
rect 19257 24361 19291 24395
rect 21097 24361 21131 24395
rect 23029 24361 23063 24395
rect 25513 24361 25547 24395
rect 10333 24293 10367 24327
rect 16221 24293 16255 24327
rect 1409 24225 1443 24259
rect 5365 24225 5399 24259
rect 6561 24225 6595 24259
rect 7757 24225 7791 24259
rect 10885 24225 10919 24259
rect 15853 24225 15887 24259
rect 16313 24225 16347 24259
rect 17233 24225 17267 24259
rect 18521 24225 18555 24259
rect 19809 24225 19843 24259
rect 21649 24225 21683 24259
rect 23581 24225 23615 24259
rect 25973 24225 26007 24259
rect 3801 24157 3835 24191
rect 3985 24157 4019 24191
rect 7849 24157 7883 24191
rect 8217 24157 8251 24191
rect 8953 24157 8987 24191
rect 9137 24157 9171 24191
rect 10057 24157 10091 24191
rect 10149 24157 10183 24191
rect 10425 24157 10459 24191
rect 11161 24157 11195 24191
rect 13185 24157 13219 24191
rect 14381 24157 14415 24191
rect 14749 24157 14783 24191
rect 16773 24157 16807 24191
rect 17049 24157 17083 24191
rect 18245 24157 18279 24191
rect 19717 24157 19751 24191
rect 20637 24157 20671 24191
rect 21557 24157 21591 24191
rect 22477 24157 22511 24191
rect 24593 24157 24627 24191
rect 25145 24157 25179 24191
rect 25329 24157 25363 24191
rect 26240 24157 26274 24191
rect 1676 24089 1710 24123
rect 5089 24089 5123 24123
rect 6285 24089 6319 24123
rect 12541 24089 12575 24123
rect 21465 24089 21499 24123
rect 23489 24089 23523 24123
rect 2789 24021 2823 24055
rect 4169 24021 4203 24055
rect 5181 24021 5215 24055
rect 6377 24021 6411 24055
rect 7941 24021 7975 24055
rect 8125 24021 8159 24055
rect 13277 24021 13311 24055
rect 14565 24021 14599 24055
rect 17325 24021 17359 24055
rect 18337 24021 18371 24055
rect 19625 24021 19659 24055
rect 20453 24021 20487 24055
rect 22293 24021 22327 24055
rect 23397 24021 23431 24055
rect 24409 24021 24443 24055
rect 27353 24021 27387 24055
rect 1961 23817 1995 23851
rect 3525 23817 3559 23851
rect 5733 23817 5767 23851
rect 6377 23817 6411 23851
rect 6745 23817 6779 23851
rect 7573 23817 7607 23851
rect 7941 23817 7975 23851
rect 11805 23817 11839 23851
rect 15685 23817 15719 23851
rect 18981 23817 19015 23851
rect 22293 23817 22327 23851
rect 23213 23817 23247 23851
rect 25053 23817 25087 23851
rect 25421 23817 25455 23851
rect 4537 23749 4571 23783
rect 8125 23749 8159 23783
rect 15485 23749 15519 23783
rect 18521 23749 18555 23783
rect 19809 23749 19843 23783
rect 25513 23749 25547 23783
rect 27169 23749 27203 23783
rect 1685 23681 1719 23715
rect 2145 23681 2179 23715
rect 3433 23681 3467 23715
rect 3801 23681 3835 23715
rect 4261 23681 4295 23715
rect 5641 23681 5675 23715
rect 6837 23681 6871 23715
rect 8861 23681 8895 23715
rect 9597 23681 9631 23715
rect 9781 23681 9815 23715
rect 9873 23681 9907 23715
rect 10149 23681 10183 23715
rect 10793 23681 10827 23715
rect 11529 23681 11563 23715
rect 12532 23681 12566 23715
rect 14381 23681 14415 23715
rect 17233 23681 17267 23715
rect 18797 23681 18831 23715
rect 19625 23681 19659 23715
rect 21833 23681 21867 23715
rect 22109 23681 22143 23715
rect 22753 23681 22787 23715
rect 23029 23681 23063 23715
rect 24041 23681 24075 23715
rect 26433 23681 26467 23715
rect 3617 23613 3651 23647
rect 4537 23613 4571 23647
rect 7021 23613 7055 23647
rect 7757 23613 7791 23647
rect 7849 23613 7883 23647
rect 8217 23613 8251 23647
rect 8953 23613 8987 23647
rect 9137 23613 9171 23647
rect 9965 23613 9999 23647
rect 11805 23613 11839 23647
rect 12265 23613 12299 23647
rect 14105 23613 14139 23647
rect 17325 23613 17359 23647
rect 18705 23613 18739 23647
rect 20269 23613 20303 23647
rect 20545 23613 20579 23647
rect 21925 23613 21959 23647
rect 22937 23613 22971 23647
rect 23765 23613 23799 23647
rect 25605 23613 25639 23647
rect 3801 23545 3835 23579
rect 10333 23545 10367 23579
rect 11621 23545 11655 23579
rect 13645 23545 13679 23579
rect 15853 23545 15887 23579
rect 26249 23545 26283 23579
rect 2789 23477 2823 23511
rect 4353 23477 4387 23511
rect 9045 23477 9079 23511
rect 10885 23477 10919 23511
rect 15669 23477 15703 23511
rect 17233 23477 17267 23511
rect 17601 23477 17635 23511
rect 18521 23477 18555 23511
rect 22017 23477 22051 23511
rect 22753 23477 22787 23511
rect 27261 23477 27295 23511
rect 2513 23273 2547 23307
rect 5917 23273 5951 23307
rect 6837 23273 6871 23307
rect 10333 23273 10367 23307
rect 12173 23273 12207 23307
rect 15209 23273 15243 23307
rect 19349 23273 19383 23307
rect 21005 23273 21039 23307
rect 22569 23273 22603 23307
rect 22753 23273 22787 23307
rect 23213 23273 23247 23307
rect 24409 23273 24443 23307
rect 7481 23205 7515 23239
rect 14657 23205 14691 23239
rect 19717 23205 19751 23239
rect 23673 23205 23707 23239
rect 3065 23137 3099 23171
rect 4353 23137 4387 23171
rect 9045 23137 9079 23171
rect 11621 23137 11655 23171
rect 12633 23137 12667 23171
rect 18429 23137 18463 23171
rect 19441 23137 19475 23171
rect 22385 23137 22419 23171
rect 23305 23137 23339 23171
rect 24961 23137 24995 23171
rect 25973 23137 26007 23171
rect 2053 23069 2087 23103
rect 2881 23069 2915 23103
rect 4169 23069 4203 23103
rect 5273 23069 5307 23103
rect 5733 23069 5767 23103
rect 6745 23069 6779 23103
rect 7665 23069 7699 23103
rect 7757 23069 7791 23103
rect 8033 23069 8067 23103
rect 8125 23069 8159 23103
rect 9321 23069 9355 23103
rect 9413 23069 9447 23103
rect 9505 23069 9539 23103
rect 9689 23069 9723 23103
rect 11069 23069 11103 23103
rect 11529 23069 11563 23103
rect 11713 23069 11747 23103
rect 12357 23069 12391 23103
rect 12449 23069 12483 23103
rect 12541 23069 12575 23103
rect 13369 23069 13403 23103
rect 13553 23069 13587 23103
rect 14381 23069 14415 23103
rect 15393 23069 15427 23103
rect 15577 23069 15611 23103
rect 15669 23069 15703 23103
rect 16589 23069 16623 23103
rect 18337 23069 18371 23103
rect 18521 23069 18555 23103
rect 19533 23069 19567 23103
rect 20729 23069 20763 23103
rect 20913 23069 20947 23103
rect 21005 23069 21039 23103
rect 21649 23069 21683 23103
rect 21833 23069 21867 23103
rect 22569 23069 22603 23103
rect 23489 23069 23523 23103
rect 24777 23069 24811 23103
rect 4997 23001 5031 23035
rect 5181 23001 5215 23035
rect 7849 23001 7883 23035
rect 10241 23001 10275 23035
rect 14105 23001 14139 23035
rect 17601 23001 17635 23035
rect 19257 23001 19291 23035
rect 22293 23001 22327 23035
rect 23213 23001 23247 23035
rect 26240 23001 26274 23035
rect 1869 22933 1903 22967
rect 2421 22933 2455 22967
rect 2973 22933 3007 22967
rect 3801 22933 3835 22967
rect 4261 22933 4295 22967
rect 5273 22933 5307 22967
rect 10885 22933 10919 22967
rect 13553 22933 13587 22967
rect 14289 22933 14323 22967
rect 14473 22933 14507 22967
rect 21189 22933 21223 22967
rect 21741 22933 21775 22967
rect 24869 22933 24903 22967
rect 27353 22933 27387 22967
rect 1777 22729 1811 22763
rect 2881 22729 2915 22763
rect 3525 22729 3559 22763
rect 4905 22729 4939 22763
rect 7849 22729 7883 22763
rect 10149 22729 10183 22763
rect 16037 22729 16071 22763
rect 19993 22729 20027 22763
rect 25513 22729 25547 22763
rect 27353 22729 27387 22763
rect 4261 22661 4295 22695
rect 6469 22661 6503 22695
rect 15117 22661 15151 22695
rect 15301 22661 15335 22695
rect 25605 22661 25639 22695
rect 1961 22593 1995 22627
rect 2789 22593 2823 22627
rect 3433 22593 3467 22627
rect 4077 22593 4111 22627
rect 5089 22593 5123 22627
rect 5181 22593 5215 22627
rect 5457 22593 5491 22627
rect 7113 22593 7147 22627
rect 7297 22593 7331 22627
rect 7757 22593 7791 22627
rect 8861 22593 8895 22627
rect 9045 22593 9079 22627
rect 9597 22593 9631 22627
rect 9781 22593 9815 22627
rect 9873 22593 9907 22627
rect 9965 22593 9999 22627
rect 10609 22593 10643 22627
rect 10793 22593 10827 22627
rect 12265 22593 12299 22627
rect 12357 22593 12391 22627
rect 14105 22593 14139 22627
rect 14197 22593 14231 22627
rect 15761 22593 15795 22627
rect 16037 22593 16071 22627
rect 16865 22593 16899 22627
rect 18337 22593 18371 22627
rect 18797 22593 18831 22627
rect 19625 22593 19659 22627
rect 20729 22593 20763 22627
rect 23673 22593 23707 22627
rect 27169 22593 27203 22627
rect 9137 22525 9171 22559
rect 12173 22525 12207 22559
rect 12449 22525 12483 22559
rect 13001 22525 13035 22559
rect 16957 22525 16991 22559
rect 18889 22525 18923 22559
rect 19717 22525 19751 22559
rect 20453 22525 20487 22559
rect 22201 22525 22235 22559
rect 22477 22525 22511 22559
rect 23949 22525 23983 22559
rect 25789 22525 25823 22559
rect 26985 22525 27019 22559
rect 10701 22457 10735 22491
rect 11989 22457 12023 22491
rect 13277 22457 13311 22491
rect 13461 22457 13495 22491
rect 18153 22457 18187 22491
rect 19165 22457 19199 22491
rect 2329 22389 2363 22423
rect 4445 22389 4479 22423
rect 5365 22389 5399 22423
rect 6561 22389 6595 22423
rect 7113 22389 7147 22423
rect 8677 22389 8711 22423
rect 14381 22389 14415 22423
rect 17141 22389 17175 22423
rect 18981 22389 19015 22423
rect 19625 22389 19659 22423
rect 25145 22389 25179 22423
rect 5089 22185 5123 22219
rect 8309 22185 8343 22219
rect 9137 22185 9171 22219
rect 11621 22185 11655 22219
rect 26249 22185 26283 22219
rect 4537 22117 4571 22151
rect 7941 22117 7975 22151
rect 9045 22117 9079 22151
rect 18153 22117 18187 22151
rect 7205 22049 7239 22083
rect 9229 22049 9263 22083
rect 9965 22049 9999 22083
rect 10057 22049 10091 22083
rect 10425 22049 10459 22083
rect 11897 22049 11931 22083
rect 12265 22049 12299 22083
rect 15853 22049 15887 22083
rect 16589 22049 16623 22083
rect 17693 22049 17727 22083
rect 20177 22049 20211 22083
rect 21925 22049 21959 22083
rect 23673 22049 23707 22083
rect 25053 22049 25087 22083
rect 26709 22049 26743 22083
rect 27077 22049 27111 22083
rect 1961 21981 1995 22015
rect 2605 21981 2639 22015
rect 3341 21981 3375 22015
rect 3617 21981 3651 22015
rect 4261 21981 4295 22015
rect 4353 21981 4387 22015
rect 4629 21981 4663 22015
rect 5089 21981 5123 22015
rect 5181 21981 5215 22015
rect 5365 21981 5399 22015
rect 5549 21981 5583 22015
rect 6837 21981 6871 22015
rect 6929 21981 6963 22015
rect 8125 21981 8159 22015
rect 8401 21981 8435 22015
rect 8953 21981 8987 22015
rect 9689 21981 9723 22015
rect 9873 21981 9907 22015
rect 10241 21981 10275 22015
rect 11805 21981 11839 22015
rect 12173 21981 12207 22015
rect 12725 21981 12759 22015
rect 12909 21981 12943 22015
rect 13553 21981 13587 22015
rect 14197 21981 14231 22015
rect 14381 21981 14415 22015
rect 17785 21981 17819 22015
rect 19257 21981 19291 22015
rect 19441 21981 19475 22015
rect 19901 21981 19935 22015
rect 21649 21981 21683 22015
rect 25697 21981 25731 22015
rect 25881 21981 25915 22015
rect 26065 21981 26099 22015
rect 26893 21981 26927 22015
rect 5457 21913 5491 21947
rect 7297 21913 7331 21947
rect 10977 21913 11011 21947
rect 14289 21913 14323 21947
rect 14933 21913 14967 21947
rect 15669 21913 15703 21947
rect 16405 21913 16439 21947
rect 23489 21913 23523 21947
rect 25973 21913 26007 21947
rect 1777 21845 1811 21879
rect 2421 21845 2455 21879
rect 2973 21845 3007 21879
rect 3433 21845 3467 21879
rect 4077 21845 4111 21879
rect 6653 21845 6687 21879
rect 11069 21845 11103 21879
rect 12081 21845 12115 21879
rect 12817 21845 12851 21879
rect 13369 21845 13403 21879
rect 15025 21845 15059 21879
rect 19441 21845 19475 21879
rect 23121 21845 23155 21879
rect 23581 21845 23615 21879
rect 24501 21845 24535 21879
rect 24869 21845 24903 21879
rect 24961 21845 24995 21879
rect 1501 21641 1535 21675
rect 4077 21641 4111 21675
rect 5457 21641 5491 21675
rect 7665 21641 7699 21675
rect 10701 21641 10735 21675
rect 10793 21641 10827 21675
rect 10977 21641 11011 21675
rect 11529 21641 11563 21675
rect 18337 21641 18371 21675
rect 19993 21641 20027 21675
rect 21281 21641 21315 21675
rect 25697 21641 25731 21675
rect 26341 21641 26375 21675
rect 3801 21573 3835 21607
rect 5181 21573 5215 21607
rect 13338 21573 13372 21607
rect 17141 21573 17175 21607
rect 20821 21573 20855 21607
rect 22017 21573 22051 21607
rect 23489 21573 23523 21607
rect 23581 21573 23615 21607
rect 25329 21573 25363 21607
rect 25421 21573 25455 21607
rect 1685 21505 1719 21539
rect 3065 21505 3099 21539
rect 3525 21505 3559 21539
rect 3709 21505 3743 21539
rect 3893 21505 3927 21539
rect 4905 21505 4939 21539
rect 5089 21505 5123 21539
rect 5273 21505 5307 21539
rect 6745 21505 6779 21539
rect 6837 21505 6871 21539
rect 7021 21505 7055 21539
rect 7113 21505 7147 21539
rect 7941 21505 7975 21539
rect 8125 21505 8159 21539
rect 8217 21505 8251 21539
rect 8401 21505 8435 21539
rect 9413 21505 9447 21539
rect 9781 21505 9815 21539
rect 9965 21505 9999 21539
rect 10609 21505 10643 21539
rect 13093 21505 13127 21539
rect 14933 21505 14967 21539
rect 15117 21505 15151 21539
rect 15945 21505 15979 21539
rect 16129 21505 16163 21539
rect 17969 21505 18003 21539
rect 18889 21505 18923 21539
rect 19533 21505 19567 21539
rect 19802 21505 19836 21539
rect 21097 21505 21131 21539
rect 22201 21505 22235 21539
rect 22293 21505 22327 21539
rect 23305 21505 23339 21539
rect 23673 21505 23707 21539
rect 24409 21505 24443 21539
rect 25145 21505 25179 21539
rect 25513 21505 25547 21539
rect 26249 21505 26283 21539
rect 26985 21505 27019 21539
rect 27169 21505 27203 21539
rect 2605 21437 2639 21471
rect 9571 21437 9605 21471
rect 10977 21437 11011 21471
rect 11713 21437 11747 21471
rect 11805 21437 11839 21471
rect 11897 21437 11931 21471
rect 11989 21437 12023 21471
rect 15025 21437 15059 21471
rect 17877 21437 17911 21471
rect 19625 21437 19659 21471
rect 20913 21437 20947 21471
rect 2881 21369 2915 21403
rect 6561 21369 6595 21403
rect 16037 21369 16071 21403
rect 22477 21369 22511 21403
rect 24593 21369 24627 21403
rect 2053 21301 2087 21335
rect 8033 21301 8067 21335
rect 9781 21301 9815 21335
rect 14473 21301 14507 21335
rect 17233 21301 17267 21335
rect 18981 21301 19015 21335
rect 19809 21301 19843 21335
rect 20913 21301 20947 21335
rect 22017 21301 22051 21335
rect 23857 21301 23891 21335
rect 26985 21301 27019 21335
rect 2421 21097 2455 21131
rect 5733 21097 5767 21131
rect 7665 21097 7699 21131
rect 7849 21097 7883 21131
rect 9965 21097 9999 21131
rect 10701 21097 10735 21131
rect 14289 21097 14323 21131
rect 16865 21097 16899 21131
rect 22385 21097 22419 21131
rect 23765 21097 23799 21131
rect 3433 21029 3467 21063
rect 10149 21029 10183 21063
rect 10977 21029 11011 21063
rect 22385 20961 22419 20995
rect 23397 20961 23431 20995
rect 25329 20961 25363 20995
rect 25973 20961 26007 20995
rect 1961 20893 1995 20927
rect 2329 20893 2363 20927
rect 2605 20893 2639 20927
rect 2973 20893 3007 20927
rect 3617 20893 3651 20927
rect 3985 20893 4019 20927
rect 4629 20893 4663 20927
rect 5181 20893 5215 20927
rect 5549 20893 5583 20927
rect 6653 20893 6687 20927
rect 6745 20893 6779 20927
rect 6837 20893 6871 20927
rect 7481 20893 7515 20927
rect 7665 20893 7699 20927
rect 8953 20893 8987 20927
rect 9137 20893 9171 20927
rect 9597 20893 9631 20927
rect 9965 20893 9999 20927
rect 10609 20893 10643 20927
rect 10793 20893 10827 20927
rect 11437 20893 11471 20927
rect 11621 20893 11655 20927
rect 12081 20893 12115 20927
rect 14105 20893 14139 20927
rect 15025 20893 15059 20927
rect 15485 20893 15519 20927
rect 17785 20893 17819 20927
rect 18521 20893 18555 20927
rect 19809 20893 19843 20927
rect 19901 20893 19935 20927
rect 20085 20893 20119 20927
rect 20177 20893 20211 20927
rect 20821 20893 20855 20927
rect 20913 20893 20947 20927
rect 21097 20893 21131 20927
rect 21189 20893 21223 20927
rect 21833 20893 21867 20927
rect 22293 20893 22327 20927
rect 22569 20893 22603 20927
rect 23581 20893 23615 20927
rect 26229 20893 26263 20927
rect 12326 20825 12360 20859
rect 15730 20825 15764 20859
rect 18705 20825 18739 20859
rect 25237 20825 25271 20859
rect 1777 20757 1811 20791
rect 2145 20757 2179 20791
rect 3249 20757 3283 20791
rect 3801 20757 3835 20791
rect 5365 20757 5399 20791
rect 7021 20757 7055 20791
rect 9137 20757 9171 20791
rect 11529 20757 11563 20791
rect 13461 20757 13495 20791
rect 14841 20757 14875 20791
rect 17877 20757 17911 20791
rect 19625 20757 19659 20791
rect 20637 20757 20671 20791
rect 21649 20757 21683 20791
rect 22753 20757 22787 20791
rect 24777 20757 24811 20791
rect 25145 20757 25179 20791
rect 27353 20757 27387 20791
rect 6929 20553 6963 20587
rect 13461 20553 13495 20587
rect 21281 20553 21315 20587
rect 23045 20553 23079 20587
rect 23213 20553 23247 20587
rect 24041 20553 24075 20587
rect 27353 20553 27387 20587
rect 13093 20485 13127 20519
rect 13309 20485 13343 20519
rect 20913 20485 20947 20519
rect 21129 20485 21163 20519
rect 22845 20485 22879 20519
rect 25513 20485 25547 20519
rect 1777 20417 1811 20451
rect 2145 20417 2179 20451
rect 2605 20417 2639 20451
rect 3617 20417 3651 20451
rect 4169 20417 4203 20451
rect 4905 20417 4939 20451
rect 5089 20417 5123 20451
rect 5365 20417 5399 20451
rect 6377 20417 6411 20451
rect 6745 20417 6779 20451
rect 7665 20417 7699 20451
rect 7941 20417 7975 20451
rect 9413 20417 9447 20451
rect 9781 20417 9815 20451
rect 10793 20417 10827 20451
rect 12173 20417 12207 20451
rect 12265 20417 12299 20451
rect 12362 20417 12396 20451
rect 12541 20417 12575 20451
rect 13921 20417 13955 20451
rect 14188 20417 14222 20451
rect 15945 20417 15979 20451
rect 16911 20417 16945 20451
rect 17049 20417 17083 20451
rect 17141 20417 17175 20451
rect 17325 20417 17359 20451
rect 18052 20417 18086 20451
rect 19625 20417 19659 20451
rect 19901 20417 19935 20451
rect 22017 20417 22051 20451
rect 22109 20417 22143 20451
rect 22293 20417 22327 20451
rect 22385 20417 22419 20451
rect 25329 20417 25363 20451
rect 25605 20417 25639 20451
rect 25697 20417 25731 20451
rect 27169 20417 27203 20451
rect 11897 20349 11931 20383
rect 17785 20349 17819 20383
rect 24133 20349 24167 20383
rect 24225 20349 24259 20383
rect 26985 20349 27019 20383
rect 4997 20281 5031 20315
rect 9965 20281 9999 20315
rect 10977 20281 11011 20315
rect 15301 20281 15335 20315
rect 25881 20281 25915 20315
rect 1593 20213 1627 20247
rect 2421 20213 2455 20247
rect 3433 20213 3467 20247
rect 4261 20213 4295 20247
rect 6653 20213 6687 20247
rect 9505 20213 9539 20247
rect 13277 20213 13311 20247
rect 15761 20213 15795 20247
rect 16681 20213 16715 20247
rect 19165 20213 19199 20247
rect 21097 20213 21131 20247
rect 21833 20213 21867 20247
rect 23029 20213 23063 20247
rect 23673 20213 23707 20247
rect 5273 20009 5307 20043
rect 6193 20009 6227 20043
rect 14105 20009 14139 20043
rect 15209 20009 15243 20043
rect 18153 20009 18187 20043
rect 19901 20009 19935 20043
rect 21373 20009 21407 20043
rect 22201 20009 22235 20043
rect 23857 20009 23891 20043
rect 1685 19941 1719 19975
rect 4445 19941 4479 19975
rect 2237 19873 2271 19907
rect 6745 19873 6779 19907
rect 12449 19873 12483 19907
rect 14381 19873 14415 19907
rect 18521 19873 18555 19907
rect 23489 19873 23523 19907
rect 25329 19873 25363 19907
rect 25973 19873 26007 19907
rect 1869 19805 1903 19839
rect 2513 19805 2547 19839
rect 3249 19805 3283 19839
rect 4997 19805 5031 19839
rect 5181 19805 5215 19839
rect 5365 19805 5399 19839
rect 6101 19805 6135 19839
rect 7021 19805 7055 19839
rect 8125 19805 8159 19839
rect 9229 19805 9263 19839
rect 9321 19805 9355 19839
rect 9413 19805 9447 19839
rect 9597 19805 9631 19839
rect 10333 19805 10367 19839
rect 12265 19805 12299 19839
rect 12357 19805 12391 19839
rect 12633 19805 12667 19839
rect 13369 19805 13403 19839
rect 14289 19805 14323 19839
rect 14473 19805 14507 19839
rect 14565 19805 14599 19839
rect 15485 19805 15519 19839
rect 15577 19805 15611 19839
rect 15669 19805 15703 19839
rect 15853 19805 15887 19839
rect 16313 19805 16347 19839
rect 16580 19805 16614 19839
rect 18337 19805 18371 19839
rect 18613 19805 18647 19839
rect 19257 19805 19291 19839
rect 19441 19805 19475 19839
rect 20177 19805 20211 19839
rect 20269 19805 20303 19839
rect 20361 19805 20395 19839
rect 20545 19805 20579 19839
rect 22477 19805 22511 19839
rect 22569 19805 22603 19839
rect 22661 19805 22695 19839
rect 22845 19805 22879 19839
rect 23673 19805 23707 19839
rect 26240 19805 26274 19839
rect 4261 19737 4295 19771
rect 8309 19737 8343 19771
rect 10600 19737 10634 19771
rect 13185 19737 13219 19771
rect 21189 19737 21223 19771
rect 2329 19669 2363 19703
rect 3065 19669 3099 19703
rect 8953 19669 8987 19703
rect 11713 19669 11747 19703
rect 12541 19669 12575 19703
rect 17693 19669 17727 19703
rect 19441 19669 19475 19703
rect 21389 19669 21423 19703
rect 21557 19669 21591 19703
rect 24777 19669 24811 19703
rect 25145 19669 25179 19703
rect 25237 19669 25271 19703
rect 27353 19669 27387 19703
rect 1685 19465 1719 19499
rect 4997 19465 5031 19499
rect 6929 19465 6963 19499
rect 13553 19465 13587 19499
rect 16129 19465 16163 19499
rect 16773 19465 16807 19499
rect 18153 19465 18187 19499
rect 22293 19465 22327 19499
rect 23305 19465 23339 19499
rect 25697 19465 25731 19499
rect 26249 19465 26283 19499
rect 27353 19465 27387 19499
rect 3884 19397 3918 19431
rect 10701 19397 10735 19431
rect 20177 19397 20211 19431
rect 21097 19397 21131 19431
rect 24133 19397 24167 19431
rect 25329 19397 25363 19431
rect 1869 19329 1903 19363
rect 2329 19329 2363 19363
rect 2513 19329 2547 19363
rect 2973 19329 3007 19363
rect 3157 19329 3191 19363
rect 3617 19329 3651 19363
rect 5549 19329 5583 19363
rect 6837 19329 6871 19363
rect 7941 19329 7975 19363
rect 8033 19329 8067 19363
rect 8125 19329 8159 19363
rect 8309 19329 8343 19363
rect 8769 19329 8803 19363
rect 9036 19329 9070 19363
rect 11759 19329 11793 19363
rect 11897 19329 11931 19363
rect 11989 19329 12023 19363
rect 12173 19329 12207 19363
rect 12633 19329 12667 19363
rect 12817 19329 12851 19363
rect 13809 19329 13843 19363
rect 13918 19329 13952 19363
rect 14013 19329 14047 19363
rect 14197 19329 14231 19363
rect 14749 19329 14783 19363
rect 15005 19329 15039 19363
rect 16681 19329 16715 19363
rect 17417 19329 17451 19363
rect 17601 19329 17635 19363
rect 17969 19329 18003 19363
rect 18889 19329 18923 19363
rect 19073 19329 19107 19363
rect 19257 19329 19291 19363
rect 19441 19329 19475 19363
rect 22477 19329 22511 19363
rect 22569 19329 22603 19363
rect 22753 19329 22787 19363
rect 22845 19329 22879 19363
rect 23489 19329 23523 19363
rect 23949 19329 23983 19363
rect 24225 19329 24259 19363
rect 24317 19329 24351 19363
rect 25145 19329 25179 19363
rect 25421 19329 25455 19363
rect 25513 19329 25547 19363
rect 26433 19329 26467 19363
rect 27169 19329 27203 19363
rect 13001 19261 13035 19295
rect 17693 19261 17727 19295
rect 17785 19261 17819 19295
rect 19165 19261 19199 19295
rect 21281 19261 21315 19295
rect 26985 19261 27019 19295
rect 2421 19125 2455 19159
rect 2973 19125 3007 19159
rect 5641 19125 5675 19159
rect 7665 19125 7699 19159
rect 10149 19125 10183 19159
rect 10793 19125 10827 19159
rect 11529 19125 11563 19159
rect 19625 19125 19659 19159
rect 20269 19125 20303 19159
rect 24501 19125 24535 19159
rect 1593 18921 1627 18955
rect 4905 18921 4939 18955
rect 9781 18921 9815 18955
rect 13553 18921 13587 18955
rect 21925 18921 21959 18955
rect 27261 18921 27295 18955
rect 2421 18853 2455 18887
rect 6837 18853 6871 18887
rect 10885 18853 10919 18887
rect 15761 18853 15795 18887
rect 18521 18853 18555 18887
rect 7573 18785 7607 18819
rect 9321 18785 9355 18819
rect 12449 18785 12483 18819
rect 14381 18785 14415 18819
rect 15669 18785 15703 18819
rect 18061 18785 18095 18819
rect 18153 18785 18187 18819
rect 22477 18785 22511 18819
rect 23581 18785 23615 18819
rect 1593 18717 1627 18751
rect 1777 18717 1811 18751
rect 2145 18717 2179 18751
rect 2605 18717 2639 18751
rect 3249 18717 3283 18751
rect 4261 18717 4295 18751
rect 4813 18717 4847 18751
rect 5457 18717 5491 18751
rect 7297 18717 7331 18751
rect 10011 18717 10045 18751
rect 10146 18717 10180 18751
rect 10241 18717 10275 18751
rect 10425 18717 10459 18751
rect 11161 18717 11195 18751
rect 11250 18714 11284 18748
rect 11366 18717 11400 18751
rect 11529 18717 11563 18751
rect 11989 18717 12023 18751
rect 12173 18717 12207 18751
rect 12541 18717 12575 18751
rect 13185 18717 13219 18751
rect 14105 18717 14139 18751
rect 15577 18717 15611 18751
rect 15853 18717 15887 18751
rect 16497 18717 16531 18751
rect 16773 18717 16807 18751
rect 17785 18717 17819 18751
rect 17969 18717 18003 18751
rect 18337 18717 18371 18751
rect 19257 18717 19291 18751
rect 19513 18717 19547 18751
rect 21281 18717 21315 18751
rect 23305 18717 23339 18751
rect 23489 18717 23523 18751
rect 24777 18717 24811 18751
rect 27077 18717 27111 18751
rect 5724 18649 5758 18683
rect 9137 18649 9171 18683
rect 13369 18649 13403 18683
rect 25044 18649 25078 18683
rect 2881 18581 2915 18615
rect 3065 18581 3099 18615
rect 4077 18581 4111 18615
rect 15393 18581 15427 18615
rect 20637 18581 20671 18615
rect 21097 18581 21131 18615
rect 22293 18581 22327 18615
rect 22385 18581 22419 18615
rect 23121 18581 23155 18615
rect 26157 18581 26191 18615
rect 7757 18377 7791 18411
rect 8309 18377 8343 18411
rect 11989 18377 12023 18411
rect 14749 18377 14783 18411
rect 16037 18377 16071 18411
rect 19441 18377 19475 18411
rect 20545 18377 20579 18411
rect 21005 18377 21039 18411
rect 21833 18377 21867 18411
rect 22201 18377 22235 18411
rect 4905 18309 4939 18343
rect 5549 18309 5583 18343
rect 12091 18309 12125 18343
rect 23296 18309 23330 18343
rect 25320 18309 25354 18343
rect 2228 18241 2262 18275
rect 4077 18241 4111 18275
rect 4537 18241 4571 18275
rect 4721 18241 4755 18275
rect 5365 18241 5399 18275
rect 6633 18241 6667 18275
rect 8217 18241 8251 18275
rect 9505 18241 9539 18275
rect 10701 18241 10735 18275
rect 10885 18241 10919 18275
rect 10977 18241 11011 18275
rect 11805 18241 11839 18275
rect 12725 18241 12759 18275
rect 12909 18241 12943 18275
rect 14105 18241 14139 18275
rect 14289 18241 14323 18275
rect 14933 18241 14967 18275
rect 15117 18241 15151 18275
rect 15209 18241 15243 18275
rect 15669 18241 15703 18275
rect 15853 18241 15887 18275
rect 17969 18241 18003 18275
rect 18153 18241 18187 18275
rect 18337 18241 18371 18275
rect 18532 18241 18566 18275
rect 19625 18241 19659 18275
rect 19809 18241 19843 18275
rect 20913 18241 20947 18275
rect 26985 18241 27019 18275
rect 27169 18241 27203 18275
rect 1961 18173 1995 18207
rect 6377 18173 6411 18207
rect 9229 18173 9263 18207
rect 13001 18173 13035 18207
rect 16681 18173 16715 18207
rect 16957 18173 16991 18207
rect 18245 18173 18279 18207
rect 19901 18173 19935 18207
rect 21097 18173 21131 18207
rect 22293 18173 22327 18207
rect 22385 18173 22419 18207
rect 23029 18173 23063 18207
rect 25053 18173 25087 18207
rect 3341 18105 3375 18139
rect 10701 18105 10735 18139
rect 3893 18037 3927 18071
rect 5733 18037 5767 18071
rect 11621 18037 11655 18071
rect 12541 18037 12575 18071
rect 18705 18037 18739 18071
rect 24409 18037 24443 18071
rect 26433 18037 26467 18071
rect 26985 18037 27019 18071
rect 6469 17833 6503 17867
rect 13001 17833 13035 17867
rect 16313 17833 16347 17867
rect 23397 17833 23431 17867
rect 15485 17765 15519 17799
rect 3801 17697 3835 17731
rect 7573 17697 7607 17731
rect 19717 17697 19751 17731
rect 21005 17697 21039 17731
rect 26709 17697 26743 17731
rect 1869 17629 1903 17663
rect 4057 17629 4091 17663
rect 5825 17629 5859 17663
rect 6745 17629 6779 17663
rect 6837 17629 6871 17663
rect 6929 17629 6963 17663
rect 7113 17629 7147 17663
rect 7849 17629 7883 17663
rect 9505 17629 9539 17663
rect 11621 17629 11655 17663
rect 14105 17629 14139 17663
rect 17325 17629 17359 17663
rect 19441 17629 19475 17663
rect 20729 17607 20763 17641
rect 20913 17629 20947 17663
rect 21097 17629 21131 17663
rect 21281 17629 21315 17663
rect 22017 17629 22051 17663
rect 24409 17629 24443 17663
rect 26433 17629 26467 17663
rect 26617 17629 26651 17663
rect 27353 17629 27387 17663
rect 2136 17561 2170 17595
rect 5641 17561 5675 17595
rect 9750 17561 9784 17595
rect 11888 17561 11922 17595
rect 14350 17561 14384 17595
rect 15945 17561 15979 17595
rect 16129 17561 16163 17595
rect 17592 17561 17626 17595
rect 22284 17561 22318 17595
rect 24654 17561 24688 17595
rect 3249 17493 3283 17527
rect 5181 17493 5215 17527
rect 6009 17493 6043 17527
rect 10885 17493 10919 17527
rect 18705 17493 18739 17527
rect 21465 17493 21499 17527
rect 25789 17493 25823 17527
rect 26249 17493 26283 17527
rect 27169 17493 27203 17527
rect 3893 17289 3927 17323
rect 9597 17289 9631 17323
rect 10885 17289 10919 17323
rect 13001 17289 13035 17323
rect 13737 17289 13771 17323
rect 17601 17289 17635 17323
rect 24225 17289 24259 17323
rect 2228 17221 2262 17255
rect 4721 17221 4755 17255
rect 5549 17221 5583 17255
rect 14933 17221 14967 17255
rect 18797 17221 18831 17255
rect 25697 17221 25731 17255
rect 27077 17221 27111 17255
rect 4077 17153 4111 17187
rect 4537 17153 4571 17187
rect 5365 17153 5399 17187
rect 5733 17153 5767 17187
rect 6633 17153 6667 17187
rect 8309 17153 8343 17187
rect 9873 17153 9907 17187
rect 9965 17153 9999 17187
rect 10057 17153 10091 17187
rect 10241 17153 10275 17187
rect 10793 17153 10827 17187
rect 11713 17153 11747 17187
rect 11989 17153 12023 17187
rect 12173 17153 12207 17187
rect 12817 17153 12851 17187
rect 13093 17153 13127 17187
rect 13993 17153 14027 17187
rect 14105 17153 14139 17187
rect 14197 17153 14231 17187
rect 14381 17153 14415 17187
rect 15117 17153 15151 17187
rect 15853 17153 15887 17187
rect 15945 17153 15979 17187
rect 16865 17153 16899 17187
rect 17785 17153 17819 17187
rect 18613 17153 18647 17187
rect 19625 17153 19659 17187
rect 21837 17153 21871 17187
rect 22017 17153 22051 17187
rect 22201 17153 22235 17187
rect 22385 17153 22419 17187
rect 23029 17153 23063 17187
rect 23213 17153 23247 17187
rect 23305 17153 23339 17187
rect 23581 17153 23615 17187
rect 23765 17153 23799 17187
rect 24409 17153 24443 17187
rect 24685 17153 24719 17187
rect 25881 17153 25915 17187
rect 1961 17085 1995 17119
rect 6377 17085 6411 17119
rect 8585 17085 8619 17119
rect 12633 17085 12667 17119
rect 15301 17085 15335 17119
rect 16681 17085 16715 17119
rect 18061 17085 18095 17119
rect 19717 17085 19751 17119
rect 19901 17085 19935 17119
rect 20453 17085 20487 17119
rect 22109 17085 22143 17119
rect 23397 17085 23431 17119
rect 24593 17085 24627 17119
rect 26065 17085 26099 17119
rect 26157 17085 26191 17119
rect 3341 17017 3375 17051
rect 11805 17017 11839 17051
rect 11897 17017 11931 17051
rect 17049 17017 17083 17051
rect 27261 17017 27295 17051
rect 4905 16949 4939 16983
rect 7757 16949 7791 16983
rect 11529 16949 11563 16983
rect 16129 16949 16163 16983
rect 17969 16949 18003 16983
rect 19257 16949 19291 16983
rect 20683 16949 20717 16983
rect 22569 16949 22603 16983
rect 4813 16745 4847 16779
rect 6285 16745 6319 16779
rect 10149 16745 10183 16779
rect 11989 16745 12023 16779
rect 18245 16745 18279 16779
rect 19809 16745 19843 16779
rect 21925 16745 21959 16779
rect 25145 16745 25179 16779
rect 13461 16677 13495 16711
rect 14749 16677 14783 16711
rect 15853 16677 15887 16711
rect 17877 16677 17911 16711
rect 7021 16609 7055 16643
rect 10609 16609 10643 16643
rect 16313 16609 16347 16643
rect 16681 16609 16715 16643
rect 17417 16609 17451 16643
rect 18337 16609 18371 16643
rect 21465 16609 21499 16643
rect 21557 16609 21591 16643
rect 22845 16609 22879 16643
rect 23121 16609 23155 16643
rect 24685 16609 24719 16643
rect 25973 16609 26007 16643
rect 1869 16541 1903 16575
rect 4353 16541 4387 16575
rect 4997 16541 5031 16575
rect 5641 16541 5675 16575
rect 6469 16541 6503 16575
rect 9137 16541 9171 16575
rect 12633 16541 12667 16575
rect 13093 16541 13127 16575
rect 14105 16541 14139 16575
rect 14198 16541 14232 16575
rect 14570 16541 14604 16575
rect 15209 16541 15243 16575
rect 15357 16541 15391 16575
rect 15674 16541 15708 16575
rect 16497 16541 16531 16575
rect 18061 16541 18095 16575
rect 20545 16541 20579 16575
rect 21189 16541 21223 16575
rect 21373 16541 21407 16575
rect 21741 16541 21775 16575
rect 24409 16541 24443 16575
rect 24593 16541 24627 16575
rect 24777 16541 24811 16575
rect 24961 16541 24995 16575
rect 26240 16541 26274 16575
rect 2136 16473 2170 16507
rect 7288 16473 7322 16507
rect 9781 16473 9815 16507
rect 9965 16473 9999 16507
rect 10876 16473 10910 16507
rect 14381 16473 14415 16507
rect 14473 16473 14507 16507
rect 15485 16473 15519 16507
rect 15577 16473 15611 16507
rect 17233 16473 17267 16507
rect 19717 16473 19751 16507
rect 3249 16405 3283 16439
rect 4169 16405 4203 16439
rect 5457 16405 5491 16439
rect 8401 16405 8435 16439
rect 8953 16405 8987 16439
rect 12449 16405 12483 16439
rect 13553 16405 13587 16439
rect 20361 16405 20395 16439
rect 27353 16405 27387 16439
rect 5457 16201 5491 16235
rect 7573 16201 7607 16235
rect 8401 16201 8435 16235
rect 25789 16201 25823 16235
rect 27261 16201 27295 16235
rect 7205 16133 7239 16167
rect 7421 16133 7455 16167
rect 8033 16133 8067 16167
rect 8249 16133 8283 16167
rect 9220 16133 9254 16167
rect 13645 16133 13679 16167
rect 2053 16065 2087 16099
rect 2513 16065 2547 16099
rect 2697 16065 2731 16099
rect 3525 16065 3559 16099
rect 4077 16065 4111 16099
rect 4344 16065 4378 16099
rect 6561 16065 6595 16099
rect 8953 16065 8987 16099
rect 10793 16065 10827 16099
rect 10977 16065 11011 16099
rect 12173 16065 12207 16099
rect 13277 16065 13311 16099
rect 13370 16065 13404 16099
rect 13553 16065 13587 16099
rect 13783 16065 13817 16099
rect 14381 16065 14415 16099
rect 16865 16065 16899 16099
rect 16957 16065 16991 16099
rect 17233 16065 17267 16099
rect 17969 16065 18003 16099
rect 18225 16065 18259 16099
rect 19809 16065 19843 16099
rect 20065 16065 20099 16099
rect 22192 16065 22226 16099
rect 24041 16065 24075 16099
rect 25053 16065 25087 16099
rect 25237 16065 25271 16099
rect 25329 16065 25363 16099
rect 25605 16065 25639 16099
rect 26433 16065 26467 16099
rect 27169 16065 27203 16099
rect 11897 15997 11931 16031
rect 16129 15997 16163 16031
rect 17141 15997 17175 16031
rect 21925 15997 21959 16031
rect 23765 15997 23799 16031
rect 25421 15997 25455 16031
rect 19349 15929 19383 15963
rect 1869 15861 1903 15895
rect 2881 15861 2915 15895
rect 3341 15861 3375 15895
rect 6377 15861 6411 15895
rect 7389 15861 7423 15895
rect 8217 15861 8251 15895
rect 10333 15861 10367 15895
rect 10793 15861 10827 15895
rect 13921 15861 13955 15895
rect 16681 15861 16715 15895
rect 21189 15861 21223 15895
rect 23305 15861 23339 15895
rect 26249 15861 26283 15895
rect 2789 15657 2823 15691
rect 4169 15657 4203 15691
rect 4997 15657 5031 15691
rect 5181 15657 5215 15691
rect 8217 15657 8251 15691
rect 10609 15657 10643 15691
rect 11805 15657 11839 15691
rect 16037 15657 16071 15691
rect 18153 15657 18187 15691
rect 19717 15657 19751 15691
rect 20821 15657 20855 15691
rect 23213 15657 23247 15691
rect 23581 15657 23615 15691
rect 27353 15657 27387 15691
rect 14105 15589 14139 15623
rect 15393 15589 15427 15623
rect 20085 15589 20119 15623
rect 1409 15521 1443 15555
rect 5641 15521 5675 15555
rect 8953 15521 8987 15555
rect 12725 15521 12759 15555
rect 21465 15521 21499 15555
rect 22385 15521 22419 15555
rect 23673 15521 23707 15555
rect 24409 15521 24443 15555
rect 24685 15521 24719 15555
rect 25973 15521 26007 15555
rect 4353 15453 4387 15487
rect 5908 15453 5942 15487
rect 9229 15453 9263 15487
rect 10241 15453 10275 15487
rect 11069 15453 11103 15487
rect 11161 15453 11195 15487
rect 11989 15453 12023 15487
rect 12449 15453 12483 15487
rect 14289 15453 14323 15487
rect 14749 15453 14783 15487
rect 14842 15453 14876 15487
rect 15025 15453 15059 15487
rect 15255 15453 15289 15487
rect 16773 15453 16807 15487
rect 19901 15453 19935 15487
rect 20177 15453 20211 15487
rect 21281 15453 21315 15487
rect 22017 15453 22051 15487
rect 22201 15453 22235 15487
rect 22293 15453 22327 15487
rect 22569 15453 22603 15487
rect 23397 15453 23431 15487
rect 16083 15419 16117 15453
rect 1676 15385 1710 15419
rect 4813 15385 4847 15419
rect 8125 15385 8159 15419
rect 10425 15385 10459 15419
rect 15117 15385 15151 15419
rect 15853 15385 15887 15419
rect 17040 15385 17074 15419
rect 26240 15385 26274 15419
rect 5023 15317 5057 15351
rect 7021 15317 7055 15351
rect 16221 15317 16255 15351
rect 21189 15317 21223 15351
rect 22753 15317 22787 15351
rect 1869 15113 1903 15147
rect 2513 15113 2547 15147
rect 5207 15113 5241 15147
rect 6577 15113 6611 15147
rect 6745 15113 6779 15147
rect 7481 15113 7515 15147
rect 8217 15113 8251 15147
rect 9137 15113 9171 15147
rect 10885 15113 10919 15147
rect 13119 15113 13153 15147
rect 14397 15113 14431 15147
rect 15869 15113 15903 15147
rect 16037 15113 16071 15147
rect 17141 15113 17175 15147
rect 19533 15113 19567 15147
rect 26249 15113 26283 15147
rect 4997 15045 5031 15079
rect 6377 15045 6411 15079
rect 9873 15045 9907 15079
rect 11529 15045 11563 15079
rect 11745 15045 11779 15079
rect 12909 15045 12943 15079
rect 14197 15045 14231 15079
rect 15669 15045 15703 15079
rect 20269 15045 20303 15079
rect 2053 14977 2087 15011
rect 2697 14961 2731 14995
rect 3424 14977 3458 15011
rect 7389 14977 7423 15011
rect 7573 14977 7607 15011
rect 8125 14977 8159 15011
rect 8769 14977 8803 15011
rect 10793 14977 10827 15011
rect 10977 14977 11011 15011
rect 15209 14977 15243 15011
rect 16773 14977 16807 15011
rect 16957 14977 16991 15011
rect 18153 14977 18187 15011
rect 18420 14977 18454 15011
rect 19993 14977 20027 15011
rect 20086 14977 20120 15011
rect 20361 14977 20395 15011
rect 20499 14977 20533 15011
rect 21281 14977 21315 15011
rect 22017 14977 22051 15011
rect 22293 14977 22327 15011
rect 23121 14977 23155 15011
rect 23213 14977 23247 15011
rect 25513 14977 25547 15011
rect 25697 14977 25731 15011
rect 26065 14977 26099 15011
rect 27169 14977 27203 15011
rect 3157 14909 3191 14943
rect 8861 14909 8895 14943
rect 23305 14909 23339 14943
rect 24225 14909 24259 14943
rect 24501 14909 24535 14943
rect 25789 14909 25823 14943
rect 25881 14909 25915 14943
rect 5365 14841 5399 14875
rect 11897 14841 11931 14875
rect 14565 14841 14599 14875
rect 22753 14841 22787 14875
rect 26985 14841 27019 14875
rect 4537 14773 4571 14807
rect 5181 14773 5215 14807
rect 6561 14773 6595 14807
rect 8953 14773 8987 14807
rect 9965 14773 9999 14807
rect 11713 14773 11747 14807
rect 13093 14773 13127 14807
rect 13277 14773 13311 14807
rect 14381 14773 14415 14807
rect 15025 14773 15059 14807
rect 15853 14773 15887 14807
rect 20637 14773 20671 14807
rect 21097 14773 21131 14807
rect 21833 14773 21867 14807
rect 22201 14773 22235 14807
rect 3801 14569 3835 14603
rect 8953 14569 8987 14603
rect 9965 14569 9999 14603
rect 12633 14569 12667 14603
rect 13277 14569 13311 14603
rect 15301 14569 15335 14603
rect 16129 14569 16163 14603
rect 22293 14569 22327 14603
rect 27353 14569 27387 14603
rect 11805 14501 11839 14535
rect 14565 14501 14599 14535
rect 6469 14433 6503 14467
rect 9045 14433 9079 14467
rect 10425 14433 10459 14467
rect 11069 14433 11103 14467
rect 22937 14433 22971 14467
rect 24409 14433 24443 14467
rect 25973 14433 26007 14467
rect 1409 14365 1443 14399
rect 3985 14365 4019 14399
rect 4629 14365 4663 14399
rect 5273 14365 5307 14399
rect 6009 14365 6043 14399
rect 9229 14365 9263 14399
rect 10149 14365 10183 14399
rect 10333 14365 10367 14399
rect 11253 14365 11287 14399
rect 11713 14365 11747 14399
rect 13461 14365 13495 14399
rect 14290 14365 14324 14399
rect 14382 14365 14416 14399
rect 14611 14365 14645 14399
rect 15945 14365 15979 14399
rect 17877 14365 17911 14399
rect 18061 14365 18095 14399
rect 20177 14365 20211 14399
rect 24685 14365 24719 14399
rect 26229 14365 26263 14399
rect 1676 14297 1710 14331
rect 6736 14297 6770 14331
rect 8953 14297 8987 14331
rect 12449 14297 12483 14331
rect 12649 14297 12683 14331
rect 14105 14297 14139 14331
rect 15117 14297 15151 14331
rect 15317 14297 15351 14331
rect 16773 14297 16807 14331
rect 19349 14297 19383 14331
rect 20422 14297 20456 14331
rect 22661 14297 22695 14331
rect 23673 14297 23707 14331
rect 23857 14297 23891 14331
rect 2789 14229 2823 14263
rect 4445 14229 4479 14263
rect 5089 14229 5123 14263
rect 5825 14229 5859 14263
rect 7849 14229 7883 14263
rect 9413 14229 9447 14263
rect 12817 14229 12851 14263
rect 15485 14229 15519 14263
rect 16865 14229 16899 14263
rect 18245 14229 18279 14263
rect 19441 14229 19475 14263
rect 21557 14229 21591 14263
rect 22753 14229 22787 14263
rect 1685 14025 1719 14059
rect 6745 14025 6779 14059
rect 9229 14025 9263 14059
rect 10793 14025 10827 14059
rect 12383 14025 12417 14059
rect 14473 14025 14507 14059
rect 15133 14025 15167 14059
rect 15301 14025 15335 14059
rect 19165 14025 19199 14059
rect 22017 14025 22051 14059
rect 26249 14025 26283 14059
rect 26985 14025 27019 14059
rect 4712 13957 4746 13991
rect 7941 13957 7975 13991
rect 8585 13957 8619 13991
rect 12173 13957 12207 13991
rect 14933 13957 14967 13991
rect 15761 13957 15795 13991
rect 15977 13957 16011 13991
rect 16948 13957 16982 13991
rect 19901 13957 19935 13991
rect 20913 13957 20947 13991
rect 21005 13957 21039 13991
rect 1869 13889 1903 13923
rect 2605 13889 2639 13923
rect 2872 13889 2906 13923
rect 6929 13889 6963 13923
rect 8732 13889 8766 13923
rect 9781 13889 9815 13923
rect 10517 13889 10551 13923
rect 11529 13889 11563 13923
rect 13360 13889 13394 13923
rect 18521 13889 18555 13923
rect 18669 13889 18703 13923
rect 18797 13889 18831 13923
rect 18889 13889 18923 13923
rect 19027 13889 19061 13923
rect 19717 13889 19751 13923
rect 20626 13889 20660 13923
rect 20730 13889 20764 13923
rect 21143 13889 21177 13923
rect 21833 13889 21867 13923
rect 22569 13889 22603 13923
rect 22753 13889 22787 13923
rect 23121 13889 23155 13923
rect 23305 13889 23339 13923
rect 23765 13889 23799 13923
rect 23937 13895 23971 13929
rect 24133 13889 24167 13923
rect 24317 13889 24351 13923
rect 24961 13889 24995 13923
rect 25145 13889 25179 13923
rect 25513 13889 25547 13923
rect 26433 13889 26467 13923
rect 27169 13889 27203 13923
rect 4445 13821 4479 13855
rect 8953 13821 8987 13855
rect 10057 13821 10091 13855
rect 10793 13821 10827 13855
rect 11621 13821 11655 13855
rect 13093 13821 13127 13855
rect 16681 13821 16715 13855
rect 22845 13821 22879 13855
rect 22937 13821 22971 13855
rect 24041 13821 24075 13855
rect 24501 13821 24535 13855
rect 25237 13821 25271 13855
rect 25329 13821 25363 13855
rect 8125 13753 8159 13787
rect 9873 13753 9907 13787
rect 10609 13753 10643 13787
rect 16129 13753 16163 13787
rect 20085 13753 20119 13787
rect 21281 13753 21315 13787
rect 3985 13685 4019 13719
rect 5825 13685 5859 13719
rect 8861 13685 8895 13719
rect 9965 13685 9999 13719
rect 12357 13685 12391 13719
rect 12541 13685 12575 13719
rect 15117 13685 15151 13719
rect 15945 13685 15979 13719
rect 18061 13685 18095 13719
rect 25697 13685 25731 13719
rect 5273 13481 5307 13515
rect 7297 13481 7331 13515
rect 8309 13481 8343 13515
rect 10701 13481 10735 13515
rect 17601 13481 17635 13515
rect 19901 13481 19935 13515
rect 27353 13481 27387 13515
rect 6745 13413 6779 13447
rect 4629 13345 4663 13379
rect 5365 13345 5399 13379
rect 11345 13345 11379 13379
rect 12173 13345 12207 13379
rect 14565 13345 14599 13379
rect 20913 13345 20947 13379
rect 25053 13345 25087 13379
rect 25145 13345 25179 13379
rect 1593 13277 1627 13311
rect 6653 13277 6687 13311
rect 6745 13277 6779 13311
rect 7205 13277 7239 13311
rect 8217 13277 8251 13311
rect 8401 13277 8435 13311
rect 8953 13277 8987 13311
rect 9229 13277 9263 13311
rect 11529 13277 11563 13311
rect 12449 13277 12483 13311
rect 14289 13277 14323 13311
rect 15577 13277 15611 13311
rect 15670 13277 15704 13311
rect 16042 13277 16076 13311
rect 16957 13277 16991 13311
rect 17105 13277 17139 13311
rect 17422 13277 17456 13311
rect 18061 13277 18095 13311
rect 18154 13277 18188 13311
rect 18429 13277 18463 13311
rect 18567 13277 18601 13311
rect 19257 13277 19291 13311
rect 19405 13277 19439 13311
rect 19633 13277 19667 13311
rect 19722 13277 19756 13311
rect 20637 13277 20671 13311
rect 22385 13277 22419 13311
rect 24777 13277 24811 13311
rect 24961 13277 24995 13311
rect 25329 13277 25363 13311
rect 25973 13277 26007 13311
rect 1860 13209 1894 13243
rect 4445 13209 4479 13243
rect 5089 13209 5123 13243
rect 5457 13209 5491 13243
rect 6469 13209 6503 13243
rect 10609 13209 10643 13243
rect 11713 13209 11747 13243
rect 15853 13209 15887 13243
rect 15945 13209 15979 13243
rect 17233 13209 17267 13243
rect 17325 13209 17359 13243
rect 18337 13209 18371 13243
rect 19533 13209 19567 13243
rect 22652 13209 22686 13243
rect 26240 13209 26274 13243
rect 2973 13141 3007 13175
rect 5181 13141 5215 13175
rect 7665 13141 7699 13175
rect 16221 13141 16255 13175
rect 18705 13141 18739 13175
rect 23765 13141 23799 13175
rect 25513 13141 25547 13175
rect 3065 12937 3099 12971
rect 6745 12937 6779 12971
rect 8309 12937 8343 12971
rect 9229 12937 9263 12971
rect 11713 12937 11747 12971
rect 13369 12937 13403 12971
rect 17785 12937 17819 12971
rect 19717 12937 19751 12971
rect 22477 12937 22511 12971
rect 22845 12937 22879 12971
rect 25053 12937 25087 12971
rect 2697 12869 2731 12903
rect 6653 12869 6687 12903
rect 10149 12869 10183 12903
rect 10241 12869 10275 12903
rect 14197 12869 14231 12903
rect 15117 12869 15151 12903
rect 18604 12869 18638 12903
rect 1777 12801 1811 12835
rect 1961 12801 1995 12835
rect 2881 12801 2915 12835
rect 3985 12801 4019 12835
rect 4252 12801 4286 12835
rect 7481 12801 7515 12835
rect 7941 12801 7975 12835
rect 8769 12801 8803 12835
rect 9085 12801 9119 12835
rect 10057 12801 10091 12835
rect 10379 12801 10413 12835
rect 11529 12801 11563 12835
rect 12265 12801 12299 12835
rect 12449 12801 12483 12835
rect 13277 12801 13311 12835
rect 14933 12801 14967 12835
rect 16129 12801 16163 12835
rect 17141 12801 17175 12835
rect 17693 12801 17727 12835
rect 20729 12801 20763 12835
rect 20913 12801 20947 12835
rect 21005 12801 21039 12835
rect 21097 12801 21131 12835
rect 22017 12801 22051 12835
rect 23673 12801 23707 12835
rect 23940 12801 23974 12835
rect 26157 12801 26191 12835
rect 27353 12801 27387 12835
rect 8033 12733 8067 12767
rect 8861 12733 8895 12767
rect 10517 12733 10551 12767
rect 13553 12733 13587 12767
rect 18337 12733 18371 12767
rect 22937 12733 22971 12767
rect 23121 12733 23155 12767
rect 26433 12733 26467 12767
rect 5365 12665 5399 12699
rect 14381 12665 14415 12699
rect 15945 12665 15979 12699
rect 25973 12665 26007 12699
rect 2145 12597 2179 12631
rect 7297 12597 7331 12631
rect 8125 12597 8159 12631
rect 8769 12597 8803 12631
rect 9873 12597 9907 12631
rect 12357 12597 12391 12631
rect 12909 12597 12943 12631
rect 16957 12597 16991 12631
rect 21281 12597 21315 12631
rect 21833 12597 21867 12631
rect 26341 12597 26375 12631
rect 27169 12597 27203 12631
rect 2053 12393 2087 12427
rect 2513 12393 2547 12427
rect 3801 12393 3835 12427
rect 7757 12393 7791 12427
rect 10333 12393 10367 12427
rect 13093 12393 13127 12427
rect 15669 12393 15703 12427
rect 17601 12393 17635 12427
rect 18429 12393 18463 12427
rect 21557 12393 21591 12427
rect 23305 12393 23339 12427
rect 25421 12393 25455 12427
rect 4261 12325 4295 12359
rect 9597 12325 9631 12359
rect 23673 12325 23707 12359
rect 7389 12257 7423 12291
rect 8309 12257 8343 12291
rect 11713 12257 11747 12291
rect 19717 12257 19751 12291
rect 23765 12257 23799 12291
rect 25513 12257 25547 12291
rect 25973 12257 26007 12291
rect 2697 12189 2731 12223
rect 3985 12189 4019 12223
rect 4077 12189 4111 12223
rect 4353 12189 4387 12223
rect 5365 12189 5399 12223
rect 5641 12189 5675 12223
rect 5733 12189 5767 12223
rect 6377 12189 6411 12223
rect 6653 12189 6687 12223
rect 6745 12189 6779 12223
rect 7573 12189 7607 12223
rect 8217 12189 8251 12223
rect 10517 12189 10551 12223
rect 10793 12189 10827 12223
rect 11980 12189 12014 12223
rect 14289 12189 14323 12223
rect 16221 12189 16255 12223
rect 18245 12189 18279 12223
rect 19349 12189 19383 12223
rect 20177 12189 20211 12223
rect 22063 12189 22097 12223
rect 22293 12189 22327 12223
rect 23489 12189 23523 12223
rect 24593 12189 24627 12223
rect 25237 12189 25271 12223
rect 26240 12189 26274 12223
rect 1685 12121 1719 12155
rect 1869 12121 1903 12155
rect 5549 12121 5583 12155
rect 6561 12121 6595 12155
rect 9413 12121 9447 12155
rect 10701 12121 10735 12155
rect 14534 12121 14568 12155
rect 16466 12121 16500 12155
rect 18061 12121 18095 12155
rect 19533 12121 19567 12155
rect 20444 12121 20478 12155
rect 5917 12053 5951 12087
rect 6929 12053 6963 12087
rect 24409 12053 24443 12087
rect 25053 12053 25087 12087
rect 27353 12053 27387 12087
rect 2789 11849 2823 11883
rect 3801 11849 3835 11883
rect 6745 11849 6779 11883
rect 9137 11849 9171 11883
rect 10977 11849 11011 11883
rect 12265 11849 12299 11883
rect 14489 11849 14523 11883
rect 14657 11849 14691 11883
rect 18613 11849 18647 11883
rect 24041 11849 24075 11883
rect 26433 11849 26467 11883
rect 5365 11781 5399 11815
rect 8002 11781 8036 11815
rect 11897 11781 11931 11815
rect 14289 11781 14323 11815
rect 15577 11781 15611 11815
rect 15793 11781 15827 11815
rect 18245 11781 18279 11815
rect 19533 11781 19567 11815
rect 2053 11713 2087 11747
rect 2973 11713 3007 11747
rect 3065 11713 3099 11747
rect 3341 11713 3375 11747
rect 3985 11713 4019 11747
rect 4077 11713 4111 11747
rect 4353 11713 4387 11747
rect 5089 11713 5123 11747
rect 5273 11713 5307 11747
rect 5457 11713 5491 11747
rect 6561 11713 6595 11747
rect 9853 11713 9887 11747
rect 12081 11713 12115 11747
rect 12725 11713 12759 11747
rect 13001 11713 13035 11747
rect 13553 11713 13587 11747
rect 16957 11713 16991 11747
rect 17233 11713 17267 11747
rect 18429 11713 18463 11747
rect 20913 11713 20947 11747
rect 21925 11713 21959 11747
rect 22109 11713 22143 11747
rect 22201 11713 22235 11747
rect 22293 11713 22327 11747
rect 23305 11713 23339 11747
rect 24225 11713 24259 11747
rect 25053 11713 25087 11747
rect 25309 11713 25343 11747
rect 27077 11713 27111 11747
rect 6377 11645 6411 11679
rect 7757 11645 7791 11679
rect 9597 11645 9631 11679
rect 19717 11645 19751 11679
rect 24501 11645 24535 11679
rect 3249 11577 3283 11611
rect 4261 11577 4295 11611
rect 13001 11577 13035 11611
rect 13737 11577 13771 11611
rect 15945 11577 15979 11611
rect 22477 11577 22511 11611
rect 27261 11577 27295 11611
rect 1869 11509 1903 11543
rect 5641 11509 5675 11543
rect 14473 11509 14507 11543
rect 15761 11509 15795 11543
rect 20729 11509 20763 11543
rect 23489 11509 23523 11543
rect 24409 11509 24443 11543
rect 6101 11305 6135 11339
rect 9321 11305 9355 11339
rect 9965 11305 9999 11339
rect 14473 11305 14507 11339
rect 18705 11305 18739 11339
rect 19809 11305 19843 11339
rect 21649 11305 21683 11339
rect 26341 11305 26375 11339
rect 7435 11237 7469 11271
rect 15393 11169 15427 11203
rect 16773 11169 16807 11203
rect 17325 11169 17359 11203
rect 22109 11169 22143 11203
rect 24501 11169 24535 11203
rect 26709 11169 26743 11203
rect 26801 11169 26835 11203
rect 1685 11101 1719 11135
rect 1952 11101 1986 11135
rect 3893 11101 3927 11135
rect 5733 11101 5767 11135
rect 5917 11101 5951 11135
rect 6745 11101 6779 11135
rect 7205 11101 7239 11135
rect 9045 11101 9079 11135
rect 9137 11101 9171 11135
rect 10609 11101 10643 11135
rect 11437 11101 11471 11135
rect 11621 11101 11655 11135
rect 11897 11101 11931 11135
rect 12725 11101 12759 11135
rect 13001 11101 13035 11135
rect 14105 11101 14139 11135
rect 14381 11101 14415 11135
rect 16497 11101 16531 11135
rect 16589 11101 16623 11135
rect 16865 11101 16899 11135
rect 20269 11101 20303 11135
rect 20525 11101 20559 11135
rect 24409 11101 24443 11135
rect 24961 11101 24995 11135
rect 25421 11101 25455 11135
rect 25605 11101 25639 11135
rect 26525 11101 26559 11135
rect 4160 11033 4194 11067
rect 9873 11033 9907 11067
rect 10793 11033 10827 11067
rect 15209 11033 15243 11067
rect 16313 11033 16347 11067
rect 17592 11033 17626 11067
rect 19441 11033 19475 11067
rect 19625 11033 19659 11067
rect 22376 11033 22410 11067
rect 3065 10965 3099 10999
rect 5273 10965 5307 10999
rect 6561 10965 6595 10999
rect 14657 10965 14691 10999
rect 23489 10965 23523 10999
rect 2237 10761 2271 10795
rect 8769 10761 8803 10795
rect 10793 10761 10827 10795
rect 12081 10761 12115 10795
rect 14841 10761 14875 10795
rect 21097 10761 21131 10795
rect 26341 10761 26375 10795
rect 1869 10693 1903 10727
rect 3065 10693 3099 10727
rect 5549 10693 5583 10727
rect 10609 10693 10643 10727
rect 16948 10693 16982 10727
rect 19984 10693 20018 10727
rect 25206 10693 25240 10727
rect 2053 10625 2087 10659
rect 3249 10625 3283 10659
rect 3341 10625 3375 10659
rect 3617 10625 3651 10659
rect 4537 10625 4571 10659
rect 4629 10625 4663 10659
rect 5273 10625 5307 10659
rect 5457 10625 5491 10659
rect 5641 10625 5675 10659
rect 6561 10625 6595 10659
rect 6828 10625 6862 10659
rect 8585 10625 8619 10659
rect 9873 10625 9907 10659
rect 10057 10625 10091 10659
rect 10885 10625 10919 10659
rect 11897 10625 11931 10659
rect 12173 10625 12207 10659
rect 12633 10625 12667 10659
rect 13728 10625 13762 10659
rect 15669 10625 15703 10659
rect 15853 10625 15887 10659
rect 15945 10625 15979 10659
rect 16681 10625 16715 10659
rect 19073 10625 19107 10659
rect 19717 10625 19751 10659
rect 22201 10625 22235 10659
rect 23029 10625 23063 10659
rect 23581 10625 23615 10659
rect 23857 10625 23891 10659
rect 24225 10625 24259 10659
rect 24961 10625 24995 10659
rect 27169 10625 27203 10659
rect 8401 10557 8435 10591
rect 10149 10557 10183 10591
rect 13461 10557 13495 10591
rect 18889 10557 18923 10591
rect 19257 10557 19291 10591
rect 23121 10557 23155 10591
rect 5825 10489 5859 10523
rect 12817 10489 12851 10523
rect 18061 10489 18095 10523
rect 3525 10421 3559 10455
rect 4813 10421 4847 10455
rect 7941 10421 7975 10455
rect 10609 10421 10643 10455
rect 11897 10421 11931 10455
rect 15485 10421 15519 10455
rect 22017 10421 22051 10455
rect 26985 10421 27019 10455
rect 4629 10217 4663 10251
rect 8125 10217 8159 10251
rect 11529 10217 11563 10251
rect 14105 10217 14139 10251
rect 16405 10217 16439 10251
rect 17233 10217 17267 10251
rect 18613 10217 18647 10251
rect 19809 10217 19843 10251
rect 20361 10217 20395 10251
rect 21005 10217 21039 10251
rect 25145 10217 25179 10251
rect 3065 10149 3099 10183
rect 6101 10149 6135 10183
rect 12909 10149 12943 10183
rect 23857 10149 23891 10183
rect 4721 10081 4755 10115
rect 10149 10081 10183 10115
rect 12449 10081 12483 10115
rect 15025 10081 15059 10115
rect 25973 10081 26007 10115
rect 1777 10013 1811 10047
rect 2421 10013 2455 10047
rect 3249 10013 3283 10047
rect 4905 10013 4939 10047
rect 5549 10013 5583 10047
rect 5825 10013 5859 10047
rect 5917 10013 5951 10047
rect 6561 10013 6595 10047
rect 6745 10013 6779 10047
rect 7573 10013 7607 10047
rect 7941 10013 7975 10047
rect 9229 10013 9263 10047
rect 9413 10013 9447 10047
rect 9505 10013 9539 10047
rect 10416 10013 10450 10047
rect 12633 10013 12667 10047
rect 14105 10013 14139 10047
rect 14381 10013 14415 10047
rect 15292 10013 15326 10047
rect 16865 10013 16899 10047
rect 17049 10013 17083 10047
rect 17877 10013 17911 10047
rect 18521 10013 18555 10047
rect 19257 10013 19291 10047
rect 19625 10013 19659 10047
rect 20545 10013 20579 10047
rect 21189 10013 21223 10047
rect 21741 10013 21775 10047
rect 21925 10013 21959 10047
rect 23673 10013 23707 10047
rect 24409 10013 24443 10047
rect 25329 10013 25363 10047
rect 3985 9945 4019 9979
rect 4629 9945 4663 9979
rect 5733 9945 5767 9979
rect 7757 9945 7791 9979
rect 7849 9945 7883 9979
rect 13001 9945 13035 9979
rect 19441 9945 19475 9979
rect 19533 9945 19567 9979
rect 22753 9945 22787 9979
rect 26240 9945 26274 9979
rect 1593 9877 1627 9911
rect 2237 9877 2271 9911
rect 4077 9877 4111 9911
rect 5089 9877 5123 9911
rect 6929 9877 6963 9911
rect 9045 9877 9079 9911
rect 14289 9877 14323 9911
rect 17693 9877 17727 9911
rect 22845 9877 22879 9911
rect 24593 9877 24627 9911
rect 27353 9877 27387 9911
rect 23213 9673 23247 9707
rect 2044 9605 2078 9639
rect 10609 9605 10643 9639
rect 10701 9605 10735 9639
rect 12173 9605 12207 9639
rect 15117 9605 15151 9639
rect 18797 9605 18831 9639
rect 18885 9605 18919 9639
rect 25881 9605 25915 9639
rect 4149 9537 4183 9571
rect 7021 9537 7055 9571
rect 8125 9537 8159 9571
rect 8769 9537 8803 9571
rect 9045 9537 9079 9571
rect 9781 9537 9815 9571
rect 10425 9537 10459 9571
rect 10793 9537 10827 9571
rect 11989 9537 12023 9571
rect 13452 9537 13486 9571
rect 15025 9537 15059 9571
rect 15853 9537 15887 9571
rect 16865 9537 16899 9571
rect 18061 9537 18095 9571
rect 18659 9537 18693 9571
rect 18981 9537 19015 9571
rect 19625 9537 19659 9571
rect 19809 9537 19843 9571
rect 20637 9537 20671 9571
rect 21281 9537 21315 9571
rect 22100 9537 22134 9571
rect 23673 9537 23707 9571
rect 23940 9537 23974 9571
rect 25697 9537 25731 9571
rect 25973 9537 26007 9571
rect 27077 9537 27111 9571
rect 1777 9469 1811 9503
rect 3893 9469 3927 9503
rect 6745 9469 6779 9503
rect 8309 9469 8343 9503
rect 13185 9469 13219 9503
rect 19993 9469 20027 9503
rect 21833 9469 21867 9503
rect 10977 9401 11011 9435
rect 15669 9401 15703 9435
rect 3157 9333 3191 9367
rect 5273 9333 5307 9367
rect 8861 9333 8895 9367
rect 9873 9333 9907 9367
rect 14565 9333 14599 9367
rect 16681 9333 16715 9367
rect 17877 9333 17911 9367
rect 19165 9333 19199 9367
rect 20453 9333 20487 9367
rect 21097 9333 21131 9367
rect 25053 9333 25087 9367
rect 25513 9333 25547 9367
rect 27261 9333 27295 9367
rect 12541 9129 12575 9163
rect 13369 9129 13403 9163
rect 18061 9129 18095 9163
rect 18521 9129 18555 9163
rect 19809 9129 19843 9163
rect 26709 9129 26743 9163
rect 1869 9061 1903 9095
rect 3157 9061 3191 9095
rect 6009 9061 6043 9095
rect 21833 9061 21867 9095
rect 23397 9061 23431 9095
rect 4261 8993 4295 9027
rect 6469 8993 6503 9027
rect 6745 8993 6779 9027
rect 9597 8993 9631 9027
rect 10333 8993 10367 9027
rect 13001 8993 13035 9027
rect 14657 8993 14691 9027
rect 24869 8993 24903 9027
rect 1501 8925 1535 8959
rect 1593 8925 1627 8959
rect 1685 8925 1719 8959
rect 2881 8925 2915 8959
rect 2973 8925 3007 8959
rect 3249 8925 3283 8959
rect 3985 8925 4019 8959
rect 10517 8925 10551 8959
rect 10701 8925 10735 8959
rect 11161 8925 11195 8959
rect 13185 8925 13219 8959
rect 16681 8925 16715 8959
rect 16948 8925 16982 8959
rect 18705 8925 18739 8959
rect 19257 8925 19291 8959
rect 19441 8925 19475 8959
rect 19533 8925 19567 8959
rect 19625 8925 19659 8959
rect 20453 8925 20487 8959
rect 20720 8925 20754 8959
rect 22477 8925 22511 8959
rect 23029 8925 23063 8959
rect 23213 8925 23247 8959
rect 23581 8925 23615 8959
rect 23765 8925 23799 8959
rect 25136 8925 25170 8959
rect 26893 8925 26927 8959
rect 27169 8925 27203 8959
rect 5825 8857 5859 8891
rect 8217 8857 8251 8891
rect 9413 8857 9447 8891
rect 11428 8857 11462 8891
rect 14924 8857 14958 8891
rect 2697 8789 2731 8823
rect 8309 8789 8343 8823
rect 16037 8789 16071 8823
rect 22293 8789 22327 8823
rect 26249 8789 26283 8823
rect 27077 8789 27111 8823
rect 2973 8585 3007 8619
rect 8309 8585 8343 8619
rect 12081 8585 12115 8619
rect 13185 8585 13219 8619
rect 13645 8585 13679 8619
rect 17049 8585 17083 8619
rect 18889 8585 18923 8619
rect 19901 8585 19935 8619
rect 23765 8585 23799 8619
rect 2605 8517 2639 8551
rect 2789 8517 2823 8551
rect 4629 8517 4663 8551
rect 8861 8517 8895 8551
rect 9505 8517 9539 8551
rect 11713 8517 11747 8551
rect 12817 8517 12851 8551
rect 12909 8517 12943 8551
rect 15669 8517 15703 8551
rect 17601 8517 17635 8551
rect 17785 8517 17819 8551
rect 22385 8517 22419 8551
rect 23121 8517 23155 8551
rect 2053 8449 2087 8483
rect 3617 8449 3651 8483
rect 5273 8449 5307 8483
rect 5549 8449 5583 8483
rect 7196 8449 7230 8483
rect 8769 8449 8803 8483
rect 11529 8449 11563 8483
rect 11805 8449 11839 8483
rect 11897 8449 11931 8483
rect 12633 8449 12667 8483
rect 13001 8449 13035 8483
rect 13829 8449 13863 8483
rect 14473 8449 14507 8483
rect 15393 8449 15427 8483
rect 15577 8449 15611 8483
rect 15761 8449 15795 8483
rect 16773 8449 16807 8483
rect 16865 8449 16899 8483
rect 18429 8449 18463 8483
rect 19073 8449 19107 8483
rect 19717 8449 19751 8483
rect 20821 8449 20855 8483
rect 23949 8449 23983 8483
rect 24593 8449 24627 8483
rect 25320 8449 25354 8483
rect 26985 8449 27019 8483
rect 5365 8381 5399 8415
rect 6929 8381 6963 8415
rect 9689 8381 9723 8415
rect 10149 8381 10183 8415
rect 10425 8381 10459 8415
rect 14289 8381 14323 8415
rect 19533 8381 19567 8415
rect 25053 8381 25087 8415
rect 3433 8313 3467 8347
rect 5733 8313 5767 8347
rect 14657 8313 14691 8347
rect 15945 8313 15979 8347
rect 18245 8313 18279 8347
rect 20637 8313 20671 8347
rect 22569 8313 22603 8347
rect 27169 8313 27203 8347
rect 1869 8245 1903 8279
rect 4721 8245 4755 8279
rect 5365 8245 5399 8279
rect 23213 8245 23247 8279
rect 24409 8245 24443 8279
rect 26433 8245 26467 8279
rect 5641 8041 5675 8075
rect 9321 8041 9355 8075
rect 13461 8041 13495 8075
rect 15117 8041 15151 8075
rect 18705 8041 18739 8075
rect 26433 8041 26467 8075
rect 6101 7973 6135 8007
rect 12081 7973 12115 8007
rect 14657 7973 14691 8007
rect 19625 7973 19659 8007
rect 5825 7905 5859 7939
rect 7665 7905 7699 7939
rect 10609 7905 10643 7939
rect 17325 7905 17359 7939
rect 1593 7837 1627 7871
rect 3801 7837 3835 7871
rect 5917 7837 5951 7871
rect 6653 7837 6687 7871
rect 6929 7837 6963 7871
rect 7021 7837 7055 7871
rect 7849 7837 7883 7871
rect 10333 7837 10367 7871
rect 11897 7837 11931 7871
rect 13277 7837 13311 7871
rect 14105 7837 14139 7871
rect 14381 7837 14415 7871
rect 14473 7837 14507 7871
rect 15301 7837 15335 7871
rect 15853 7837 15887 7871
rect 16221 7837 16255 7871
rect 17592 7837 17626 7871
rect 20177 7837 20211 7871
rect 20433 7837 20467 7871
rect 22477 7837 22511 7871
rect 24501 7837 24535 7871
rect 24757 7837 24791 7871
rect 26617 7837 26651 7871
rect 26893 7837 26927 7871
rect 1860 7769 1894 7803
rect 4046 7769 4080 7803
rect 5641 7769 5675 7803
rect 6837 7769 6871 7803
rect 8953 7769 8987 7803
rect 9137 7769 9171 7803
rect 12633 7769 12667 7803
rect 12817 7769 12851 7803
rect 14289 7769 14323 7803
rect 16037 7769 16071 7803
rect 16129 7769 16163 7803
rect 19257 7769 19291 7803
rect 19441 7769 19475 7803
rect 22744 7769 22778 7803
rect 2973 7701 3007 7735
rect 5181 7701 5215 7735
rect 7205 7701 7239 7735
rect 8033 7701 8067 7735
rect 16405 7701 16439 7735
rect 21557 7701 21591 7735
rect 23857 7701 23891 7735
rect 25881 7701 25915 7735
rect 26801 7701 26835 7735
rect 2237 7497 2271 7531
rect 10517 7497 10551 7531
rect 17141 7497 17175 7531
rect 18889 7497 18923 7531
rect 23970 7497 24004 7531
rect 24133 7497 24167 7531
rect 24961 7497 24995 7531
rect 26433 7497 26467 7531
rect 27195 7497 27229 7531
rect 1869 7429 1903 7463
rect 2973 7429 3007 7463
rect 5549 7429 5583 7463
rect 7481 7429 7515 7463
rect 8462 7429 8496 7463
rect 10149 7429 10183 7463
rect 11529 7429 11563 7463
rect 12633 7429 12667 7463
rect 17969 7429 18003 7463
rect 22293 7429 22327 7463
rect 23765 7429 23799 7463
rect 24593 7429 24627 7463
rect 26065 7429 26099 7463
rect 26281 7429 26315 7463
rect 26985 7429 27019 7463
rect 24823 7395 24857 7429
rect 2053 7361 2087 7395
rect 3157 7361 3191 7395
rect 3249 7361 3283 7395
rect 3525 7361 3559 7395
rect 4353 7361 4387 7395
rect 5273 7361 5307 7395
rect 5457 7361 5491 7395
rect 5641 7361 5675 7395
rect 6469 7361 6503 7395
rect 6561 7361 6595 7395
rect 7297 7361 7331 7395
rect 10333 7361 10367 7395
rect 11713 7361 11747 7395
rect 11805 7361 11839 7395
rect 12081 7361 12115 7395
rect 13461 7361 13495 7395
rect 14105 7361 14139 7395
rect 14749 7361 14783 7395
rect 15301 7361 15335 7395
rect 16129 7361 16163 7395
rect 16773 7361 16807 7395
rect 16957 7361 16991 7395
rect 17601 7361 17635 7395
rect 17785 7361 17819 7395
rect 19073 7361 19107 7395
rect 19165 7361 19199 7395
rect 19441 7361 19475 7395
rect 19901 7361 19935 7395
rect 20085 7361 20119 7395
rect 20913 7361 20947 7395
rect 23121 7361 23155 7395
rect 25605 7361 25639 7395
rect 8217 7293 8251 7327
rect 11989 7293 12023 7327
rect 15485 7293 15519 7327
rect 5825 7225 5859 7259
rect 13277 7225 13311 7259
rect 20269 7225 20303 7259
rect 27353 7225 27387 7259
rect 3433 7157 3467 7191
rect 4445 7157 4479 7191
rect 6745 7157 6779 7191
rect 9597 7157 9631 7191
rect 12725 7157 12759 7191
rect 13921 7157 13955 7191
rect 14565 7157 14599 7191
rect 15945 7157 15979 7191
rect 19349 7157 19383 7191
rect 20729 7157 20763 7191
rect 22385 7157 22419 7191
rect 22937 7157 22971 7191
rect 23949 7157 23983 7191
rect 24777 7157 24811 7191
rect 25421 7157 25455 7191
rect 26249 7157 26283 7191
rect 27169 7157 27203 7191
rect 6745 6953 6779 6987
rect 12725 6953 12759 6987
rect 24593 6953 24627 6987
rect 27353 6953 27387 6987
rect 19717 6885 19751 6919
rect 24777 6885 24811 6919
rect 3801 6817 3835 6851
rect 8953 6817 8987 6851
rect 10425 6817 10459 6851
rect 19257 6817 19291 6851
rect 25973 6817 26007 6851
rect 3249 6749 3283 6783
rect 4077 6749 4111 6783
rect 5273 6749 5307 6783
rect 6101 6749 6135 6783
rect 7573 6749 7607 6783
rect 7849 6749 7883 6783
rect 9229 6749 9263 6783
rect 10692 6749 10726 6783
rect 12449 6749 12483 6783
rect 12601 6749 12635 6783
rect 12817 6749 12851 6783
rect 13461 6749 13495 6783
rect 14565 6749 14599 6783
rect 15025 6749 15059 6783
rect 17233 6749 17267 6783
rect 17500 6749 17534 6783
rect 19441 6749 19475 6783
rect 19533 6749 19567 6783
rect 19809 6749 19843 6783
rect 20545 6749 20579 6783
rect 22845 6749 22879 6783
rect 23581 6749 23615 6783
rect 25237 6749 25271 6783
rect 1961 6681 1995 6715
rect 2145 6681 2179 6715
rect 5089 6681 5123 6715
rect 5457 6681 5491 6715
rect 6653 6681 6687 6715
rect 15292 6681 15326 6715
rect 20790 6681 20824 6715
rect 24409 6681 24443 6715
rect 26218 6681 26252 6715
rect 2329 6613 2363 6647
rect 3065 6613 3099 6647
rect 5917 6613 5951 6647
rect 11805 6613 11839 6647
rect 12265 6613 12299 6647
rect 13277 6613 13311 6647
rect 14381 6613 14415 6647
rect 16405 6613 16439 6647
rect 18613 6613 18647 6647
rect 21925 6613 21959 6647
rect 23029 6613 23063 6647
rect 23765 6613 23799 6647
rect 24619 6613 24653 6647
rect 25421 6613 25455 6647
rect 3341 6409 3375 6443
rect 5457 6409 5491 6443
rect 9137 6409 9171 6443
rect 10517 6409 10551 6443
rect 16037 6409 16071 6443
rect 16957 6409 16991 6443
rect 24317 6409 24351 6443
rect 27185 6409 27219 6443
rect 27353 6409 27387 6443
rect 1768 6341 1802 6375
rect 8493 6341 8527 6375
rect 13084 6341 13118 6375
rect 14657 6341 14691 6375
rect 15669 6341 15703 6375
rect 20168 6341 20202 6375
rect 23949 6341 23983 6375
rect 24165 6341 24199 6375
rect 25044 6341 25078 6375
rect 26985 6341 27019 6375
rect 3525 6273 3559 6307
rect 4344 6273 4378 6307
rect 6377 6273 6411 6307
rect 6633 6273 6667 6307
rect 9321 6273 9355 6307
rect 9413 6273 9447 6307
rect 9689 6273 9723 6307
rect 10149 6273 10183 6307
rect 10333 6273 10367 6307
rect 12817 6273 12851 6307
rect 14841 6273 14875 6307
rect 14933 6273 14967 6307
rect 15191 6273 15225 6307
rect 15853 6273 15887 6307
rect 17141 6273 17175 6307
rect 17233 6273 17267 6307
rect 17509 6273 17543 6307
rect 18153 6273 18187 6307
rect 18797 6273 18831 6307
rect 19441 6273 19475 6307
rect 19901 6273 19935 6307
rect 22109 6273 22143 6307
rect 22376 6273 22410 6307
rect 24777 6273 24811 6307
rect 1501 6205 1535 6239
rect 4077 6205 4111 6239
rect 11529 6205 11563 6239
rect 11805 6205 11839 6239
rect 19257 6137 19291 6171
rect 2881 6069 2915 6103
rect 7757 6069 7791 6103
rect 8585 6069 8619 6103
rect 9597 6069 9631 6103
rect 14197 6069 14231 6103
rect 15117 6069 15151 6103
rect 17417 6069 17451 6103
rect 17969 6069 18003 6103
rect 18613 6069 18647 6103
rect 21281 6069 21315 6103
rect 23489 6069 23523 6103
rect 24133 6069 24167 6103
rect 26157 6069 26191 6103
rect 27169 6069 27203 6103
rect 2697 5865 2731 5899
rect 3157 5865 3191 5899
rect 5089 5865 5123 5899
rect 13461 5865 13495 5899
rect 20821 5865 20855 5899
rect 21005 5865 21039 5899
rect 22293 5865 22327 5899
rect 22477 5865 22511 5899
rect 24593 5865 24627 5899
rect 1409 5797 1443 5831
rect 5549 5797 5583 5831
rect 14749 5797 14783 5831
rect 15669 5797 15703 5831
rect 16681 5797 16715 5831
rect 21465 5797 21499 5831
rect 25421 5797 25455 5831
rect 3801 5729 3835 5763
rect 9413 5729 9447 5763
rect 10517 5729 10551 5763
rect 17325 5729 17359 5763
rect 25973 5729 26007 5763
rect 1593 5661 1627 5695
rect 2237 5661 2271 5695
rect 2881 5661 2915 5695
rect 2973 5661 3007 5695
rect 3249 5661 3283 5695
rect 4077 5661 4111 5695
rect 5273 5661 5307 5695
rect 5365 5661 5399 5695
rect 5641 5661 5675 5695
rect 7849 5661 7883 5695
rect 8953 5661 8987 5695
rect 9137 5661 9171 5695
rect 9229 5661 9263 5695
rect 9505 5661 9539 5695
rect 10784 5661 10818 5695
rect 12541 5661 12575 5695
rect 13168 5661 13202 5695
rect 13277 5661 13311 5695
rect 13553 5661 13587 5695
rect 14381 5661 14415 5695
rect 15209 5661 15243 5695
rect 15393 5661 15427 5695
rect 15485 5661 15519 5695
rect 15761 5661 15795 5695
rect 16405 5661 16439 5695
rect 16497 5661 16531 5695
rect 16773 5661 16807 5695
rect 17581 5661 17615 5695
rect 19441 5661 19475 5695
rect 20085 5661 20119 5695
rect 21649 5661 21683 5695
rect 23121 5661 23155 5695
rect 23581 5661 23615 5695
rect 25237 5661 25271 5695
rect 26240 5661 26274 5695
rect 6653 5593 6687 5627
rect 6837 5593 6871 5627
rect 8033 5593 8067 5627
rect 14565 5593 14599 5627
rect 20637 5593 20671 5627
rect 22109 5593 22143 5627
rect 24409 5593 24443 5627
rect 2053 5525 2087 5559
rect 7021 5525 7055 5559
rect 8217 5525 8251 5559
rect 11897 5525 11931 5559
rect 12357 5525 12391 5559
rect 13001 5525 13035 5559
rect 16221 5525 16255 5559
rect 18705 5525 18739 5559
rect 19257 5525 19291 5559
rect 19901 5525 19935 5559
rect 20837 5525 20871 5559
rect 22309 5525 22343 5559
rect 22937 5525 22971 5559
rect 23765 5525 23799 5559
rect 24609 5525 24643 5559
rect 24777 5525 24811 5559
rect 27353 5525 27387 5559
rect 3065 5321 3099 5355
rect 6653 5321 6687 5355
rect 9229 5321 9263 5355
rect 9965 5321 9999 5355
rect 15669 5321 15703 5355
rect 20637 5321 20671 5355
rect 23949 5321 23983 5355
rect 24777 5321 24811 5355
rect 2697 5253 2731 5287
rect 3801 5253 3835 5287
rect 4997 5253 5031 5287
rect 11529 5253 11563 5287
rect 12449 5253 12483 5287
rect 13461 5253 13495 5287
rect 14534 5253 14568 5287
rect 20269 5253 20303 5287
rect 22201 5253 22235 5287
rect 23581 5253 23615 5287
rect 23797 5253 23831 5287
rect 24409 5253 24443 5287
rect 24609 5253 24643 5287
rect 26985 5253 27019 5287
rect 27185 5253 27219 5287
rect 20499 5219 20533 5253
rect 1869 5185 1903 5219
rect 2053 5185 2087 5219
rect 2881 5185 2915 5219
rect 3985 5185 4019 5219
rect 4077 5185 4111 5219
rect 4353 5185 4387 5219
rect 5181 5185 5215 5219
rect 6837 5185 6871 5219
rect 6929 5185 6963 5219
rect 7205 5185 7239 5219
rect 8105 5185 8139 5219
rect 10149 5185 10183 5219
rect 10241 5185 10275 5219
rect 10517 5185 10551 5219
rect 11805 5185 11839 5219
rect 12633 5185 12667 5219
rect 12817 5185 12851 5219
rect 13645 5185 13679 5219
rect 14289 5185 14323 5219
rect 16681 5185 16715 5219
rect 16937 5185 16971 5219
rect 18797 5185 18831 5219
rect 19533 5185 19567 5219
rect 21281 5185 21315 5219
rect 22063 5185 22097 5219
rect 22293 5185 22327 5219
rect 22845 5185 22879 5219
rect 7849 5117 7883 5151
rect 11621 5117 11655 5151
rect 25605 5117 25639 5151
rect 25881 5117 25915 5151
rect 4261 5049 4295 5083
rect 13829 5049 13863 5083
rect 27353 5049 27387 5083
rect 2237 4981 2271 5015
rect 5365 4981 5399 5015
rect 7113 4981 7147 5015
rect 10425 4981 10459 5015
rect 11805 4981 11839 5015
rect 11989 4981 12023 5015
rect 18061 4981 18095 5015
rect 18613 4981 18647 5015
rect 19717 4981 19751 5015
rect 20453 4981 20487 5015
rect 21097 4981 21131 5015
rect 21833 4981 21867 5015
rect 23029 4981 23063 5015
rect 23765 4981 23799 5015
rect 24584 4981 24618 5015
rect 27169 4981 27203 5015
rect 3801 4777 3835 4811
rect 7757 4777 7791 4811
rect 8217 4777 8251 4811
rect 9597 4777 9631 4811
rect 13553 4777 13587 4811
rect 17141 4777 17175 4811
rect 26893 4777 26927 4811
rect 6929 4709 6963 4743
rect 10471 4709 10505 4743
rect 27077 4709 27111 4743
rect 4261 4641 4295 4675
rect 7849 4641 7883 4675
rect 19257 4641 19291 4675
rect 1409 4573 1443 4607
rect 3985 4573 4019 4607
rect 4077 4573 4111 4607
rect 4353 4573 4387 4607
rect 5089 4573 5123 4607
rect 7113 4573 7147 4607
rect 7757 4573 7791 4607
rect 8033 4573 8067 4607
rect 9321 4573 9355 4607
rect 9505 4573 9539 4607
rect 9597 4573 9631 4607
rect 10241 4573 10275 4607
rect 11713 4573 11747 4607
rect 12173 4573 12207 4607
rect 14289 4573 14323 4607
rect 14749 4573 14783 4607
rect 15485 4573 15519 4607
rect 16773 4573 16807 4607
rect 17601 4573 17635 4607
rect 18337 4573 18371 4607
rect 21097 4573 21131 4607
rect 23121 4573 23155 4607
rect 23397 4573 23431 4607
rect 24593 4573 24627 4607
rect 1676 4505 1710 4539
rect 5356 4505 5390 4539
rect 12418 4505 12452 4539
rect 16957 4505 16991 4539
rect 19524 4505 19558 4539
rect 21364 4505 21398 4539
rect 24860 4505 24894 4539
rect 26709 4505 26743 4539
rect 26925 4505 26959 4539
rect 2789 4437 2823 4471
rect 6469 4437 6503 4471
rect 9781 4437 9815 4471
rect 11529 4437 11563 4471
rect 14105 4437 14139 4471
rect 14933 4437 14967 4471
rect 15669 4437 15703 4471
rect 17785 4437 17819 4471
rect 18521 4437 18555 4471
rect 20637 4437 20671 4471
rect 22477 4437 22511 4471
rect 22937 4437 22971 4471
rect 23305 4437 23339 4471
rect 25973 4437 26007 4471
rect 1685 4233 1719 4267
rect 4905 4233 4939 4267
rect 5365 4233 5399 4267
rect 7849 4233 7883 4267
rect 23857 4233 23891 4267
rect 24777 4233 24811 4267
rect 26341 4233 26375 4267
rect 27185 4233 27219 4267
rect 4445 4165 4479 4199
rect 12909 4165 12943 4199
rect 15761 4165 15795 4199
rect 18705 4165 18739 4199
rect 22744 4165 22778 4199
rect 26249 4165 26283 4199
rect 26985 4165 27019 4199
rect 1869 4097 1903 4131
rect 2605 4097 2639 4131
rect 2872 4097 2906 4131
rect 4721 4097 4755 4131
rect 5549 4097 5583 4131
rect 6469 4097 6503 4131
rect 6653 4097 6687 4131
rect 6745 4097 6779 4131
rect 7021 4097 7055 4131
rect 7573 4097 7607 4131
rect 7665 4097 7699 4131
rect 8309 4097 8343 4131
rect 8565 4097 8599 4131
rect 11529 4097 11563 4131
rect 11713 4097 11747 4131
rect 11801 4097 11835 4131
rect 11943 4097 11977 4131
rect 12725 4097 12759 4131
rect 13369 4097 13403 4131
rect 14105 4097 14139 4131
rect 14841 4097 14875 4131
rect 16681 4097 16715 4131
rect 17785 4097 17819 4131
rect 19625 4097 19659 4131
rect 20545 4097 20579 4131
rect 21005 4097 21039 4131
rect 22017 4097 22051 4131
rect 24593 4097 24627 4131
rect 24869 4097 24903 4131
rect 25329 4097 25363 4131
rect 4629 4029 4663 4063
rect 6929 4029 6963 4063
rect 10149 4029 10183 4063
rect 10425 4029 10459 4063
rect 12541 4029 12575 4063
rect 18245 4029 18279 4063
rect 19165 4029 19199 4063
rect 22477 4029 22511 4063
rect 9689 3961 9723 3995
rect 12081 3961 12115 3995
rect 15025 3961 15059 3995
rect 16865 3961 16899 3995
rect 18153 3961 18187 3995
rect 18981 3961 19015 3995
rect 20361 3961 20395 3995
rect 21189 3961 21223 3995
rect 24409 3961 24443 3995
rect 25513 3961 25547 3995
rect 27353 3961 27387 3995
rect 3985 3893 4019 3927
rect 4445 3893 4479 3927
rect 13553 3893 13587 3927
rect 14289 3893 14323 3927
rect 15853 3893 15887 3927
rect 19809 3893 19843 3927
rect 21833 3893 21867 3927
rect 27169 3893 27203 3927
rect 2421 3689 2455 3723
rect 7297 3689 7331 3723
rect 7481 3689 7515 3723
rect 10149 3689 10183 3723
rect 15485 3689 15519 3723
rect 16497 3689 16531 3723
rect 17325 3689 17359 3723
rect 18613 3689 18647 3723
rect 21097 3689 21131 3723
rect 21281 3689 21315 3723
rect 26157 3689 26191 3723
rect 26985 3689 27019 3723
rect 3065 3621 3099 3655
rect 11989 3621 12023 3655
rect 12817 3621 12851 3655
rect 20453 3621 20487 3655
rect 25329 3621 25363 3655
rect 26341 3621 26375 3655
rect 27169 3621 27203 3655
rect 5549 3553 5583 3587
rect 7941 3553 7975 3587
rect 16129 3553 16163 3587
rect 16957 3553 16991 3587
rect 18245 3553 18279 3587
rect 19625 3553 19659 3587
rect 20085 3553 20119 3587
rect 1961 3485 1995 3519
rect 2605 3485 2639 3519
rect 3249 3485 3283 3519
rect 4261 3485 4295 3519
rect 4721 3485 4755 3519
rect 4905 3487 4939 3521
rect 5733 3485 5767 3519
rect 6561 3485 6595 3519
rect 7205 3485 7239 3519
rect 7297 3485 7331 3519
rect 8125 3485 8159 3519
rect 9137 3485 9171 3519
rect 9597 3485 9631 3519
rect 9873 3485 9907 3519
rect 9965 3485 9999 3519
rect 10977 3485 11011 3519
rect 11437 3485 11471 3519
rect 11713 3485 11747 3519
rect 11805 3485 11839 3519
rect 12449 3485 12483 3519
rect 12633 3485 12667 3519
rect 13277 3485 13311 3519
rect 14105 3485 14139 3519
rect 14372 3485 14406 3519
rect 16313 3485 16347 3519
rect 17141 3485 17175 3519
rect 18429 3485 18463 3519
rect 19257 3485 19291 3519
rect 19441 3485 19475 3519
rect 20269 3485 20303 3519
rect 21741 3485 21775 3519
rect 22017 3485 22051 3519
rect 23213 3485 23247 3519
rect 23489 3485 23523 3519
rect 24593 3485 24627 3519
rect 24869 3485 24903 3519
rect 25513 3485 25547 3519
rect 5089 3417 5123 3451
rect 7021 3417 7055 3451
rect 9781 3417 9815 3451
rect 11621 3417 11655 3451
rect 20913 3417 20947 3451
rect 25973 3417 26007 3451
rect 26801 3417 26835 3451
rect 1777 3349 1811 3383
rect 4077 3349 4111 3383
rect 5917 3349 5951 3383
rect 6377 3349 6411 3383
rect 8309 3349 8343 3383
rect 8953 3349 8987 3383
rect 10793 3349 10827 3383
rect 13461 3349 13495 3383
rect 21113 3349 21147 3383
rect 23029 3349 23063 3383
rect 23397 3349 23431 3383
rect 24409 3349 24443 3383
rect 24777 3349 24811 3383
rect 26173 3349 26207 3383
rect 27001 3349 27035 3383
rect 9597 3145 9631 3179
rect 10609 3145 10643 3179
rect 14197 3145 14231 3179
rect 15209 3145 15243 3179
rect 18705 3145 18739 3179
rect 25513 3145 25547 3179
rect 26183 3145 26217 3179
rect 27185 3145 27219 3179
rect 5365 3077 5399 3111
rect 5457 3077 5491 3111
rect 8484 3077 8518 3111
rect 10241 3077 10275 3111
rect 20637 3077 20671 3111
rect 20853 3077 20887 3111
rect 24400 3077 24434 3111
rect 25973 3077 26007 3111
rect 26985 3077 27019 3111
rect 1501 3009 1535 3043
rect 1768 3009 1802 3043
rect 3341 3009 3375 3043
rect 3608 3009 3642 3043
rect 5181 3009 5215 3043
rect 5549 3009 5583 3043
rect 6377 3009 6411 3043
rect 6633 3009 6667 3043
rect 8217 3009 8251 3043
rect 10057 3009 10091 3043
rect 10333 3009 10367 3043
rect 10425 3009 10459 3043
rect 11529 3009 11563 3043
rect 11796 3009 11830 3043
rect 13553 3009 13587 3043
rect 13737 3009 13771 3043
rect 14381 3009 14415 3043
rect 15025 3009 15059 3043
rect 15853 3009 15887 3043
rect 16773 3009 16807 3043
rect 16865 3009 16899 3043
rect 17693 3009 17727 3043
rect 18541 3009 18575 3043
rect 19717 3009 19751 3043
rect 22109 3009 22143 3043
rect 22376 3009 22410 3043
rect 24133 3009 24167 3043
rect 13369 2941 13403 2975
rect 14841 2941 14875 2975
rect 15669 2941 15703 2975
rect 17509 2941 17543 2975
rect 18337 2941 18371 2975
rect 20177 2941 20211 2975
rect 5733 2873 5767 2907
rect 17049 2873 17083 2907
rect 20085 2873 20119 2907
rect 26341 2873 26375 2907
rect 27353 2873 27387 2907
rect 2881 2805 2915 2839
rect 4721 2805 4755 2839
rect 7757 2805 7791 2839
rect 12909 2805 12943 2839
rect 16037 2805 16071 2839
rect 17877 2805 17911 2839
rect 20821 2805 20855 2839
rect 21005 2805 21039 2839
rect 23489 2805 23523 2839
rect 26157 2805 26191 2839
rect 27169 2805 27203 2839
rect 3801 2601 3835 2635
rect 5273 2601 5307 2635
rect 8125 2601 8159 2635
rect 8953 2601 8987 2635
rect 14749 2601 14783 2635
rect 15393 2601 15427 2635
rect 15945 2601 15979 2635
rect 21097 2601 21131 2635
rect 22017 2601 22051 2635
rect 22201 2601 22235 2635
rect 23581 2601 23615 2635
rect 7297 2533 7331 2567
rect 10701 2533 10735 2567
rect 13185 2533 13219 2567
rect 20177 2533 20211 2567
rect 22845 2533 22879 2567
rect 25329 2533 25363 2567
rect 11529 2465 11563 2499
rect 12817 2465 12851 2499
rect 2697 2397 2731 2431
rect 3985 2397 4019 2431
rect 4721 2397 4755 2431
rect 4997 2397 5031 2431
rect 5089 2397 5123 2431
rect 6745 2397 6779 2431
rect 7113 2397 7147 2431
rect 7849 2397 7883 2431
rect 7941 2397 7975 2431
rect 9137 2397 9171 2431
rect 10149 2397 10183 2431
rect 10333 2397 10367 2431
rect 10517 2397 10551 2431
rect 11713 2397 11747 2431
rect 13001 2397 13035 2431
rect 14381 2397 14415 2431
rect 14565 2397 14599 2431
rect 15209 2397 15243 2431
rect 16129 2397 16163 2431
rect 16681 2397 16715 2431
rect 17417 2397 17451 2431
rect 18153 2397 18187 2431
rect 19257 2397 19291 2431
rect 19993 2397 20027 2431
rect 22661 2397 22695 2431
rect 23397 2397 23431 2431
rect 24409 2397 24443 2431
rect 25145 2397 25179 2431
rect 25881 2397 25915 2431
rect 1869 2329 1903 2363
rect 4905 2329 4939 2363
rect 6929 2329 6963 2363
rect 7021 2329 7055 2363
rect 10425 2329 10459 2363
rect 20913 2329 20947 2363
rect 21113 2329 21147 2363
rect 21833 2329 21867 2363
rect 27169 2329 27203 2363
rect 2145 2261 2179 2295
rect 2881 2261 2915 2295
rect 11897 2261 11931 2295
rect 16865 2261 16899 2295
rect 17601 2261 17635 2295
rect 18337 2261 18371 2295
rect 19441 2261 19475 2295
rect 21281 2261 21315 2295
rect 22033 2261 22067 2295
rect 24593 2261 24627 2295
rect 26065 2261 26099 2295
rect 27261 2261 27295 2295
<< metal1 >>
rect 1104 28858 28060 28880
rect 1104 28806 5442 28858
rect 5494 28806 5506 28858
rect 5558 28806 5570 28858
rect 5622 28806 5634 28858
rect 5686 28806 5698 28858
rect 5750 28806 14428 28858
rect 14480 28806 14492 28858
rect 14544 28806 14556 28858
rect 14608 28806 14620 28858
rect 14672 28806 14684 28858
rect 14736 28806 23413 28858
rect 23465 28806 23477 28858
rect 23529 28806 23541 28858
rect 23593 28806 23605 28858
rect 23657 28806 23669 28858
rect 23721 28806 28060 28858
rect 1104 28784 28060 28806
rect 10137 28747 10195 28753
rect 10137 28713 10149 28747
rect 10183 28744 10195 28747
rect 12802 28744 12808 28756
rect 10183 28716 12808 28744
rect 10183 28713 10195 28716
rect 10137 28707 10195 28713
rect 12802 28704 12808 28716
rect 12860 28704 12866 28756
rect 15746 28744 15752 28756
rect 12912 28716 15752 28744
rect 8113 28679 8171 28685
rect 8113 28645 8125 28679
rect 8159 28676 8171 28679
rect 9122 28676 9128 28688
rect 8159 28648 9128 28676
rect 8159 28645 8171 28648
rect 8113 28639 8171 28645
rect 9122 28636 9128 28648
rect 9180 28636 9186 28688
rect 12912 28608 12940 28716
rect 15746 28704 15752 28716
rect 15804 28704 15810 28756
rect 16666 28704 16672 28756
rect 16724 28744 16730 28756
rect 23109 28747 23167 28753
rect 23109 28744 23121 28747
rect 16724 28716 23121 28744
rect 16724 28704 16730 28716
rect 23109 28713 23121 28716
rect 23155 28713 23167 28747
rect 23109 28707 23167 28713
rect 13538 28636 13544 28688
rect 13596 28676 13602 28688
rect 13725 28679 13783 28685
rect 13725 28676 13737 28679
rect 13596 28648 13737 28676
rect 13596 28636 13602 28648
rect 13725 28645 13737 28648
rect 13771 28645 13783 28679
rect 13725 28639 13783 28645
rect 18322 28636 18328 28688
rect 18380 28676 18386 28688
rect 20073 28679 20131 28685
rect 20073 28676 20085 28679
rect 18380 28648 20085 28676
rect 18380 28636 18386 28648
rect 20073 28645 20085 28648
rect 20119 28645 20131 28679
rect 20073 28639 20131 28645
rect 20162 28636 20168 28688
rect 20220 28676 20226 28688
rect 21453 28679 21511 28685
rect 20220 28648 20392 28676
rect 20220 28636 20226 28648
rect 13556 28608 13584 28636
rect 10336 28580 12940 28608
rect 13004 28580 13584 28608
rect 13909 28611 13967 28617
rect 8113 28543 8171 28549
rect 8113 28509 8125 28543
rect 8159 28540 8171 28543
rect 8294 28540 8300 28552
rect 8159 28512 8300 28540
rect 8159 28509 8171 28512
rect 8113 28503 8171 28509
rect 8294 28500 8300 28512
rect 8352 28500 8358 28552
rect 8386 28500 8392 28552
rect 8444 28540 8450 28552
rect 10336 28549 10364 28580
rect 9493 28543 9551 28549
rect 8444 28512 8489 28540
rect 8444 28500 8450 28512
rect 9493 28509 9505 28543
rect 9539 28540 9551 28543
rect 10321 28543 10379 28549
rect 10321 28540 10333 28543
rect 9539 28512 10333 28540
rect 9539 28509 9551 28512
rect 9493 28503 9551 28509
rect 10321 28509 10333 28512
rect 10367 28509 10379 28543
rect 10321 28503 10379 28509
rect 10502 28500 10508 28552
rect 10560 28540 10566 28552
rect 10965 28543 11023 28549
rect 10965 28540 10977 28543
rect 10560 28512 10977 28540
rect 10560 28500 10566 28512
rect 10965 28509 10977 28512
rect 11011 28509 11023 28543
rect 11330 28540 11336 28552
rect 11291 28512 11336 28540
rect 10965 28503 11023 28509
rect 11330 28500 11336 28512
rect 11388 28500 11394 28552
rect 13004 28549 13032 28580
rect 13909 28577 13921 28611
rect 13955 28608 13967 28611
rect 13998 28608 14004 28620
rect 13955 28580 14004 28608
rect 13955 28577 13967 28580
rect 13909 28571 13967 28577
rect 13998 28568 14004 28580
rect 14056 28568 14062 28620
rect 19242 28568 19248 28620
rect 19300 28608 19306 28620
rect 19705 28611 19763 28617
rect 19705 28608 19717 28611
rect 19300 28580 19717 28608
rect 19300 28568 19306 28580
rect 19705 28577 19717 28580
rect 19751 28608 19763 28611
rect 20364 28608 20392 28648
rect 21453 28645 21465 28679
rect 21499 28676 21511 28679
rect 22094 28676 22100 28688
rect 21499 28648 22100 28676
rect 21499 28645 21511 28648
rect 21453 28639 21511 28645
rect 22094 28636 22100 28648
rect 22152 28636 22158 28688
rect 19751 28580 20300 28608
rect 20364 28580 22094 28608
rect 19751 28577 19763 28580
rect 19705 28571 19763 28577
rect 12345 28543 12403 28549
rect 12345 28540 12357 28543
rect 11992 28512 12357 28540
rect 8570 28472 8576 28484
rect 8531 28444 8576 28472
rect 8570 28432 8576 28444
rect 8628 28432 8634 28484
rect 8754 28472 8760 28484
rect 8715 28444 8760 28472
rect 8754 28432 8760 28444
rect 8812 28432 8818 28484
rect 9861 28475 9919 28481
rect 9861 28441 9873 28475
rect 9907 28472 9919 28475
rect 10520 28472 10548 28500
rect 9907 28444 10548 28472
rect 9907 28441 9919 28444
rect 9861 28435 9919 28441
rect 11992 28416 12020 28512
rect 12345 28509 12357 28512
rect 12391 28509 12403 28543
rect 12345 28503 12403 28509
rect 12989 28543 13047 28549
rect 12989 28509 13001 28543
rect 13035 28509 13047 28543
rect 13170 28540 13176 28552
rect 13131 28512 13176 28540
rect 12989 28503 13047 28509
rect 13170 28500 13176 28512
rect 13228 28500 13234 28552
rect 13633 28543 13691 28549
rect 13633 28509 13645 28543
rect 13679 28540 13691 28543
rect 13722 28540 13728 28552
rect 13679 28512 13728 28540
rect 13679 28509 13691 28512
rect 13633 28503 13691 28509
rect 13722 28500 13728 28512
rect 13780 28500 13786 28552
rect 14553 28543 14611 28549
rect 14553 28509 14565 28543
rect 14599 28540 14611 28543
rect 15010 28540 15016 28552
rect 14599 28512 15016 28540
rect 14599 28509 14611 28512
rect 14553 28503 14611 28509
rect 15010 28500 15016 28512
rect 15068 28500 15074 28552
rect 16025 28543 16083 28549
rect 16025 28540 16037 28543
rect 15580 28512 16037 28540
rect 15580 28416 15608 28512
rect 16025 28509 16037 28512
rect 16071 28509 16083 28543
rect 16482 28540 16488 28552
rect 16443 28512 16488 28540
rect 16025 28503 16083 28509
rect 16482 28500 16488 28512
rect 16540 28500 16546 28552
rect 17037 28543 17095 28549
rect 17037 28509 17049 28543
rect 17083 28540 17095 28543
rect 17497 28543 17555 28549
rect 17497 28540 17509 28543
rect 17083 28512 17509 28540
rect 17083 28509 17095 28512
rect 17037 28503 17095 28509
rect 17497 28509 17509 28512
rect 17543 28540 17555 28543
rect 17586 28540 17592 28552
rect 17543 28512 17592 28540
rect 17543 28509 17555 28512
rect 17497 28503 17555 28509
rect 17586 28500 17592 28512
rect 17644 28500 17650 28552
rect 18138 28540 18144 28552
rect 18099 28512 18144 28540
rect 18138 28500 18144 28512
rect 18196 28500 18202 28552
rect 18690 28540 18696 28552
rect 18651 28512 18696 28540
rect 18690 28500 18696 28512
rect 18748 28500 18754 28552
rect 18877 28543 18935 28549
rect 18877 28509 18889 28543
rect 18923 28540 18935 28543
rect 19794 28540 19800 28552
rect 18923 28512 19800 28540
rect 18923 28509 18935 28512
rect 18877 28503 18935 28509
rect 19794 28500 19800 28512
rect 19852 28500 19858 28552
rect 20272 28549 20300 28580
rect 20257 28543 20315 28549
rect 20257 28509 20269 28543
rect 20303 28509 20315 28543
rect 20257 28503 20315 28509
rect 20622 28500 20628 28552
rect 20680 28540 20686 28552
rect 20901 28543 20959 28549
rect 20901 28540 20913 28543
rect 20680 28512 20913 28540
rect 20680 28500 20686 28512
rect 20901 28509 20913 28512
rect 20947 28540 20959 28543
rect 21177 28543 21235 28549
rect 21177 28540 21189 28543
rect 20947 28512 21189 28540
rect 20947 28509 20959 28512
rect 20901 28503 20959 28509
rect 21177 28509 21189 28512
rect 21223 28509 21235 28543
rect 21634 28540 21640 28552
rect 21595 28512 21640 28540
rect 21177 28503 21235 28509
rect 21634 28500 21640 28512
rect 21692 28500 21698 28552
rect 22066 28540 22094 28580
rect 22189 28543 22247 28549
rect 22189 28540 22201 28543
rect 22066 28512 22201 28540
rect 22189 28509 22201 28512
rect 22235 28540 22247 28543
rect 22649 28543 22707 28549
rect 22649 28540 22661 28543
rect 22235 28512 22661 28540
rect 22235 28509 22247 28512
rect 22189 28503 22247 28509
rect 22649 28509 22661 28512
rect 22695 28509 22707 28543
rect 22649 28503 22707 28509
rect 22922 28500 22928 28552
rect 22980 28540 22986 28552
rect 23293 28543 23351 28549
rect 23293 28540 23305 28543
rect 22980 28512 23305 28540
rect 22980 28500 22986 28512
rect 23293 28509 23305 28512
rect 23339 28540 23351 28543
rect 23569 28543 23627 28549
rect 23569 28540 23581 28543
rect 23339 28512 23581 28540
rect 23339 28509 23351 28512
rect 23293 28503 23351 28509
rect 23569 28509 23581 28512
rect 23615 28509 23627 28543
rect 27338 28540 27344 28552
rect 27299 28512 27344 28540
rect 23569 28503 23627 28509
rect 27338 28500 27344 28512
rect 27396 28500 27402 28552
rect 21818 28472 21824 28484
rect 15856 28444 21824 28472
rect 4338 28364 4344 28416
rect 4396 28404 4402 28416
rect 7098 28404 7104 28416
rect 4396 28376 7104 28404
rect 4396 28364 4402 28376
rect 7098 28364 7104 28376
rect 7156 28364 7162 28416
rect 7466 28364 7472 28416
rect 7524 28404 7530 28416
rect 8297 28407 8355 28413
rect 8297 28404 8309 28407
rect 7524 28376 8309 28404
rect 7524 28364 7530 28376
rect 8297 28373 8309 28376
rect 8343 28404 8355 28407
rect 10410 28404 10416 28416
rect 8343 28376 10416 28404
rect 8343 28373 8355 28376
rect 8297 28367 8355 28373
rect 10410 28364 10416 28376
rect 10468 28364 10474 28416
rect 10781 28407 10839 28413
rect 10781 28373 10793 28407
rect 10827 28404 10839 28407
rect 10962 28404 10968 28416
rect 10827 28376 10968 28404
rect 10827 28373 10839 28376
rect 10781 28367 10839 28373
rect 10962 28364 10968 28376
rect 11020 28364 11026 28416
rect 11146 28404 11152 28416
rect 11107 28376 11152 28404
rect 11146 28364 11152 28376
rect 11204 28364 11210 28416
rect 11885 28407 11943 28413
rect 11885 28373 11897 28407
rect 11931 28404 11943 28407
rect 11974 28404 11980 28416
rect 11931 28376 11980 28404
rect 11931 28373 11943 28376
rect 11885 28367 11943 28373
rect 11974 28364 11980 28376
rect 12032 28364 12038 28416
rect 12158 28404 12164 28416
rect 12119 28376 12164 28404
rect 12158 28364 12164 28376
rect 12216 28364 12222 28416
rect 13078 28404 13084 28416
rect 13039 28376 13084 28404
rect 13078 28364 13084 28376
rect 13136 28364 13142 28416
rect 13814 28364 13820 28416
rect 13872 28404 13878 28416
rect 13909 28407 13967 28413
rect 13909 28404 13921 28407
rect 13872 28376 13921 28404
rect 13872 28364 13878 28376
rect 13909 28373 13921 28376
rect 13955 28373 13967 28407
rect 14826 28404 14832 28416
rect 14787 28376 14832 28404
rect 13909 28367 13967 28373
rect 14826 28364 14832 28376
rect 14884 28364 14890 28416
rect 15562 28404 15568 28416
rect 15523 28376 15568 28404
rect 15562 28364 15568 28376
rect 15620 28364 15626 28416
rect 15856 28413 15884 28444
rect 21818 28432 21824 28444
rect 21876 28432 21882 28484
rect 15841 28407 15899 28413
rect 15841 28373 15853 28407
rect 15887 28373 15899 28407
rect 15841 28367 15899 28373
rect 16301 28407 16359 28413
rect 16301 28373 16313 28407
rect 16347 28404 16359 28407
rect 16850 28404 16856 28416
rect 16347 28376 16856 28404
rect 16347 28373 16359 28376
rect 16301 28367 16359 28373
rect 16850 28364 16856 28376
rect 16908 28364 16914 28416
rect 17310 28404 17316 28416
rect 17271 28376 17316 28404
rect 17310 28364 17316 28376
rect 17368 28364 17374 28416
rect 17957 28407 18015 28413
rect 17957 28373 17969 28407
rect 18003 28404 18015 28407
rect 18598 28404 18604 28416
rect 18003 28376 18604 28404
rect 18003 28373 18015 28376
rect 17957 28367 18015 28373
rect 18598 28364 18604 28376
rect 18656 28364 18662 28416
rect 19061 28407 19119 28413
rect 19061 28373 19073 28407
rect 19107 28404 19119 28407
rect 19610 28404 19616 28416
rect 19107 28376 19616 28404
rect 19107 28373 19119 28376
rect 19061 28367 19119 28373
rect 19610 28364 19616 28376
rect 19668 28364 19674 28416
rect 20714 28404 20720 28416
rect 20675 28376 20720 28404
rect 20714 28364 20720 28376
rect 20772 28364 20778 28416
rect 22186 28364 22192 28416
rect 22244 28404 22250 28416
rect 22465 28407 22523 28413
rect 22465 28404 22477 28407
rect 22244 28376 22477 28404
rect 22244 28364 22250 28376
rect 22465 28373 22477 28376
rect 22511 28373 22523 28407
rect 22465 28367 22523 28373
rect 27062 28364 27068 28416
rect 27120 28404 27126 28416
rect 27157 28407 27215 28413
rect 27157 28404 27169 28407
rect 27120 28376 27169 28404
rect 27120 28364 27126 28376
rect 27157 28373 27169 28376
rect 27203 28373 27215 28407
rect 27157 28367 27215 28373
rect 1104 28314 28060 28336
rect 1104 28262 9935 28314
rect 9987 28262 9999 28314
rect 10051 28262 10063 28314
rect 10115 28262 10127 28314
rect 10179 28262 10191 28314
rect 10243 28262 18920 28314
rect 18972 28262 18984 28314
rect 19036 28262 19048 28314
rect 19100 28262 19112 28314
rect 19164 28262 19176 28314
rect 19228 28262 28060 28314
rect 1104 28240 28060 28262
rect 4338 28200 4344 28212
rect 4299 28172 4344 28200
rect 4338 28160 4344 28172
rect 4396 28160 4402 28212
rect 5902 28160 5908 28212
rect 5960 28200 5966 28212
rect 5960 28172 6684 28200
rect 5960 28160 5966 28172
rect 4246 28092 4252 28144
rect 4304 28132 4310 28144
rect 6656 28132 6684 28172
rect 12802 28160 12808 28212
rect 12860 28200 12866 28212
rect 16114 28200 16120 28212
rect 12860 28172 16120 28200
rect 12860 28160 12866 28172
rect 16114 28160 16120 28172
rect 16172 28160 16178 28212
rect 7438 28135 7496 28141
rect 7438 28132 7450 28135
rect 4304 28104 6592 28132
rect 6656 28104 7450 28132
rect 4304 28092 4310 28104
rect 4448 28073 4476 28104
rect 2685 28067 2743 28073
rect 2685 28033 2697 28067
rect 2731 28064 2743 28067
rect 3145 28067 3203 28073
rect 3145 28064 3157 28067
rect 2731 28036 3157 28064
rect 2731 28033 2743 28036
rect 2685 28027 2743 28033
rect 3145 28033 3157 28036
rect 3191 28064 3203 28067
rect 4433 28067 4491 28073
rect 3191 28036 4384 28064
rect 3191 28033 3203 28036
rect 3145 28027 3203 28033
rect 2961 27863 3019 27869
rect 2961 27829 2973 27863
rect 3007 27860 3019 27863
rect 3878 27860 3884 27872
rect 3007 27832 3884 27860
rect 3007 27829 3019 27832
rect 2961 27823 3019 27829
rect 3878 27820 3884 27832
rect 3936 27820 3942 27872
rect 4356 27860 4384 28036
rect 4433 28033 4445 28067
rect 4479 28033 4491 28067
rect 4433 28027 4491 28033
rect 4700 28067 4758 28073
rect 4700 28033 4712 28067
rect 4746 28064 4758 28067
rect 5258 28064 5264 28076
rect 4746 28036 5264 28064
rect 4746 28033 4758 28036
rect 4700 28027 4758 28033
rect 5258 28024 5264 28036
rect 5316 28024 5322 28076
rect 6564 28008 6592 28104
rect 7438 28101 7450 28104
rect 7484 28101 7496 28135
rect 9674 28132 9680 28144
rect 7438 28095 7496 28101
rect 9600 28104 9680 28132
rect 9600 28073 9628 28104
rect 9674 28092 9680 28104
rect 9732 28092 9738 28144
rect 11900 28104 14320 28132
rect 9858 28073 9864 28076
rect 9585 28067 9643 28073
rect 9585 28033 9597 28067
rect 9631 28033 9643 28067
rect 9585 28027 9643 28033
rect 9852 28027 9864 28073
rect 9916 28064 9922 28076
rect 9916 28036 9952 28064
rect 9858 28024 9864 28027
rect 9916 28024 9922 28036
rect 6546 27956 6552 28008
rect 6604 27996 6610 28008
rect 7193 27999 7251 28005
rect 7193 27996 7205 27999
rect 6604 27968 7205 27996
rect 6604 27956 6610 27968
rect 7193 27965 7205 27968
rect 7239 27965 7251 27999
rect 7193 27959 7251 27965
rect 10962 27956 10968 28008
rect 11020 27996 11026 28008
rect 11900 28005 11928 28104
rect 12152 28067 12210 28073
rect 12152 28033 12164 28067
rect 12198 28064 12210 28067
rect 12526 28064 12532 28076
rect 12198 28036 12532 28064
rect 12198 28033 12210 28036
rect 12152 28027 12210 28033
rect 12526 28024 12532 28036
rect 12584 28024 12590 28076
rect 14292 28073 14320 28104
rect 16776 28104 18552 28132
rect 16776 28076 16804 28104
rect 14277 28067 14335 28073
rect 14277 28033 14289 28067
rect 14323 28033 14335 28067
rect 14533 28067 14591 28073
rect 14533 28064 14545 28067
rect 14277 28027 14335 28033
rect 14384 28036 14545 28064
rect 11885 27999 11943 28005
rect 11885 27996 11897 27999
rect 11020 27968 11897 27996
rect 11020 27956 11026 27968
rect 11885 27965 11897 27968
rect 11931 27965 11943 27999
rect 11885 27959 11943 27965
rect 13906 27956 13912 28008
rect 13964 27996 13970 28008
rect 14384 27996 14412 28036
rect 14533 28033 14545 28036
rect 14579 28033 14591 28067
rect 14533 28027 14591 28033
rect 16669 28067 16727 28073
rect 16669 28033 16681 28067
rect 16715 28064 16727 28067
rect 16758 28064 16764 28076
rect 16715 28036 16764 28064
rect 16715 28033 16727 28036
rect 16669 28027 16727 28033
rect 16758 28024 16764 28036
rect 16816 28024 16822 28076
rect 16942 28073 16948 28076
rect 16936 28064 16948 28073
rect 16903 28036 16948 28064
rect 16936 28027 16948 28036
rect 16942 28024 16948 28027
rect 17000 28024 17006 28076
rect 18524 28073 18552 28104
rect 19702 28092 19708 28144
rect 19760 28132 19766 28144
rect 19760 28104 27016 28132
rect 19760 28092 19766 28104
rect 18509 28067 18567 28073
rect 18509 28033 18521 28067
rect 18555 28033 18567 28067
rect 18509 28027 18567 28033
rect 18598 28024 18604 28076
rect 18656 28064 18662 28076
rect 18765 28067 18823 28073
rect 18765 28064 18777 28067
rect 18656 28036 18777 28064
rect 18656 28024 18662 28036
rect 18765 28033 18777 28036
rect 18811 28033 18823 28067
rect 18765 28027 18823 28033
rect 19610 28024 19616 28076
rect 19668 28064 19674 28076
rect 20533 28067 20591 28073
rect 20533 28064 20545 28067
rect 19668 28036 20545 28064
rect 19668 28024 19674 28036
rect 20533 28033 20545 28036
rect 20579 28033 20591 28067
rect 20533 28027 20591 28033
rect 21177 28067 21235 28073
rect 21177 28033 21189 28067
rect 21223 28064 21235 28067
rect 21223 28036 22094 28064
rect 21223 28033 21235 28036
rect 21177 28027 21235 28033
rect 13964 27968 14412 27996
rect 22066 27996 22094 28036
rect 22278 28024 22284 28076
rect 22336 28064 22342 28076
rect 22557 28067 22615 28073
rect 22557 28064 22569 28067
rect 22336 28036 22569 28064
rect 22336 28024 22342 28036
rect 22557 28033 22569 28036
rect 22603 28033 22615 28067
rect 22557 28027 22615 28033
rect 23290 28024 23296 28076
rect 23348 28064 23354 28076
rect 23845 28067 23903 28073
rect 23845 28064 23857 28067
rect 23348 28036 23857 28064
rect 23348 28024 23354 28036
rect 23845 28033 23857 28036
rect 23891 28033 23903 28067
rect 23845 28027 23903 28033
rect 26421 28067 26479 28073
rect 26421 28033 26433 28067
rect 26467 28064 26479 28067
rect 26878 28064 26884 28076
rect 26467 28036 26884 28064
rect 26467 28033 26479 28036
rect 26421 28027 26479 28033
rect 26878 28024 26884 28036
rect 26936 28024 26942 28076
rect 26988 28073 27016 28104
rect 26973 28067 27031 28073
rect 26973 28033 26985 28067
rect 27019 28033 27031 28067
rect 27154 28064 27160 28076
rect 27115 28036 27160 28064
rect 26973 28027 27031 28033
rect 27154 28024 27160 28036
rect 27212 28024 27218 28076
rect 27798 27996 27804 28008
rect 22066 27968 27804 27996
rect 13964 27956 13970 27968
rect 27798 27956 27804 27968
rect 27856 27956 27862 28008
rect 6822 27928 6828 27940
rect 5368 27900 6828 27928
rect 5368 27860 5396 27900
rect 6822 27888 6828 27900
rect 6880 27888 6886 27940
rect 25866 27888 25872 27940
rect 25924 27928 25930 27940
rect 26973 27931 27031 27937
rect 26973 27928 26985 27931
rect 25924 27900 26985 27928
rect 25924 27888 25930 27900
rect 26973 27897 26985 27900
rect 27019 27897 27031 27931
rect 26973 27891 27031 27897
rect 5810 27860 5816 27872
rect 4356 27832 5396 27860
rect 5771 27832 5816 27860
rect 5810 27820 5816 27832
rect 5868 27820 5874 27872
rect 8570 27860 8576 27872
rect 8483 27832 8576 27860
rect 8570 27820 8576 27832
rect 8628 27860 8634 27872
rect 9214 27860 9220 27872
rect 8628 27832 9220 27860
rect 8628 27820 8634 27832
rect 9214 27820 9220 27832
rect 9272 27820 9278 27872
rect 10686 27820 10692 27872
rect 10744 27860 10750 27872
rect 10965 27863 11023 27869
rect 10965 27860 10977 27863
rect 10744 27832 10977 27860
rect 10744 27820 10750 27832
rect 10965 27829 10977 27832
rect 11011 27829 11023 27863
rect 10965 27823 11023 27829
rect 13170 27820 13176 27872
rect 13228 27860 13234 27872
rect 13265 27863 13323 27869
rect 13265 27860 13277 27863
rect 13228 27832 13277 27860
rect 13228 27820 13234 27832
rect 13265 27829 13277 27832
rect 13311 27829 13323 27863
rect 13265 27823 13323 27829
rect 13538 27820 13544 27872
rect 13596 27860 13602 27872
rect 15286 27860 15292 27872
rect 13596 27832 15292 27860
rect 13596 27820 13602 27832
rect 15286 27820 15292 27832
rect 15344 27860 15350 27872
rect 15657 27863 15715 27869
rect 15657 27860 15669 27863
rect 15344 27832 15669 27860
rect 15344 27820 15350 27832
rect 15657 27829 15669 27832
rect 15703 27829 15715 27863
rect 18046 27860 18052 27872
rect 18007 27832 18052 27860
rect 15657 27823 15715 27829
rect 18046 27820 18052 27832
rect 18104 27820 18110 27872
rect 19426 27820 19432 27872
rect 19484 27860 19490 27872
rect 19889 27863 19947 27869
rect 19889 27860 19901 27863
rect 19484 27832 19901 27860
rect 19484 27820 19490 27832
rect 19889 27829 19901 27832
rect 19935 27829 19947 27863
rect 20346 27860 20352 27872
rect 20307 27832 20352 27860
rect 19889 27823 19947 27829
rect 20346 27820 20352 27832
rect 20404 27820 20410 27872
rect 20990 27860 20996 27872
rect 20951 27832 20996 27860
rect 20990 27820 20996 27832
rect 21048 27820 21054 27872
rect 22370 27860 22376 27872
rect 22331 27832 22376 27860
rect 22370 27820 22376 27832
rect 22428 27820 22434 27872
rect 22738 27820 22744 27872
rect 22796 27860 22802 27872
rect 23290 27860 23296 27872
rect 22796 27832 23296 27860
rect 22796 27820 22802 27832
rect 23290 27820 23296 27832
rect 23348 27820 23354 27872
rect 23661 27863 23719 27869
rect 23661 27829 23673 27863
rect 23707 27860 23719 27863
rect 23842 27860 23848 27872
rect 23707 27832 23848 27860
rect 23707 27829 23719 27832
rect 23661 27823 23719 27829
rect 23842 27820 23848 27832
rect 23900 27820 23906 27872
rect 26237 27863 26295 27869
rect 26237 27829 26249 27863
rect 26283 27860 26295 27863
rect 26602 27860 26608 27872
rect 26283 27832 26608 27860
rect 26283 27829 26295 27832
rect 26237 27823 26295 27829
rect 26602 27820 26608 27832
rect 26660 27820 26666 27872
rect 1104 27770 28060 27792
rect 1104 27718 5442 27770
rect 5494 27718 5506 27770
rect 5558 27718 5570 27770
rect 5622 27718 5634 27770
rect 5686 27718 5698 27770
rect 5750 27718 14428 27770
rect 14480 27718 14492 27770
rect 14544 27718 14556 27770
rect 14608 27718 14620 27770
rect 14672 27718 14684 27770
rect 14736 27718 23413 27770
rect 23465 27718 23477 27770
rect 23529 27718 23541 27770
rect 23593 27718 23605 27770
rect 23657 27718 23669 27770
rect 23721 27718 28060 27770
rect 1104 27696 28060 27718
rect 6638 27656 6644 27668
rect 3988 27628 4476 27656
rect 1765 27591 1823 27597
rect 1765 27557 1777 27591
rect 1811 27588 1823 27591
rect 3988 27588 4016 27628
rect 4338 27588 4344 27600
rect 1811 27560 4016 27588
rect 4080 27560 4344 27588
rect 1811 27557 1823 27560
rect 1765 27551 1823 27557
rect 4080 27520 4108 27560
rect 4338 27548 4344 27560
rect 4396 27548 4402 27600
rect 4448 27588 4476 27628
rect 6472 27628 6644 27656
rect 5442 27588 5448 27600
rect 4448 27560 5448 27588
rect 5442 27548 5448 27560
rect 5500 27548 5506 27600
rect 5534 27548 5540 27600
rect 5592 27588 5598 27600
rect 5810 27588 5816 27600
rect 5592 27560 5816 27588
rect 5592 27548 5598 27560
rect 5810 27548 5816 27560
rect 5868 27588 5874 27600
rect 6472 27588 6500 27628
rect 6638 27616 6644 27628
rect 6696 27616 6702 27668
rect 9674 27656 9680 27668
rect 8956 27628 9680 27656
rect 5868 27560 6500 27588
rect 5868 27548 5874 27560
rect 1964 27492 4108 27520
rect 1964 27461 1992 27492
rect 4154 27480 4160 27532
rect 4212 27520 4218 27532
rect 4433 27523 4491 27529
rect 4433 27520 4445 27523
rect 4212 27492 4445 27520
rect 4212 27480 4218 27492
rect 4433 27489 4445 27492
rect 4479 27520 4491 27523
rect 4982 27520 4988 27532
rect 4479 27492 4988 27520
rect 4479 27489 4491 27492
rect 4433 27483 4491 27489
rect 4982 27480 4988 27492
rect 5040 27480 5046 27532
rect 6472 27520 6500 27560
rect 6472 27492 6592 27520
rect 1949 27455 2007 27461
rect 1949 27421 1961 27455
rect 1995 27421 2007 27455
rect 2590 27452 2596 27464
rect 2551 27424 2596 27452
rect 1949 27415 2007 27421
rect 2590 27412 2596 27424
rect 2648 27412 2654 27464
rect 3237 27455 3295 27461
rect 3237 27421 3249 27455
rect 3283 27452 3295 27455
rect 3694 27452 3700 27464
rect 3283 27424 3700 27452
rect 3283 27421 3295 27424
rect 3237 27415 3295 27421
rect 3694 27412 3700 27424
rect 3752 27412 3758 27464
rect 4525 27455 4583 27461
rect 4525 27421 4537 27455
rect 4571 27421 4583 27455
rect 4706 27452 4712 27464
rect 4667 27424 4712 27452
rect 4525 27415 4583 27421
rect 4540 27384 4568 27415
rect 4706 27412 4712 27424
rect 4764 27412 4770 27464
rect 5353 27455 5411 27461
rect 5353 27421 5365 27455
rect 5399 27452 5411 27455
rect 5813 27455 5871 27461
rect 5813 27452 5825 27455
rect 5399 27424 5825 27452
rect 5399 27421 5411 27424
rect 5353 27415 5411 27421
rect 5813 27421 5825 27424
rect 5859 27452 5871 27455
rect 5994 27452 6000 27464
rect 5859 27424 6000 27452
rect 5859 27421 5871 27424
rect 5813 27415 5871 27421
rect 5994 27412 6000 27424
rect 6052 27412 6058 27464
rect 6454 27452 6460 27464
rect 6415 27424 6460 27452
rect 6454 27412 6460 27424
rect 6512 27412 6518 27464
rect 6564 27452 6592 27492
rect 8110 27452 8116 27464
rect 6564 27424 8116 27452
rect 8110 27412 8116 27424
rect 8168 27412 8174 27464
rect 8956 27461 8984 27628
rect 9674 27616 9680 27628
rect 9732 27656 9738 27668
rect 10962 27656 10968 27668
rect 9732 27628 10968 27656
rect 9732 27616 9738 27628
rect 10962 27616 10968 27628
rect 11020 27616 11026 27668
rect 12989 27659 13047 27665
rect 12989 27625 13001 27659
rect 13035 27656 13047 27659
rect 13078 27656 13084 27668
rect 13035 27628 13084 27656
rect 13035 27625 13047 27628
rect 12989 27619 13047 27625
rect 13078 27616 13084 27628
rect 13136 27616 13142 27668
rect 18138 27616 18144 27668
rect 18196 27656 18202 27668
rect 18693 27659 18751 27665
rect 18693 27656 18705 27659
rect 18196 27628 18705 27656
rect 18196 27616 18202 27628
rect 18693 27625 18705 27628
rect 18739 27625 18751 27659
rect 18693 27619 18751 27625
rect 21634 27616 21640 27668
rect 21692 27656 21698 27668
rect 21729 27659 21787 27665
rect 21729 27656 21741 27659
rect 21692 27628 21741 27656
rect 21692 27616 21698 27628
rect 21729 27625 21741 27628
rect 21775 27625 21787 27659
rect 21729 27619 21787 27625
rect 21818 27616 21824 27668
rect 21876 27656 21882 27668
rect 27614 27656 27620 27668
rect 21876 27628 27620 27656
rect 21876 27616 21882 27628
rect 27614 27616 27620 27628
rect 27672 27616 27678 27668
rect 13265 27591 13323 27597
rect 13265 27557 13277 27591
rect 13311 27588 13323 27591
rect 13906 27588 13912 27600
rect 13311 27560 13912 27588
rect 13311 27557 13323 27560
rect 13265 27551 13323 27557
rect 13906 27548 13912 27560
rect 13964 27548 13970 27600
rect 15933 27591 15991 27597
rect 15933 27557 15945 27591
rect 15979 27588 15991 27591
rect 18230 27588 18236 27600
rect 15979 27560 18236 27588
rect 15979 27557 15991 27560
rect 15933 27551 15991 27557
rect 18230 27548 18236 27560
rect 18288 27548 18294 27600
rect 23293 27591 23351 27597
rect 23293 27557 23305 27591
rect 23339 27588 23351 27591
rect 25222 27588 25228 27600
rect 23339 27560 25228 27588
rect 23339 27557 23351 27560
rect 23293 27551 23351 27557
rect 25222 27548 25228 27560
rect 25280 27548 25286 27600
rect 27154 27548 27160 27600
rect 27212 27548 27218 27600
rect 13173 27523 13231 27529
rect 13173 27520 13185 27523
rect 12084 27492 13185 27520
rect 8941 27455 8999 27461
rect 8941 27421 8953 27455
rect 8987 27421 8999 27455
rect 8941 27415 8999 27421
rect 9208 27455 9266 27461
rect 9208 27421 9220 27455
rect 9254 27421 9266 27455
rect 9208 27415 9266 27421
rect 5166 27384 5172 27396
rect 4540 27356 5172 27384
rect 5166 27344 5172 27356
rect 5224 27344 5230 27396
rect 6362 27344 6368 27396
rect 6420 27384 6426 27396
rect 6702 27387 6760 27393
rect 6702 27384 6714 27387
rect 6420 27356 6714 27384
rect 6420 27344 6426 27356
rect 6702 27353 6714 27356
rect 6748 27353 6760 27387
rect 6702 27347 6760 27353
rect 9122 27344 9128 27396
rect 9180 27384 9186 27396
rect 9232 27384 9260 27415
rect 10962 27412 10968 27464
rect 11020 27452 11026 27464
rect 11057 27455 11115 27461
rect 11057 27452 11069 27455
rect 11020 27424 11069 27452
rect 11020 27412 11026 27424
rect 11057 27421 11069 27424
rect 11103 27421 11115 27455
rect 11057 27415 11115 27421
rect 11146 27412 11152 27464
rect 11204 27452 11210 27464
rect 11313 27455 11371 27461
rect 11313 27452 11325 27455
rect 11204 27424 11325 27452
rect 11204 27412 11210 27424
rect 11313 27421 11325 27424
rect 11359 27421 11371 27455
rect 11313 27415 11371 27421
rect 12084 27384 12112 27492
rect 13173 27489 13185 27492
rect 13219 27489 13231 27523
rect 13998 27520 14004 27532
rect 13173 27483 13231 27489
rect 13648 27492 14004 27520
rect 12897 27455 12955 27461
rect 12897 27421 12909 27455
rect 12943 27421 12955 27455
rect 13538 27452 13544 27464
rect 13499 27424 13544 27452
rect 12897 27415 12955 27421
rect 9180 27356 9260 27384
rect 9324 27356 12112 27384
rect 12912 27384 12940 27415
rect 13538 27412 13544 27424
rect 13596 27412 13602 27464
rect 13648 27461 13676 27492
rect 13998 27480 14004 27492
rect 14056 27480 14062 27532
rect 18325 27523 18383 27529
rect 18325 27489 18337 27523
rect 18371 27520 18383 27523
rect 18690 27520 18696 27532
rect 18371 27492 18696 27520
rect 18371 27489 18383 27492
rect 18325 27483 18383 27489
rect 18690 27480 18696 27492
rect 18748 27480 18754 27532
rect 21818 27520 21824 27532
rect 21008 27492 21824 27520
rect 13633 27455 13691 27461
rect 13633 27421 13645 27455
rect 13679 27421 13691 27455
rect 13633 27415 13691 27421
rect 13725 27455 13783 27461
rect 13725 27421 13737 27455
rect 13771 27452 13783 27455
rect 13814 27452 13820 27464
rect 13771 27424 13820 27452
rect 13771 27421 13783 27424
rect 13725 27415 13783 27421
rect 13814 27412 13820 27424
rect 13872 27412 13878 27464
rect 13906 27412 13912 27464
rect 13964 27452 13970 27464
rect 15381 27455 15439 27461
rect 15381 27452 15393 27455
rect 13964 27424 14009 27452
rect 14936 27424 15393 27452
rect 13964 27412 13970 27424
rect 14090 27384 14096 27396
rect 12912 27356 14096 27384
rect 9180 27344 9186 27356
rect 2409 27319 2467 27325
rect 2409 27285 2421 27319
rect 2455 27316 2467 27319
rect 2498 27316 2504 27328
rect 2455 27288 2504 27316
rect 2455 27285 2467 27288
rect 2409 27279 2467 27285
rect 2498 27276 2504 27288
rect 2556 27276 2562 27328
rect 3050 27316 3056 27328
rect 3011 27288 3056 27316
rect 3050 27276 3056 27288
rect 3108 27276 3114 27328
rect 3694 27276 3700 27328
rect 3752 27316 3758 27328
rect 3973 27319 4031 27325
rect 3973 27316 3985 27319
rect 3752 27288 3985 27316
rect 3752 27276 3758 27288
rect 3973 27285 3985 27288
rect 4019 27285 4031 27319
rect 3973 27279 4031 27285
rect 4338 27276 4344 27328
rect 4396 27316 4402 27328
rect 4617 27319 4675 27325
rect 4617 27316 4629 27319
rect 4396 27288 4629 27316
rect 4396 27276 4402 27288
rect 4617 27285 4629 27288
rect 4663 27285 4675 27319
rect 4617 27279 4675 27285
rect 5629 27319 5687 27325
rect 5629 27285 5641 27319
rect 5675 27316 5687 27319
rect 6822 27316 6828 27328
rect 5675 27288 6828 27316
rect 5675 27285 5687 27288
rect 5629 27279 5687 27285
rect 6822 27276 6828 27288
rect 6880 27276 6886 27328
rect 7834 27316 7840 27328
rect 7795 27288 7840 27316
rect 7834 27276 7840 27288
rect 7892 27276 7898 27328
rect 8018 27276 8024 27328
rect 8076 27316 8082 27328
rect 9324 27316 9352 27356
rect 14090 27344 14096 27356
rect 14148 27344 14154 27396
rect 14936 27328 14964 27424
rect 15381 27421 15393 27424
rect 15427 27421 15439 27455
rect 15381 27415 15439 27421
rect 15841 27455 15899 27461
rect 15841 27421 15853 27455
rect 15887 27452 15899 27455
rect 16022 27452 16028 27464
rect 15887 27424 16028 27452
rect 15887 27421 15899 27424
rect 15841 27415 15899 27421
rect 16022 27412 16028 27424
rect 16080 27412 16086 27464
rect 16117 27455 16175 27461
rect 16117 27421 16129 27455
rect 16163 27452 16175 27455
rect 17405 27455 17463 27461
rect 16163 27424 16528 27452
rect 16163 27421 16175 27424
rect 16117 27415 16175 27421
rect 10318 27316 10324 27328
rect 8076 27288 9352 27316
rect 10279 27288 10324 27316
rect 8076 27276 8082 27288
rect 10318 27276 10324 27288
rect 10376 27276 10382 27328
rect 12434 27276 12440 27328
rect 12492 27316 12498 27328
rect 12492 27288 12537 27316
rect 12492 27276 12498 27288
rect 12710 27276 12716 27328
rect 12768 27316 12774 27328
rect 13173 27319 13231 27325
rect 13173 27316 13185 27319
rect 12768 27288 13185 27316
rect 12768 27276 12774 27288
rect 13173 27285 13185 27288
rect 13219 27285 13231 27319
rect 14918 27316 14924 27328
rect 14879 27288 14924 27316
rect 13173 27279 13231 27285
rect 14918 27276 14924 27288
rect 14976 27276 14982 27328
rect 15194 27316 15200 27328
rect 15155 27288 15200 27316
rect 15194 27276 15200 27288
rect 15252 27276 15258 27328
rect 15654 27316 15660 27328
rect 15615 27288 15660 27316
rect 15654 27276 15660 27288
rect 15712 27276 15718 27328
rect 16500 27325 16528 27424
rect 17405 27421 17417 27455
rect 17451 27421 17463 27455
rect 18506 27452 18512 27464
rect 18467 27424 18512 27452
rect 17405 27415 17463 27421
rect 16945 27387 17003 27393
rect 16945 27353 16957 27387
rect 16991 27384 17003 27387
rect 17126 27384 17132 27396
rect 16991 27356 17132 27384
rect 16991 27353 17003 27356
rect 16945 27347 17003 27353
rect 17126 27344 17132 27356
rect 17184 27384 17190 27396
rect 17420 27384 17448 27415
rect 18506 27412 18512 27424
rect 18564 27412 18570 27464
rect 19245 27455 19303 27461
rect 19245 27421 19257 27455
rect 19291 27452 19303 27455
rect 19886 27452 19892 27464
rect 19291 27424 19892 27452
rect 19291 27421 19303 27424
rect 19245 27415 19303 27421
rect 19886 27412 19892 27424
rect 19944 27452 19950 27464
rect 21008 27452 21036 27492
rect 21818 27480 21824 27492
rect 21876 27480 21882 27532
rect 23198 27480 23204 27532
rect 23256 27520 23262 27532
rect 27172 27520 27200 27548
rect 23256 27492 27200 27520
rect 23256 27480 23262 27492
rect 19944 27424 21036 27452
rect 19944 27412 19950 27424
rect 21174 27412 21180 27464
rect 21232 27452 21238 27464
rect 22094 27461 22100 27464
rect 21361 27455 21419 27461
rect 21361 27452 21373 27455
rect 21232 27424 21373 27452
rect 21232 27412 21238 27424
rect 21361 27421 21373 27424
rect 21407 27421 21419 27455
rect 21361 27415 21419 27421
rect 21545 27455 21603 27461
rect 21545 27421 21557 27455
rect 21591 27421 21603 27455
rect 21545 27415 21603 27421
rect 22088 27415 22100 27461
rect 22152 27452 22158 27464
rect 23492 27461 23520 27492
rect 23293 27455 23351 27461
rect 23293 27452 23305 27455
rect 22152 27424 22188 27452
rect 22572 27424 23305 27452
rect 17184 27356 17448 27384
rect 19512 27387 19570 27393
rect 17184 27344 17190 27356
rect 19512 27353 19524 27387
rect 19558 27384 19570 27387
rect 20346 27384 20352 27396
rect 19558 27356 20352 27384
rect 19558 27353 19570 27356
rect 19512 27347 19570 27353
rect 20346 27344 20352 27356
rect 20404 27344 20410 27396
rect 21560 27384 21588 27415
rect 22094 27412 22100 27415
rect 22152 27412 22158 27424
rect 22462 27384 22468 27396
rect 21560 27356 22468 27384
rect 22462 27344 22468 27356
rect 22520 27344 22526 27396
rect 16485 27319 16543 27325
rect 16485 27285 16497 27319
rect 16531 27316 16543 27319
rect 16574 27316 16580 27328
rect 16531 27288 16580 27316
rect 16531 27285 16543 27288
rect 16485 27279 16543 27285
rect 16574 27276 16580 27288
rect 16632 27276 16638 27328
rect 17034 27276 17040 27328
rect 17092 27316 17098 27328
rect 17221 27319 17279 27325
rect 17221 27316 17233 27319
rect 17092 27288 17233 27316
rect 17092 27276 17098 27288
rect 17221 27285 17233 27288
rect 17267 27285 17279 27319
rect 17221 27279 17279 27285
rect 20070 27276 20076 27328
rect 20128 27316 20134 27328
rect 20625 27319 20683 27325
rect 20625 27316 20637 27319
rect 20128 27288 20637 27316
rect 20128 27276 20134 27288
rect 20625 27285 20637 27288
rect 20671 27285 20683 27319
rect 20625 27279 20683 27285
rect 21542 27276 21548 27328
rect 21600 27316 21606 27328
rect 22572 27316 22600 27424
rect 23293 27421 23305 27424
rect 23339 27421 23351 27455
rect 23293 27415 23351 27421
rect 23477 27455 23535 27461
rect 23477 27421 23489 27455
rect 23523 27421 23535 27455
rect 23477 27415 23535 27421
rect 23308 27384 23336 27415
rect 23750 27412 23756 27464
rect 23808 27452 23814 27464
rect 23845 27455 23903 27461
rect 23845 27452 23857 27455
rect 23808 27424 23857 27452
rect 23808 27412 23814 27424
rect 23845 27421 23857 27424
rect 23891 27421 23903 27455
rect 24578 27452 24584 27464
rect 24539 27424 24584 27452
rect 23845 27415 23903 27421
rect 24578 27412 24584 27424
rect 24636 27412 24642 27464
rect 25225 27455 25283 27461
rect 25225 27421 25237 27455
rect 25271 27421 25283 27455
rect 25225 27415 25283 27421
rect 25961 27455 26019 27461
rect 25961 27421 25973 27455
rect 26007 27452 26019 27455
rect 26050 27452 26056 27464
rect 26007 27424 26056 27452
rect 26007 27421 26019 27424
rect 25961 27415 26019 27421
rect 24210 27384 24216 27396
rect 23308 27356 24216 27384
rect 24210 27344 24216 27356
rect 24268 27344 24274 27396
rect 24302 27344 24308 27396
rect 24360 27384 24366 27396
rect 25240 27384 25268 27415
rect 26050 27412 26056 27424
rect 26108 27412 26114 27464
rect 26605 27455 26663 27461
rect 26605 27421 26617 27455
rect 26651 27452 26663 27455
rect 26970 27452 26976 27464
rect 26651 27424 26976 27452
rect 26651 27421 26663 27424
rect 26605 27415 26663 27421
rect 26970 27412 26976 27424
rect 27028 27412 27034 27464
rect 27065 27455 27123 27461
rect 27065 27421 27077 27455
rect 27111 27452 27123 27455
rect 27154 27452 27160 27464
rect 27111 27424 27160 27452
rect 27111 27421 27123 27424
rect 27065 27415 27123 27421
rect 27154 27412 27160 27424
rect 27212 27412 27218 27464
rect 24360 27356 25268 27384
rect 24360 27344 24366 27356
rect 21600 27288 22600 27316
rect 21600 27276 21606 27288
rect 23014 27276 23020 27328
rect 23072 27316 23078 27328
rect 23201 27319 23259 27325
rect 23201 27316 23213 27319
rect 23072 27288 23213 27316
rect 23072 27276 23078 27288
rect 23201 27285 23213 27288
rect 23247 27285 23259 27319
rect 23201 27279 23259 27285
rect 23661 27319 23719 27325
rect 23661 27285 23673 27319
rect 23707 27316 23719 27319
rect 23934 27316 23940 27328
rect 23707 27288 23940 27316
rect 23707 27285 23719 27288
rect 23661 27279 23719 27285
rect 23934 27276 23940 27288
rect 23992 27276 23998 27328
rect 24397 27319 24455 27325
rect 24397 27285 24409 27319
rect 24443 27316 24455 27319
rect 24486 27316 24492 27328
rect 24443 27288 24492 27316
rect 24443 27285 24455 27288
rect 24397 27279 24455 27285
rect 24486 27276 24492 27288
rect 24544 27276 24550 27328
rect 25041 27319 25099 27325
rect 25041 27285 25053 27319
rect 25087 27316 25099 27319
rect 25130 27316 25136 27328
rect 25087 27288 25136 27316
rect 25087 27285 25099 27288
rect 25041 27279 25099 27285
rect 25130 27276 25136 27288
rect 25188 27276 25194 27328
rect 25774 27316 25780 27328
rect 25735 27288 25780 27316
rect 25774 27276 25780 27288
rect 25832 27276 25838 27328
rect 26326 27276 26332 27328
rect 26384 27316 26390 27328
rect 26421 27319 26479 27325
rect 26421 27316 26433 27319
rect 26384 27288 26433 27316
rect 26384 27276 26390 27288
rect 26421 27285 26433 27288
rect 26467 27285 26479 27319
rect 27246 27316 27252 27328
rect 27207 27288 27252 27316
rect 26421 27279 26479 27285
rect 27246 27276 27252 27288
rect 27304 27276 27310 27328
rect 1104 27226 28060 27248
rect 1104 27174 9935 27226
rect 9987 27174 9999 27226
rect 10051 27174 10063 27226
rect 10115 27174 10127 27226
rect 10179 27174 10191 27226
rect 10243 27174 18920 27226
rect 18972 27174 18984 27226
rect 19036 27174 19048 27226
rect 19100 27174 19112 27226
rect 19164 27174 19176 27226
rect 19228 27174 28060 27226
rect 1104 27152 28060 27174
rect 2590 27072 2596 27124
rect 2648 27112 2654 27124
rect 4062 27112 4068 27124
rect 2648 27084 4068 27112
rect 2648 27072 2654 27084
rect 4062 27072 4068 27084
rect 4120 27072 4126 27124
rect 4154 27072 4160 27124
rect 4212 27112 4218 27124
rect 5258 27112 5264 27124
rect 4212 27084 4844 27112
rect 5219 27084 5264 27112
rect 4212 27072 4218 27084
rect 3329 27047 3387 27053
rect 3329 27044 3341 27047
rect 1596 27016 3341 27044
rect 1394 26936 1400 26988
rect 1452 26976 1458 26988
rect 1596 26985 1624 27016
rect 3329 27013 3341 27016
rect 3375 27013 3387 27047
rect 4246 27044 4252 27056
rect 3329 27007 3387 27013
rect 3804 27016 4252 27044
rect 1581 26979 1639 26985
rect 1581 26976 1593 26979
rect 1452 26948 1593 26976
rect 1452 26936 1458 26948
rect 1581 26945 1593 26948
rect 1627 26945 1639 26979
rect 1581 26939 1639 26945
rect 2317 26979 2375 26985
rect 2317 26945 2329 26979
rect 2363 26976 2375 26979
rect 2866 26976 2872 26988
rect 2363 26948 2872 26976
rect 2363 26945 2375 26948
rect 2317 26939 2375 26945
rect 2866 26936 2872 26948
rect 2924 26936 2930 26988
rect 3804 26985 3832 27016
rect 4246 27004 4252 27016
rect 4304 27004 4310 27056
rect 3789 26979 3847 26985
rect 3789 26945 3801 26979
rect 3835 26945 3847 26979
rect 3789 26939 3847 26945
rect 4056 26979 4114 26985
rect 4056 26945 4068 26979
rect 4102 26976 4114 26979
rect 4522 26976 4528 26988
rect 4102 26948 4528 26976
rect 4102 26945 4114 26948
rect 4056 26939 4114 26945
rect 1854 26868 1860 26920
rect 1912 26908 1918 26920
rect 3804 26908 3832 26939
rect 4522 26936 4528 26948
rect 4580 26936 4586 26988
rect 1912 26880 3832 26908
rect 4816 26908 4844 27084
rect 5258 27072 5264 27084
rect 5316 27072 5322 27124
rect 5810 27072 5816 27124
rect 5868 27072 5874 27124
rect 6362 27112 6368 27124
rect 6323 27084 6368 27112
rect 6362 27072 6368 27084
rect 6420 27072 6426 27124
rect 7006 27112 7012 27124
rect 6564 27084 7012 27112
rect 5534 26976 5540 26988
rect 5495 26948 5540 26976
rect 5534 26936 5540 26948
rect 5592 26936 5598 26988
rect 5626 26979 5684 26985
rect 5626 26945 5638 26979
rect 5672 26945 5684 26979
rect 5626 26939 5684 26945
rect 5726 26979 5784 26985
rect 5726 26945 5738 26979
rect 5772 26976 5784 26979
rect 5828 26976 5856 27072
rect 5772 26948 5856 26976
rect 5905 26979 5963 26985
rect 5772 26945 5784 26948
rect 5726 26939 5784 26945
rect 5905 26945 5917 26979
rect 5951 26976 5963 26979
rect 6086 26976 6092 26988
rect 5951 26948 6092 26976
rect 5951 26945 5963 26948
rect 5905 26939 5963 26945
rect 5641 26908 5669 26939
rect 6086 26936 6092 26948
rect 6144 26936 6150 26988
rect 6564 26979 6592 27084
rect 7006 27072 7012 27084
rect 7064 27112 7070 27124
rect 8159 27115 8217 27121
rect 8159 27112 8171 27115
rect 7064 27084 8171 27112
rect 7064 27072 7070 27084
rect 8159 27081 8171 27084
rect 8205 27081 8217 27115
rect 8159 27075 8217 27081
rect 11330 27072 11336 27124
rect 11388 27112 11394 27124
rect 11885 27115 11943 27121
rect 11885 27112 11897 27115
rect 11388 27084 11897 27112
rect 11388 27072 11394 27084
rect 11885 27081 11897 27084
rect 11931 27081 11943 27115
rect 12526 27112 12532 27124
rect 12487 27084 12532 27112
rect 11885 27075 11943 27081
rect 12526 27072 12532 27084
rect 12584 27072 12590 27124
rect 15654 27072 15660 27124
rect 15712 27112 15718 27124
rect 15712 27084 16804 27112
rect 15712 27072 15718 27084
rect 7282 27044 7288 27056
rect 6932 27016 7288 27044
rect 6846 26985 6904 26991
rect 6641 26979 6699 26985
rect 6564 26951 6653 26979
rect 6641 26945 6653 26951
rect 6687 26945 6699 26979
rect 6641 26939 6699 26945
rect 6733 26979 6791 26985
rect 6733 26945 6745 26979
rect 6779 26945 6791 26979
rect 6846 26951 6858 26985
rect 6892 26982 6904 26985
rect 6932 26982 6960 27016
rect 7282 27004 7288 27016
rect 7340 27004 7346 27056
rect 7558 27004 7564 27056
rect 7616 27044 7622 27056
rect 10870 27044 10876 27056
rect 7616 27016 10876 27044
rect 7616 27004 7622 27016
rect 10870 27004 10876 27016
rect 10928 27004 10934 27056
rect 12894 27044 12900 27056
rect 12820 27016 12900 27044
rect 6892 26954 6960 26982
rect 7009 26979 7067 26985
rect 6892 26951 6904 26954
rect 6846 26945 6904 26951
rect 7009 26945 7021 26979
rect 7055 26976 7067 26979
rect 7190 26976 7196 26988
rect 7055 26948 7196 26976
rect 7055 26945 7067 26948
rect 6733 26939 6791 26945
rect 7009 26939 7067 26945
rect 6178 26908 6184 26920
rect 4816 26880 6184 26908
rect 1912 26868 1918 26880
rect 6178 26868 6184 26880
rect 6236 26868 6242 26920
rect 6748 26908 6776 26939
rect 7190 26936 7196 26948
rect 7248 26976 7254 26988
rect 8570 26976 8576 26988
rect 7248 26948 8576 26976
rect 7248 26936 7254 26948
rect 8570 26936 8576 26948
rect 8628 26936 8634 26988
rect 9214 26976 9220 26988
rect 9175 26948 9220 26976
rect 9214 26936 9220 26948
rect 9272 26936 9278 26988
rect 9398 26936 9404 26988
rect 9456 26976 9462 26988
rect 10137 26979 10195 26985
rect 10137 26976 10149 26979
rect 9456 26948 10149 26976
rect 9456 26936 9462 26948
rect 10137 26945 10149 26948
rect 10183 26976 10195 26979
rect 10686 26976 10692 26988
rect 10183 26948 10692 26976
rect 10183 26945 10195 26948
rect 10137 26939 10195 26945
rect 10686 26936 10692 26948
rect 10744 26936 10750 26988
rect 11514 26976 11520 26988
rect 11475 26948 11520 26976
rect 11514 26936 11520 26948
rect 11572 26936 11578 26988
rect 11701 26979 11759 26985
rect 11701 26945 11713 26979
rect 11747 26945 11759 26979
rect 12710 26976 12716 26988
rect 12671 26948 12716 26976
rect 11701 26939 11759 26945
rect 7466 26908 7472 26920
rect 6748 26880 7472 26908
rect 7466 26868 7472 26880
rect 7524 26868 7530 26920
rect 7834 26868 7840 26920
rect 7892 26908 7898 26920
rect 7929 26911 7987 26917
rect 7929 26908 7941 26911
rect 7892 26880 7941 26908
rect 7892 26868 7898 26880
rect 7929 26877 7941 26880
rect 7975 26877 7987 26911
rect 7929 26871 7987 26877
rect 2133 26843 2191 26849
rect 2133 26809 2145 26843
rect 2179 26840 2191 26843
rect 7558 26840 7564 26852
rect 2179 26812 3832 26840
rect 2179 26809 2191 26812
rect 2133 26803 2191 26809
rect 1397 26775 1455 26781
rect 1397 26741 1409 26775
rect 1443 26772 1455 26775
rect 1670 26772 1676 26784
rect 1443 26744 1676 26772
rect 1443 26741 1455 26744
rect 1397 26735 1455 26741
rect 1670 26732 1676 26744
rect 1728 26732 1734 26784
rect 2685 26775 2743 26781
rect 2685 26741 2697 26775
rect 2731 26772 2743 26775
rect 2866 26772 2872 26784
rect 2731 26744 2872 26772
rect 2731 26741 2743 26744
rect 2685 26735 2743 26741
rect 2866 26732 2872 26744
rect 2924 26772 2930 26784
rect 2961 26775 3019 26781
rect 2961 26772 2973 26775
rect 2924 26744 2973 26772
rect 2924 26732 2930 26744
rect 2961 26741 2973 26744
rect 3007 26741 3019 26775
rect 3804 26772 3832 26812
rect 4816 26812 7564 26840
rect 4816 26772 4844 26812
rect 7558 26800 7564 26812
rect 7616 26800 7622 26852
rect 7944 26840 7972 26871
rect 8110 26868 8116 26920
rect 8168 26908 8174 26920
rect 9309 26911 9367 26917
rect 9309 26908 9321 26911
rect 8168 26880 9321 26908
rect 8168 26868 8174 26880
rect 9309 26877 9321 26880
rect 9355 26877 9367 26911
rect 9309 26871 9367 26877
rect 10413 26911 10471 26917
rect 10413 26877 10425 26911
rect 10459 26908 10471 26911
rect 10594 26908 10600 26920
rect 10459 26880 10600 26908
rect 10459 26877 10471 26880
rect 10413 26871 10471 26877
rect 10594 26868 10600 26880
rect 10652 26868 10658 26920
rect 11422 26868 11428 26920
rect 11480 26908 11486 26920
rect 11716 26908 11744 26939
rect 12710 26936 12716 26948
rect 12768 26936 12774 26988
rect 12820 26985 12848 27016
rect 12894 27004 12900 27016
rect 12952 27044 12958 27056
rect 16776 27044 16804 27084
rect 18506 27072 18512 27124
rect 18564 27112 18570 27124
rect 19061 27115 19119 27121
rect 19061 27112 19073 27115
rect 18564 27084 19073 27112
rect 18564 27072 18570 27084
rect 19061 27081 19073 27084
rect 19107 27081 19119 27115
rect 27154 27112 27160 27124
rect 19061 27075 19119 27081
rect 19720 27084 24716 27112
rect 27115 27084 27160 27112
rect 16914 27047 16972 27053
rect 16914 27044 16926 27047
rect 12952 27016 14044 27044
rect 12952 27004 12958 27016
rect 14016 26988 14044 27016
rect 14476 27016 16712 27044
rect 16776 27016 16926 27044
rect 12805 26979 12863 26985
rect 12805 26945 12817 26979
rect 12851 26945 12863 26979
rect 12805 26939 12863 26945
rect 12989 26979 13047 26985
rect 12989 26945 13001 26979
rect 13035 26945 13047 26979
rect 12989 26939 13047 26945
rect 13081 26979 13139 26985
rect 13081 26945 13093 26979
rect 13127 26976 13139 26979
rect 13725 26979 13783 26985
rect 13127 26948 13308 26976
rect 13127 26945 13139 26948
rect 13081 26939 13139 26945
rect 11480 26880 11744 26908
rect 13004 26908 13032 26939
rect 13170 26908 13176 26920
rect 13004 26880 13176 26908
rect 11480 26868 11486 26880
rect 13170 26868 13176 26880
rect 13228 26868 13234 26920
rect 13280 26852 13308 26948
rect 13725 26945 13737 26979
rect 13771 26945 13783 26979
rect 13725 26939 13783 26945
rect 13740 26908 13768 26939
rect 13814 26936 13820 26988
rect 13872 26976 13878 26988
rect 13909 26979 13967 26985
rect 13909 26976 13921 26979
rect 13872 26948 13921 26976
rect 13872 26936 13878 26948
rect 13909 26945 13921 26948
rect 13955 26945 13967 26979
rect 13909 26939 13967 26945
rect 13998 26936 14004 26988
rect 14056 26976 14062 26988
rect 14476 26985 14504 27016
rect 14734 26985 14740 26988
rect 14461 26979 14519 26985
rect 14056 26948 14101 26976
rect 14056 26936 14062 26948
rect 14461 26945 14473 26979
rect 14507 26945 14519 26979
rect 14461 26939 14519 26945
rect 14728 26939 14740 26985
rect 14792 26976 14798 26988
rect 16684 26985 16712 27016
rect 16914 27013 16926 27016
rect 16960 27013 16972 27047
rect 16914 27007 16972 27013
rect 18785 27047 18843 27053
rect 18785 27013 18797 27047
rect 18831 27044 18843 27047
rect 19334 27044 19340 27056
rect 18831 27016 19340 27044
rect 18831 27013 18843 27016
rect 18785 27007 18843 27013
rect 19334 27004 19340 27016
rect 19392 27004 19398 27056
rect 16669 26979 16727 26985
rect 14792 26948 14828 26976
rect 14734 26936 14740 26939
rect 14792 26936 14798 26948
rect 16669 26945 16681 26979
rect 16715 26976 16727 26979
rect 16758 26976 16764 26988
rect 16715 26948 16764 26976
rect 16715 26945 16727 26948
rect 16669 26939 16727 26945
rect 16758 26936 16764 26948
rect 16816 26936 16822 26988
rect 17678 26936 17684 26988
rect 17736 26976 17742 26988
rect 18509 26979 18567 26985
rect 18509 26976 18521 26979
rect 17736 26948 18521 26976
rect 17736 26936 17742 26948
rect 18509 26945 18521 26948
rect 18555 26945 18567 26979
rect 18690 26976 18696 26988
rect 18651 26948 18696 26976
rect 18509 26939 18567 26945
rect 18690 26936 18696 26948
rect 18748 26936 18754 26988
rect 18877 26979 18935 26985
rect 18877 26945 18889 26979
rect 18923 26945 18935 26979
rect 18877 26939 18935 26945
rect 13740 26880 14412 26908
rect 13262 26840 13268 26852
rect 7944 26812 8892 26840
rect 3804 26744 4844 26772
rect 2961 26735 3019 26741
rect 4890 26732 4896 26784
rect 4948 26772 4954 26784
rect 5074 26772 5080 26784
rect 4948 26744 5080 26772
rect 4948 26732 4954 26744
rect 5074 26732 5080 26744
rect 5132 26772 5138 26784
rect 5169 26775 5227 26781
rect 5169 26772 5181 26775
rect 5132 26744 5181 26772
rect 5132 26732 5138 26744
rect 5169 26741 5181 26744
rect 5215 26741 5227 26775
rect 5169 26735 5227 26741
rect 5350 26732 5356 26784
rect 5408 26772 5414 26784
rect 8662 26772 8668 26784
rect 5408 26744 8668 26772
rect 5408 26732 5414 26744
rect 8662 26732 8668 26744
rect 8720 26732 8726 26784
rect 8864 26772 8892 26812
rect 11992 26812 13268 26840
rect 9217 26775 9275 26781
rect 9217 26772 9229 26775
rect 8864 26744 9229 26772
rect 9217 26741 9229 26744
rect 9263 26741 9275 26775
rect 9217 26735 9275 26741
rect 9585 26775 9643 26781
rect 9585 26741 9597 26775
rect 9631 26772 9643 26775
rect 9674 26772 9680 26784
rect 9631 26744 9680 26772
rect 9631 26741 9643 26744
rect 9585 26735 9643 26741
rect 9674 26732 9680 26744
rect 9732 26732 9738 26784
rect 11146 26732 11152 26784
rect 11204 26772 11210 26784
rect 11992 26772 12020 26812
rect 13262 26800 13268 26812
rect 13320 26800 13326 26852
rect 13740 26840 13768 26880
rect 13648 26812 13768 26840
rect 11204 26744 12020 26772
rect 11204 26732 11210 26744
rect 12066 26732 12072 26784
rect 12124 26772 12130 26784
rect 13648 26772 13676 26812
rect 12124 26744 13676 26772
rect 13725 26775 13783 26781
rect 12124 26732 12130 26744
rect 13725 26741 13737 26775
rect 13771 26772 13783 26775
rect 14274 26772 14280 26784
rect 13771 26744 14280 26772
rect 13771 26741 13783 26744
rect 13725 26735 13783 26741
rect 14274 26732 14280 26744
rect 14332 26732 14338 26784
rect 14384 26772 14412 26880
rect 17954 26868 17960 26920
rect 18012 26908 18018 26920
rect 18892 26908 18920 26939
rect 19610 26908 19616 26920
rect 18012 26880 19616 26908
rect 18012 26868 18018 26880
rect 19610 26868 19616 26880
rect 19668 26868 19674 26920
rect 19720 26840 19748 27084
rect 20346 27004 20352 27056
rect 20404 27044 20410 27056
rect 21913 27047 21971 27053
rect 21913 27044 21925 27047
rect 20404 27016 21925 27044
rect 20404 27004 20410 27016
rect 21913 27013 21925 27016
rect 21959 27013 21971 27047
rect 24688 27044 24716 27084
rect 27154 27072 27160 27084
rect 27212 27072 27218 27124
rect 21913 27007 21971 27013
rect 22020 27016 24624 27044
rect 24688 27016 27384 27044
rect 22020 26988 22048 27016
rect 19886 26976 19892 26988
rect 19847 26948 19892 26976
rect 19886 26936 19892 26948
rect 19944 26936 19950 26988
rect 20156 26979 20214 26985
rect 20156 26945 20168 26979
rect 20202 26976 20214 26979
rect 20202 26948 21128 26976
rect 20202 26945 20214 26948
rect 20156 26939 20214 26945
rect 21100 26908 21128 26948
rect 21266 26936 21272 26988
rect 21324 26976 21330 26988
rect 21821 26979 21879 26985
rect 21821 26976 21833 26979
rect 21324 26948 21833 26976
rect 21324 26936 21330 26948
rect 21821 26945 21833 26948
rect 21867 26945 21879 26979
rect 21821 26939 21879 26945
rect 22002 26936 22008 26988
rect 22060 26976 22066 26988
rect 22646 26976 22652 26988
rect 22060 26948 22153 26976
rect 22607 26948 22652 26976
rect 22060 26936 22066 26948
rect 22646 26936 22652 26948
rect 22704 26936 22710 26988
rect 22830 26936 22836 26988
rect 22888 26976 22894 26988
rect 23293 26979 23351 26985
rect 23293 26976 23305 26979
rect 22888 26948 23305 26976
rect 22888 26936 22894 26948
rect 23293 26945 23305 26948
rect 23339 26945 23351 26979
rect 23293 26939 23351 26945
rect 23842 26936 23848 26988
rect 23900 26976 23906 26988
rect 23937 26979 23995 26985
rect 23937 26976 23949 26979
rect 23900 26948 23949 26976
rect 23900 26936 23906 26948
rect 23937 26945 23949 26948
rect 23983 26945 23995 26979
rect 23937 26939 23995 26945
rect 24210 26936 24216 26988
rect 24268 26976 24274 26988
rect 24596 26985 24624 27016
rect 24397 26979 24455 26985
rect 24397 26976 24409 26979
rect 24268 26948 24409 26976
rect 24268 26936 24274 26948
rect 24397 26945 24409 26948
rect 24443 26945 24455 26979
rect 24397 26939 24455 26945
rect 24581 26979 24639 26985
rect 24581 26945 24593 26979
rect 24627 26945 24639 26979
rect 24581 26939 24639 26945
rect 25777 26979 25835 26985
rect 25777 26945 25789 26979
rect 25823 26976 25835 26979
rect 25958 26976 25964 26988
rect 25823 26948 25964 26976
rect 25823 26945 25835 26948
rect 25777 26939 25835 26945
rect 25958 26936 25964 26948
rect 26016 26936 26022 26988
rect 26418 26976 26424 26988
rect 26379 26948 26424 26976
rect 26418 26936 26424 26948
rect 26476 26936 26482 26988
rect 27356 26985 27384 27016
rect 27341 26979 27399 26985
rect 27341 26945 27353 26979
rect 27387 26945 27399 26979
rect 27341 26939 27399 26945
rect 21100 26880 22508 26908
rect 17604 26812 19748 26840
rect 15378 26772 15384 26784
rect 14384 26744 15384 26772
rect 15378 26732 15384 26744
rect 15436 26732 15442 26784
rect 15838 26772 15844 26784
rect 15799 26744 15844 26772
rect 15838 26732 15844 26744
rect 15896 26732 15902 26784
rect 15930 26732 15936 26784
rect 15988 26772 15994 26784
rect 17604 26772 17632 26812
rect 21450 26800 21456 26852
rect 21508 26840 21514 26852
rect 22278 26840 22284 26852
rect 21508 26812 22284 26840
rect 21508 26800 21514 26812
rect 22278 26800 22284 26812
rect 22336 26800 22342 26852
rect 22480 26849 22508 26880
rect 22465 26843 22523 26849
rect 22465 26809 22477 26843
rect 22511 26809 22523 26843
rect 24397 26843 24455 26849
rect 24397 26840 24409 26843
rect 22465 26803 22523 26809
rect 23032 26812 24409 26840
rect 15988 26744 17632 26772
rect 18049 26775 18107 26781
rect 15988 26732 15994 26744
rect 18049 26741 18061 26775
rect 18095 26772 18107 26775
rect 18138 26772 18144 26784
rect 18095 26744 18144 26772
rect 18095 26741 18107 26744
rect 18049 26735 18107 26741
rect 18138 26732 18144 26744
rect 18196 26732 18202 26784
rect 20806 26732 20812 26784
rect 20864 26772 20870 26784
rect 21269 26775 21327 26781
rect 21269 26772 21281 26775
rect 20864 26744 21281 26772
rect 20864 26732 20870 26744
rect 21269 26741 21281 26744
rect 21315 26741 21327 26775
rect 21269 26735 21327 26741
rect 21634 26732 21640 26784
rect 21692 26772 21698 26784
rect 23032 26772 23060 26812
rect 24397 26809 24409 26812
rect 24443 26809 24455 26843
rect 24397 26803 24455 26809
rect 21692 26744 23060 26772
rect 21692 26732 21698 26744
rect 23106 26732 23112 26784
rect 23164 26772 23170 26784
rect 23753 26775 23811 26781
rect 23164 26744 23209 26772
rect 23164 26732 23170 26744
rect 23753 26741 23765 26775
rect 23799 26772 23811 26775
rect 24210 26772 24216 26784
rect 23799 26744 24216 26772
rect 23799 26741 23811 26744
rect 23753 26735 23811 26741
rect 24210 26732 24216 26744
rect 24268 26732 24274 26784
rect 25593 26775 25651 26781
rect 25593 26741 25605 26775
rect 25639 26772 25651 26775
rect 25682 26772 25688 26784
rect 25639 26744 25688 26772
rect 25639 26741 25651 26744
rect 25593 26735 25651 26741
rect 25682 26732 25688 26744
rect 25740 26732 25746 26784
rect 26234 26772 26240 26784
rect 26195 26744 26240 26772
rect 26234 26732 26240 26744
rect 26292 26732 26298 26784
rect 1104 26682 28060 26704
rect 1104 26630 5442 26682
rect 5494 26630 5506 26682
rect 5558 26630 5570 26682
rect 5622 26630 5634 26682
rect 5686 26630 5698 26682
rect 5750 26630 14428 26682
rect 14480 26630 14492 26682
rect 14544 26630 14556 26682
rect 14608 26630 14620 26682
rect 14672 26630 14684 26682
rect 14736 26630 23413 26682
rect 23465 26630 23477 26682
rect 23529 26630 23541 26682
rect 23593 26630 23605 26682
rect 23657 26630 23669 26682
rect 23721 26630 28060 26682
rect 1104 26608 28060 26630
rect 4522 26568 4528 26580
rect 4483 26540 4528 26568
rect 4522 26528 4528 26540
rect 4580 26528 4586 26580
rect 5537 26571 5595 26577
rect 5537 26537 5549 26571
rect 5583 26568 5595 26571
rect 5810 26568 5816 26580
rect 5583 26540 5816 26568
rect 5583 26537 5595 26540
rect 5537 26531 5595 26537
rect 5810 26528 5816 26540
rect 5868 26528 5874 26580
rect 7466 26528 7472 26580
rect 7524 26568 7530 26580
rect 8202 26568 8208 26580
rect 7524 26540 8208 26568
rect 7524 26528 7530 26540
rect 8202 26528 8208 26540
rect 8260 26528 8266 26580
rect 8294 26528 8300 26580
rect 8352 26568 8358 26580
rect 9033 26571 9091 26577
rect 9033 26568 9045 26571
rect 8352 26540 9045 26568
rect 8352 26528 8358 26540
rect 9033 26537 9045 26540
rect 9079 26537 9091 26571
rect 9033 26531 9091 26537
rect 9858 26528 9864 26580
rect 9916 26568 9922 26580
rect 9953 26571 10011 26577
rect 9953 26568 9965 26571
rect 9916 26540 9965 26568
rect 9916 26528 9922 26540
rect 9953 26537 9965 26540
rect 9999 26537 10011 26571
rect 9953 26531 10011 26537
rect 10042 26528 10048 26580
rect 10100 26568 10106 26580
rect 11422 26568 11428 26580
rect 10100 26540 11428 26568
rect 10100 26528 10106 26540
rect 11422 26528 11428 26540
rect 11480 26528 11486 26580
rect 14274 26528 14280 26580
rect 14332 26568 14338 26580
rect 14461 26571 14519 26577
rect 14461 26568 14473 26571
rect 14332 26540 14473 26568
rect 14332 26528 14338 26540
rect 14461 26537 14473 26540
rect 14507 26537 14519 26571
rect 14461 26531 14519 26537
rect 14553 26571 14611 26577
rect 14553 26537 14565 26571
rect 14599 26568 14611 26571
rect 14826 26568 14832 26580
rect 14599 26540 14832 26568
rect 14599 26537 14611 26540
rect 14553 26531 14611 26537
rect 14826 26528 14832 26540
rect 14884 26528 14890 26580
rect 16022 26528 16028 26580
rect 16080 26568 16086 26580
rect 16669 26571 16727 26577
rect 16669 26568 16681 26571
rect 16080 26540 16681 26568
rect 16080 26528 16086 26540
rect 16669 26537 16681 26540
rect 16715 26537 16727 26571
rect 19794 26568 19800 26580
rect 19755 26540 19800 26568
rect 16669 26531 16727 26537
rect 19794 26528 19800 26540
rect 19852 26528 19858 26580
rect 21450 26568 21456 26580
rect 21411 26540 21456 26568
rect 21450 26528 21456 26540
rect 21508 26528 21514 26580
rect 22646 26568 22652 26580
rect 21560 26540 22652 26568
rect 1578 26460 1584 26512
rect 1636 26500 1642 26512
rect 1857 26503 1915 26509
rect 1857 26500 1869 26503
rect 1636 26472 1869 26500
rect 1636 26460 1642 26472
rect 1857 26469 1869 26472
rect 1903 26469 1915 26503
rect 3418 26500 3424 26512
rect 1857 26463 1915 26469
rect 3068 26472 3424 26500
rect 3068 26373 3096 26472
rect 3418 26460 3424 26472
rect 3476 26500 3482 26512
rect 3476 26472 5120 26500
rect 3476 26460 3482 26472
rect 3145 26435 3203 26441
rect 3145 26401 3157 26435
rect 3191 26432 3203 26435
rect 4065 26435 4123 26441
rect 3191 26404 4016 26432
rect 3191 26401 3203 26404
rect 3145 26395 3203 26401
rect 2041 26367 2099 26373
rect 2041 26333 2053 26367
rect 2087 26364 2099 26367
rect 3053 26367 3111 26373
rect 2087 26336 2452 26364
rect 2087 26333 2099 26336
rect 2041 26327 2099 26333
rect 2424 26305 2452 26336
rect 3053 26333 3065 26367
rect 3099 26333 3111 26367
rect 3053 26327 3111 26333
rect 3237 26367 3295 26373
rect 3237 26333 3249 26367
rect 3283 26364 3295 26367
rect 3510 26364 3516 26376
rect 3283 26336 3516 26364
rect 3283 26333 3295 26336
rect 3237 26327 3295 26333
rect 3510 26324 3516 26336
rect 3568 26324 3574 26376
rect 3988 26373 4016 26404
rect 4065 26401 4077 26435
rect 4111 26432 4123 26435
rect 4617 26435 4675 26441
rect 4617 26432 4629 26435
rect 4111 26404 4629 26432
rect 4111 26401 4123 26404
rect 4065 26395 4123 26401
rect 4617 26401 4629 26404
rect 4663 26401 4675 26435
rect 4890 26432 4896 26444
rect 4617 26395 4675 26401
rect 4724 26404 4896 26432
rect 3789 26367 3847 26373
rect 3789 26333 3801 26367
rect 3835 26333 3847 26367
rect 3789 26327 3847 26333
rect 3973 26367 4031 26373
rect 3973 26333 3985 26367
rect 4019 26333 4031 26367
rect 4154 26364 4160 26376
rect 4115 26336 4160 26364
rect 3973 26327 4031 26333
rect 2409 26299 2467 26305
rect 2409 26265 2421 26299
rect 2455 26296 2467 26299
rect 2682 26296 2688 26308
rect 2455 26268 2688 26296
rect 2455 26265 2467 26268
rect 2409 26259 2467 26265
rect 2682 26256 2688 26268
rect 2740 26256 2746 26308
rect 3804 26296 3832 26327
rect 4154 26324 4160 26336
rect 4212 26324 4218 26376
rect 4341 26367 4399 26373
rect 4341 26333 4353 26367
rect 4387 26364 4399 26367
rect 4724 26364 4752 26404
rect 4890 26392 4896 26404
rect 4948 26392 4954 26444
rect 4387 26336 4752 26364
rect 4387 26333 4399 26336
rect 4341 26327 4399 26333
rect 4798 26324 4804 26376
rect 4856 26364 4862 26376
rect 5092 26373 5120 26472
rect 5166 26460 5172 26512
rect 5224 26500 5230 26512
rect 7745 26503 7803 26509
rect 5224 26472 7696 26500
rect 5224 26460 5230 26472
rect 5350 26432 5356 26444
rect 5184 26404 5356 26432
rect 5077 26367 5135 26373
rect 4856 26336 4901 26364
rect 4856 26324 4862 26336
rect 5077 26333 5089 26367
rect 5123 26333 5135 26367
rect 5077 26327 5135 26333
rect 4062 26296 4068 26308
rect 3804 26268 4068 26296
rect 4062 26256 4068 26268
rect 4120 26296 4126 26308
rect 5184 26296 5212 26404
rect 5350 26392 5356 26404
rect 5408 26392 5414 26444
rect 5442 26392 5448 26444
rect 5500 26432 5506 26444
rect 5500 26404 7604 26432
rect 5500 26392 5506 26404
rect 5258 26324 5264 26376
rect 5316 26364 5322 26376
rect 5316 26336 5361 26364
rect 5537 26345 5595 26351
rect 5316 26324 5322 26336
rect 5537 26311 5549 26345
rect 5583 26340 5595 26345
rect 5626 26340 5632 26376
rect 5583 26324 5632 26340
rect 5684 26364 5690 26376
rect 5997 26367 6055 26373
rect 5684 26336 5777 26364
rect 5684 26324 5690 26336
rect 5583 26312 5678 26324
rect 5583 26311 5595 26312
rect 5537 26305 5595 26311
rect 5445 26299 5503 26305
rect 5445 26296 5457 26299
rect 4120 26268 5212 26296
rect 4120 26256 4126 26268
rect 5440 26265 5457 26296
rect 5491 26265 5503 26299
rect 5727 26296 5755 26336
rect 5997 26333 6009 26367
rect 6043 26364 6055 26367
rect 6086 26364 6092 26376
rect 6043 26336 6092 26364
rect 6043 26333 6055 26336
rect 5997 26327 6055 26333
rect 6086 26324 6092 26336
rect 6144 26324 6150 26376
rect 6178 26324 6184 26376
rect 6236 26364 6242 26376
rect 7377 26367 7435 26373
rect 6236 26336 6281 26364
rect 6236 26324 6242 26336
rect 7377 26333 7389 26367
rect 7423 26364 7435 26367
rect 7466 26364 7472 26376
rect 7423 26336 7472 26364
rect 7423 26333 7435 26336
rect 7377 26327 7435 26333
rect 7466 26324 7472 26336
rect 7524 26324 7530 26376
rect 7576 26373 7604 26404
rect 7668 26373 7696 26472
rect 7745 26469 7757 26503
rect 7791 26500 7803 26503
rect 8386 26500 8392 26512
rect 7791 26472 8392 26500
rect 7791 26469 7803 26472
rect 7745 26463 7803 26469
rect 8386 26460 8392 26472
rect 8444 26460 8450 26512
rect 10318 26500 10324 26512
rect 9140 26472 10324 26500
rect 7837 26435 7895 26441
rect 7837 26401 7849 26435
rect 7883 26432 7895 26435
rect 8018 26432 8024 26444
rect 7883 26404 8024 26432
rect 7883 26401 7895 26404
rect 7837 26395 7895 26401
rect 8018 26392 8024 26404
rect 8076 26392 8082 26444
rect 7561 26367 7619 26373
rect 7561 26333 7573 26367
rect 7607 26333 7619 26367
rect 7561 26327 7619 26333
rect 7653 26367 7711 26373
rect 7653 26333 7665 26367
rect 7699 26333 7711 26367
rect 7653 26327 7711 26333
rect 7929 26367 7987 26373
rect 7929 26333 7941 26367
rect 7975 26364 7987 26367
rect 9140 26364 9168 26472
rect 10318 26460 10324 26472
rect 10376 26460 10382 26512
rect 13998 26460 14004 26512
rect 14056 26500 14062 26512
rect 15841 26503 15899 26509
rect 14056 26472 14228 26500
rect 14056 26460 14062 26472
rect 10042 26432 10048 26444
rect 9232 26404 10048 26432
rect 9232 26373 9260 26404
rect 10042 26392 10048 26404
rect 10100 26392 10106 26444
rect 11057 26435 11115 26441
rect 11057 26432 11069 26435
rect 10152 26404 11069 26432
rect 10152 26373 10180 26404
rect 11057 26401 11069 26404
rect 11103 26401 11115 26435
rect 11057 26395 11115 26401
rect 11425 26435 11483 26441
rect 11425 26401 11437 26435
rect 11471 26432 11483 26435
rect 12526 26432 12532 26444
rect 11471 26404 12532 26432
rect 11471 26401 11483 26404
rect 11425 26395 11483 26401
rect 12526 26392 12532 26404
rect 12584 26392 12590 26444
rect 12894 26392 12900 26444
rect 12952 26432 12958 26444
rect 12952 26404 12997 26432
rect 12952 26392 12958 26404
rect 7975 26336 9168 26364
rect 9217 26367 9275 26373
rect 7975 26333 7987 26336
rect 7929 26327 7987 26333
rect 9217 26333 9229 26367
rect 9263 26333 9275 26367
rect 9493 26367 9551 26373
rect 9493 26364 9505 26367
rect 9217 26327 9275 26333
rect 9324 26336 9505 26364
rect 6733 26299 6791 26305
rect 5727 26268 6592 26296
rect 5440 26259 5503 26265
rect 2958 26188 2964 26240
rect 3016 26228 3022 26240
rect 4890 26228 4896 26240
rect 3016 26200 4896 26228
rect 3016 26188 3022 26200
rect 4890 26188 4896 26200
rect 4948 26188 4954 26240
rect 4985 26231 5043 26237
rect 4985 26197 4997 26231
rect 5031 26228 5043 26231
rect 5440 26228 5468 26259
rect 5902 26228 5908 26240
rect 5031 26200 5908 26228
rect 5031 26197 5043 26200
rect 4985 26191 5043 26197
rect 5902 26188 5908 26200
rect 5960 26188 5966 26240
rect 6089 26231 6147 26237
rect 6089 26197 6101 26231
rect 6135 26228 6147 26231
rect 6454 26228 6460 26240
rect 6135 26200 6460 26228
rect 6135 26197 6147 26200
rect 6089 26191 6147 26197
rect 6454 26188 6460 26200
rect 6512 26188 6518 26240
rect 6564 26228 6592 26268
rect 6733 26265 6745 26299
rect 6779 26296 6791 26299
rect 8662 26296 8668 26308
rect 6779 26268 8668 26296
rect 6779 26265 6791 26268
rect 6733 26259 6791 26265
rect 8662 26256 8668 26268
rect 8720 26256 8726 26308
rect 9324 26296 9352 26336
rect 9493 26333 9505 26336
rect 9539 26364 9551 26367
rect 10137 26367 10195 26373
rect 9539 26336 9996 26364
rect 9539 26333 9551 26336
rect 9493 26327 9551 26333
rect 8772 26268 9352 26296
rect 9968 26296 9996 26336
rect 10137 26333 10149 26367
rect 10183 26333 10195 26367
rect 10410 26364 10416 26376
rect 10323 26336 10416 26364
rect 10137 26327 10195 26333
rect 10410 26324 10416 26336
rect 10468 26364 10474 26376
rect 10468 26336 10548 26364
rect 10468 26324 10474 26336
rect 9968 26268 10456 26296
rect 6825 26231 6883 26237
rect 6825 26228 6837 26231
rect 6564 26200 6837 26228
rect 6825 26197 6837 26200
rect 6871 26228 6883 26231
rect 7190 26228 7196 26240
rect 6871 26200 7196 26228
rect 6871 26197 6883 26200
rect 6825 26191 6883 26197
rect 7190 26188 7196 26200
rect 7248 26188 7254 26240
rect 7466 26188 7472 26240
rect 7524 26228 7530 26240
rect 8772 26228 8800 26268
rect 10428 26240 10456 26268
rect 7524 26200 8800 26228
rect 9401 26231 9459 26237
rect 7524 26188 7530 26200
rect 9401 26197 9413 26231
rect 9447 26228 9459 26231
rect 9766 26228 9772 26240
rect 9447 26200 9772 26228
rect 9447 26197 9459 26200
rect 9401 26191 9459 26197
rect 9766 26188 9772 26200
rect 9824 26188 9830 26240
rect 10410 26188 10416 26240
rect 10468 26188 10474 26240
rect 10520 26228 10548 26336
rect 10594 26324 10600 26376
rect 10652 26364 10658 26376
rect 10652 26336 10697 26364
rect 10652 26324 10658 26336
rect 10870 26324 10876 26376
rect 10928 26364 10934 26376
rect 11241 26367 11299 26373
rect 11241 26364 11253 26367
rect 10928 26336 11253 26364
rect 10928 26324 10934 26336
rect 11241 26333 11253 26336
rect 11287 26333 11299 26367
rect 11241 26327 11299 26333
rect 11333 26367 11391 26373
rect 11333 26333 11345 26367
rect 11379 26333 11391 26367
rect 11517 26367 11575 26373
rect 11333 26327 11391 26333
rect 10612 26296 10640 26324
rect 11348 26296 11376 26327
rect 11422 26314 11428 26366
rect 11480 26364 11486 26366
rect 11517 26364 11529 26367
rect 11480 26336 11529 26364
rect 11480 26314 11486 26336
rect 11517 26333 11529 26336
rect 11563 26333 11575 26367
rect 11517 26327 11575 26333
rect 12250 26324 12256 26376
rect 12308 26364 12314 26376
rect 12621 26367 12679 26373
rect 12621 26364 12633 26367
rect 12308 26336 12633 26364
rect 12308 26324 12314 26336
rect 12621 26333 12633 26336
rect 12667 26333 12679 26367
rect 14090 26364 14096 26376
rect 14051 26336 14096 26364
rect 12621 26327 12679 26333
rect 14090 26324 14096 26336
rect 14148 26324 14154 26376
rect 14200 26373 14228 26472
rect 15841 26469 15853 26503
rect 15887 26500 15899 26503
rect 16482 26500 16488 26512
rect 15887 26472 16488 26500
rect 15887 26469 15899 26472
rect 15841 26463 15899 26469
rect 16482 26460 16488 26472
rect 16540 26460 16546 26512
rect 18141 26503 18199 26509
rect 18141 26469 18153 26503
rect 18187 26469 18199 26503
rect 20625 26503 20683 26509
rect 18141 26463 18199 26469
rect 19306 26472 20300 26500
rect 18156 26432 18184 26463
rect 15672 26404 18184 26432
rect 14185 26367 14243 26373
rect 14185 26333 14197 26367
rect 14231 26333 14243 26367
rect 14550 26364 14556 26376
rect 14511 26336 14556 26364
rect 14185 26327 14243 26333
rect 14550 26324 14556 26336
rect 14608 26324 14614 26376
rect 15672 26373 15700 26404
rect 18782 26392 18788 26444
rect 18840 26432 18846 26444
rect 19306 26432 19334 26472
rect 20272 26441 20300 26472
rect 20625 26469 20637 26503
rect 20671 26500 20683 26503
rect 21560 26500 21588 26540
rect 22646 26528 22652 26540
rect 22704 26528 22710 26580
rect 26237 26571 26295 26577
rect 26237 26537 26249 26571
rect 26283 26568 26295 26571
rect 27706 26568 27712 26580
rect 26283 26540 27712 26568
rect 26283 26537 26295 26540
rect 26237 26531 26295 26537
rect 27706 26528 27712 26540
rect 27764 26528 27770 26580
rect 20671 26472 21588 26500
rect 20671 26469 20683 26472
rect 20625 26463 20683 26469
rect 26510 26460 26516 26512
rect 26568 26500 26574 26512
rect 26881 26503 26939 26509
rect 26881 26500 26893 26503
rect 26568 26472 26893 26500
rect 26568 26460 26574 26472
rect 26881 26469 26893 26472
rect 26927 26469 26939 26503
rect 26881 26463 26939 26469
rect 18840 26404 19334 26432
rect 20257 26435 20315 26441
rect 18840 26392 18846 26404
rect 20257 26401 20269 26435
rect 20303 26432 20315 26435
rect 20530 26432 20536 26444
rect 20303 26404 20536 26432
rect 20303 26401 20315 26404
rect 20257 26395 20315 26401
rect 20530 26392 20536 26404
rect 20588 26432 20594 26444
rect 20588 26404 21220 26432
rect 20588 26392 20594 26404
rect 21192 26376 21220 26404
rect 21818 26392 21824 26444
rect 21876 26432 21882 26444
rect 21913 26435 21971 26441
rect 21913 26432 21925 26435
rect 21876 26404 21925 26432
rect 21876 26392 21882 26404
rect 21913 26401 21925 26404
rect 21959 26401 21971 26435
rect 21913 26395 21971 26401
rect 15473 26367 15531 26373
rect 15473 26333 15485 26367
rect 15519 26333 15531 26367
rect 15473 26327 15531 26333
rect 15657 26367 15715 26373
rect 15657 26333 15669 26367
rect 15703 26333 15715 26367
rect 15657 26327 15715 26333
rect 16301 26367 16359 26373
rect 16301 26333 16313 26367
rect 16347 26333 16359 26367
rect 16301 26327 16359 26333
rect 16485 26367 16543 26373
rect 16485 26333 16497 26367
rect 16531 26364 16543 26367
rect 17494 26364 17500 26376
rect 16531 26336 17500 26364
rect 16531 26333 16543 26336
rect 16485 26327 16543 26333
rect 10612 26268 11376 26296
rect 13354 26256 13360 26308
rect 13412 26296 13418 26308
rect 15488 26296 15516 26327
rect 16316 26296 16344 26327
rect 17494 26324 17500 26336
rect 17552 26324 17558 26376
rect 17589 26367 17647 26373
rect 17589 26333 17601 26367
rect 17635 26364 17647 26367
rect 17678 26364 17684 26376
rect 17635 26336 17684 26364
rect 17635 26333 17647 26336
rect 17589 26327 17647 26333
rect 17678 26324 17684 26336
rect 17736 26324 17742 26376
rect 17954 26364 17960 26376
rect 17915 26336 17960 26364
rect 17954 26324 17960 26336
rect 18012 26324 18018 26376
rect 19245 26367 19303 26373
rect 19245 26333 19257 26367
rect 19291 26333 19303 26367
rect 19426 26364 19432 26376
rect 19387 26336 19432 26364
rect 19245 26327 19303 26333
rect 17770 26296 17776 26308
rect 13412 26268 16344 26296
rect 17731 26268 17776 26296
rect 13412 26256 13418 26268
rect 17770 26256 17776 26268
rect 17828 26256 17834 26308
rect 17865 26299 17923 26305
rect 17865 26265 17877 26299
rect 17911 26296 17923 26299
rect 18046 26296 18052 26308
rect 17911 26268 18052 26296
rect 17911 26265 17923 26268
rect 17865 26259 17923 26265
rect 18046 26256 18052 26268
rect 18104 26296 18110 26308
rect 18414 26296 18420 26308
rect 18104 26268 18420 26296
rect 18104 26256 18110 26268
rect 18414 26256 18420 26268
rect 18472 26256 18478 26308
rect 19260 26240 19288 26327
rect 19426 26324 19432 26336
rect 19484 26324 19490 26376
rect 19610 26364 19616 26376
rect 19571 26336 19616 26364
rect 19610 26324 19616 26336
rect 19668 26364 19674 26376
rect 19794 26364 19800 26376
rect 19668 26336 19800 26364
rect 19668 26324 19674 26336
rect 19794 26324 19800 26336
rect 19852 26324 19858 26376
rect 20438 26364 20444 26376
rect 20399 26336 20444 26364
rect 20438 26324 20444 26336
rect 20496 26324 20502 26376
rect 21174 26364 21180 26376
rect 21135 26336 21180 26364
rect 21174 26324 21180 26336
rect 21232 26324 21238 26376
rect 21269 26367 21327 26373
rect 21269 26333 21281 26367
rect 21315 26333 21327 26367
rect 21928 26364 21956 26395
rect 24397 26367 24455 26373
rect 24397 26364 24409 26367
rect 21928 26336 24409 26364
rect 21269 26327 21327 26333
rect 24397 26333 24409 26336
rect 24443 26364 24455 26367
rect 25406 26364 25412 26376
rect 24443 26336 25412 26364
rect 24443 26333 24455 26336
rect 24397 26327 24455 26333
rect 19521 26299 19579 26305
rect 19521 26265 19533 26299
rect 19567 26296 19579 26299
rect 20070 26296 20076 26308
rect 19567 26268 20076 26296
rect 19567 26265 19579 26268
rect 19521 26259 19579 26265
rect 20070 26256 20076 26268
rect 20128 26256 20134 26308
rect 21284 26296 21312 26327
rect 25406 26324 25412 26336
rect 25464 26324 25470 26376
rect 26421 26367 26479 26373
rect 26421 26333 26433 26367
rect 26467 26364 26479 26367
rect 26694 26364 26700 26376
rect 26467 26336 26700 26364
rect 26467 26333 26479 26336
rect 26421 26327 26479 26333
rect 26694 26324 26700 26336
rect 26752 26324 26758 26376
rect 27065 26367 27123 26373
rect 27065 26333 27077 26367
rect 27111 26333 27123 26367
rect 27065 26327 27123 26333
rect 22180 26299 22238 26305
rect 21284 26268 22140 26296
rect 10778 26228 10784 26240
rect 10520 26200 10784 26228
rect 10778 26188 10784 26200
rect 10836 26188 10842 26240
rect 11422 26188 11428 26240
rect 11480 26228 11486 26240
rect 13998 26228 14004 26240
rect 11480 26200 14004 26228
rect 11480 26188 11486 26200
rect 13998 26188 14004 26200
rect 14056 26188 14062 26240
rect 14277 26231 14335 26237
rect 14277 26197 14289 26231
rect 14323 26228 14335 26231
rect 15378 26228 15384 26240
rect 14323 26200 15384 26228
rect 14323 26197 14335 26200
rect 14277 26191 14335 26197
rect 15378 26188 15384 26200
rect 15436 26228 15442 26240
rect 15930 26228 15936 26240
rect 15436 26200 15936 26228
rect 15436 26188 15442 26200
rect 15930 26188 15936 26200
rect 15988 26188 15994 26240
rect 17678 26188 17684 26240
rect 17736 26228 17742 26240
rect 19242 26228 19248 26240
rect 17736 26200 19248 26228
rect 17736 26188 17742 26200
rect 19242 26188 19248 26200
rect 19300 26188 19306 26240
rect 22112 26228 22140 26268
rect 22180 26265 22192 26299
rect 22226 26296 22238 26299
rect 22370 26296 22376 26308
rect 22226 26268 22376 26296
rect 22226 26265 22238 26268
rect 22180 26259 22238 26265
rect 22370 26256 22376 26268
rect 22428 26256 22434 26308
rect 24486 26256 24492 26308
rect 24544 26296 24550 26308
rect 24642 26299 24700 26305
rect 24642 26296 24654 26299
rect 24544 26268 24654 26296
rect 24544 26256 24550 26268
rect 24642 26265 24654 26268
rect 24688 26265 24700 26299
rect 24642 26259 24700 26265
rect 25498 26256 25504 26308
rect 25556 26296 25562 26308
rect 27080 26296 27108 26327
rect 25556 26268 27108 26296
rect 25556 26256 25562 26268
rect 22278 26228 22284 26240
rect 22112 26200 22284 26228
rect 22278 26188 22284 26200
rect 22336 26188 22342 26240
rect 22738 26188 22744 26240
rect 22796 26228 22802 26240
rect 23293 26231 23351 26237
rect 23293 26228 23305 26231
rect 22796 26200 23305 26228
rect 22796 26188 22802 26200
rect 23293 26197 23305 26200
rect 23339 26197 23351 26231
rect 23293 26191 23351 26197
rect 24026 26188 24032 26240
rect 24084 26228 24090 26240
rect 25777 26231 25835 26237
rect 25777 26228 25789 26231
rect 24084 26200 25789 26228
rect 24084 26188 24090 26200
rect 25777 26197 25789 26200
rect 25823 26197 25835 26231
rect 25777 26191 25835 26197
rect 1104 26138 28060 26160
rect 1104 26086 9935 26138
rect 9987 26086 9999 26138
rect 10051 26086 10063 26138
rect 10115 26086 10127 26138
rect 10179 26086 10191 26138
rect 10243 26086 18920 26138
rect 18972 26086 18984 26138
rect 19036 26086 19048 26138
rect 19100 26086 19112 26138
rect 19164 26086 19176 26138
rect 19228 26086 28060 26138
rect 1104 26064 28060 26086
rect 4798 25984 4804 26036
rect 4856 26024 4862 26036
rect 4856 25996 5764 26024
rect 4856 25984 4862 25996
rect 2124 25959 2182 25965
rect 2124 25925 2136 25959
rect 2170 25956 2182 25959
rect 4709 25959 4767 25965
rect 4709 25956 4721 25959
rect 2170 25928 4721 25956
rect 2170 25925 2182 25928
rect 2124 25919 2182 25925
rect 4709 25925 4721 25928
rect 4755 25925 4767 25959
rect 4709 25919 4767 25925
rect 3973 25891 4031 25897
rect 3973 25857 3985 25891
rect 4019 25888 4031 25891
rect 4062 25888 4068 25900
rect 4019 25860 4068 25888
rect 4019 25857 4031 25860
rect 3973 25851 4031 25857
rect 4062 25848 4068 25860
rect 4120 25848 4126 25900
rect 4154 25848 4160 25900
rect 4212 25888 4218 25900
rect 4212 25860 4257 25888
rect 4212 25848 4218 25860
rect 4522 25848 4528 25900
rect 4580 25888 4586 25900
rect 5184 25888 5212 25996
rect 5258 25916 5264 25968
rect 5316 25956 5322 25968
rect 5736 25956 5764 25996
rect 7190 25984 7196 26036
rect 7248 26024 7254 26036
rect 7834 26024 7840 26036
rect 7248 25996 7840 26024
rect 7248 25984 7254 25996
rect 7834 25984 7840 25996
rect 7892 25984 7898 26036
rect 8662 26024 8668 26036
rect 8623 25996 8668 26024
rect 8662 25984 8668 25996
rect 8720 26024 8726 26036
rect 10870 26024 10876 26036
rect 8720 25996 10876 26024
rect 8720 25984 8726 25996
rect 7466 25956 7472 25968
rect 5316 25928 5678 25956
rect 5736 25928 7472 25956
rect 5316 25916 5322 25928
rect 5353 25891 5411 25897
rect 5353 25888 5365 25891
rect 4580 25860 4625 25888
rect 5184 25860 5365 25888
rect 4580 25848 4586 25860
rect 5353 25857 5365 25860
rect 5399 25857 5411 25891
rect 5353 25851 5411 25857
rect 5442 25848 5448 25900
rect 5500 25888 5506 25900
rect 5650 25897 5678 25928
rect 7466 25916 7472 25928
rect 7524 25916 7530 25968
rect 10520 25965 10548 25996
rect 10870 25984 10876 25996
rect 10928 25984 10934 26036
rect 11514 25984 11520 26036
rect 11572 26024 11578 26036
rect 11977 26027 12035 26033
rect 11977 26024 11989 26027
rect 11572 25996 11989 26024
rect 11572 25984 11578 25996
rect 11977 25993 11989 25996
rect 12023 25993 12035 26027
rect 11977 25987 12035 25993
rect 12434 25984 12440 26036
rect 12492 26024 12498 26036
rect 12492 25996 12572 26024
rect 12492 25984 12498 25996
rect 8113 25959 8171 25965
rect 8113 25925 8125 25959
rect 8159 25956 8171 25959
rect 9033 25959 9091 25965
rect 9033 25956 9045 25959
rect 8159 25928 9045 25956
rect 8159 25925 8171 25928
rect 8113 25919 8171 25925
rect 9033 25925 9045 25928
rect 9079 25956 9091 25959
rect 10505 25959 10563 25965
rect 9079 25928 10088 25956
rect 9079 25925 9091 25928
rect 9033 25919 9091 25925
rect 5537 25891 5595 25897
rect 5537 25888 5549 25891
rect 5500 25860 5549 25888
rect 5500 25848 5506 25860
rect 5537 25857 5549 25860
rect 5583 25857 5595 25891
rect 5537 25851 5595 25857
rect 5629 25891 5687 25897
rect 5629 25857 5641 25891
rect 5675 25857 5687 25891
rect 5629 25851 5687 25857
rect 6365 25891 6423 25897
rect 6365 25857 6377 25891
rect 6411 25857 6423 25891
rect 6365 25851 6423 25857
rect 1394 25780 1400 25832
rect 1452 25820 1458 25832
rect 1854 25820 1860 25832
rect 1452 25792 1860 25820
rect 1452 25780 1458 25792
rect 1854 25780 1860 25792
rect 1912 25780 1918 25832
rect 4249 25823 4307 25829
rect 4249 25789 4261 25823
rect 4295 25789 4307 25823
rect 4249 25783 4307 25789
rect 4341 25823 4399 25829
rect 4341 25789 4353 25823
rect 4387 25820 4399 25823
rect 4430 25820 4436 25832
rect 4387 25792 4436 25820
rect 4387 25789 4399 25792
rect 4341 25783 4399 25789
rect 4264 25752 4292 25783
rect 4430 25780 4436 25792
rect 4488 25780 4494 25832
rect 4614 25780 4620 25832
rect 4672 25820 4678 25832
rect 6380 25820 6408 25851
rect 7558 25848 7564 25900
rect 7616 25888 7622 25900
rect 7929 25891 7987 25897
rect 7929 25888 7941 25891
rect 7616 25860 7941 25888
rect 7616 25848 7622 25860
rect 7929 25857 7941 25860
rect 7975 25857 7987 25891
rect 7929 25851 7987 25857
rect 8205 25891 8263 25897
rect 8205 25857 8217 25891
rect 8251 25857 8263 25891
rect 8846 25888 8852 25900
rect 8807 25860 8852 25888
rect 8205 25851 8263 25857
rect 4672 25792 6408 25820
rect 6641 25823 6699 25829
rect 4672 25780 4678 25792
rect 6641 25789 6653 25823
rect 6687 25789 6699 25823
rect 7944 25820 7972 25851
rect 8220 25820 8248 25851
rect 8846 25848 8852 25860
rect 8904 25848 8910 25900
rect 9125 25891 9183 25897
rect 9125 25857 9137 25891
rect 9171 25857 9183 25891
rect 9582 25888 9588 25900
rect 9543 25860 9588 25888
rect 9125 25851 9183 25857
rect 9140 25820 9168 25851
rect 9582 25848 9588 25860
rect 9640 25848 9646 25900
rect 9674 25848 9680 25900
rect 9732 25888 9738 25900
rect 9732 25860 9777 25888
rect 9732 25848 9738 25860
rect 7944 25792 8156 25820
rect 8220 25792 9996 25820
rect 6641 25783 6699 25789
rect 5169 25755 5227 25761
rect 5169 25752 5181 25755
rect 4264 25724 5181 25752
rect 5169 25721 5181 25724
rect 5215 25721 5227 25755
rect 6656 25752 6684 25783
rect 6822 25752 6828 25764
rect 6656 25724 6828 25752
rect 5169 25715 5227 25721
rect 6822 25712 6828 25724
rect 6880 25752 6886 25764
rect 7929 25755 7987 25761
rect 7929 25752 7941 25755
rect 6880 25724 7941 25752
rect 6880 25712 6886 25724
rect 7929 25721 7941 25724
rect 7975 25721 7987 25755
rect 8128 25752 8156 25792
rect 8846 25752 8852 25764
rect 8128 25724 8852 25752
rect 7929 25715 7987 25721
rect 8846 25712 8852 25724
rect 8904 25712 8910 25764
rect 9968 25761 9996 25792
rect 9953 25755 10011 25761
rect 9953 25721 9965 25755
rect 9999 25721 10011 25755
rect 10060 25752 10088 25928
rect 10505 25925 10517 25959
rect 10551 25925 10563 25959
rect 10505 25919 10563 25925
rect 10689 25959 10747 25965
rect 10689 25925 10701 25959
rect 10735 25956 10747 25959
rect 10778 25956 10784 25968
rect 10735 25928 10784 25956
rect 10735 25925 10747 25928
rect 10689 25919 10747 25925
rect 10778 25916 10784 25928
rect 10836 25916 10842 25968
rect 12161 25891 12219 25897
rect 12161 25857 12173 25891
rect 12207 25857 12219 25891
rect 12161 25851 12219 25857
rect 12253 25891 12311 25897
rect 12253 25857 12265 25891
rect 12299 25888 12311 25891
rect 12434 25888 12440 25900
rect 12299 25860 12440 25888
rect 12299 25857 12311 25860
rect 12253 25851 12311 25857
rect 12176 25820 12204 25851
rect 12434 25848 12440 25860
rect 12492 25848 12498 25900
rect 12544 25897 12572 25996
rect 12802 25984 12808 26036
rect 12860 26024 12866 26036
rect 13173 26027 13231 26033
rect 13173 26024 13185 26027
rect 12860 25996 13185 26024
rect 12860 25984 12866 25996
rect 13173 25993 13185 25996
rect 13219 25993 13231 26027
rect 13173 25987 13231 25993
rect 13814 25984 13820 26036
rect 13872 25984 13878 26036
rect 14090 26024 14096 26036
rect 14051 25996 14096 26024
rect 14090 25984 14096 25996
rect 14148 25984 14154 26036
rect 15121 26027 15179 26033
rect 15121 26024 15133 26027
rect 14292 25996 15133 26024
rect 12618 25916 12624 25968
rect 12676 25956 12682 25968
rect 13725 25959 13783 25965
rect 13725 25956 13737 25959
rect 12676 25928 13737 25956
rect 12676 25916 12682 25928
rect 13725 25925 13737 25928
rect 13771 25956 13783 25959
rect 13832 25956 13860 25984
rect 14292 25968 14320 25996
rect 15121 25993 15133 25996
rect 15167 25993 15179 26027
rect 15121 25987 15179 25993
rect 17494 25984 17500 26036
rect 17552 26024 17558 26036
rect 18141 26027 18199 26033
rect 18141 26024 18153 26027
rect 17552 25996 18153 26024
rect 17552 25984 17558 25996
rect 18141 25993 18153 25996
rect 18187 25993 18199 26027
rect 19334 26024 19340 26036
rect 18141 25987 18199 25993
rect 18800 25996 19340 26024
rect 14274 25956 14280 25968
rect 13771 25928 14280 25956
rect 13771 25925 13783 25928
rect 13725 25919 13783 25925
rect 14274 25916 14280 25928
rect 14332 25916 14338 25968
rect 14921 25959 14979 25965
rect 14921 25925 14933 25959
rect 14967 25925 14979 25959
rect 14921 25919 14979 25925
rect 17773 25959 17831 25965
rect 17773 25925 17785 25959
rect 17819 25956 17831 25959
rect 18690 25956 18696 25968
rect 17819 25928 18696 25956
rect 17819 25925 17831 25928
rect 17773 25919 17831 25925
rect 12529 25891 12587 25897
rect 12529 25857 12541 25891
rect 12575 25888 12587 25891
rect 12986 25888 12992 25900
rect 12575 25860 12848 25888
rect 12947 25860 12992 25888
rect 12575 25857 12587 25860
rect 12529 25851 12587 25857
rect 12820 25820 12848 25860
rect 12986 25848 12992 25860
rect 13044 25848 13050 25900
rect 13262 25888 13268 25900
rect 13223 25860 13268 25888
rect 13262 25848 13268 25860
rect 13320 25848 13326 25900
rect 13906 25888 13912 25900
rect 13867 25860 13912 25888
rect 13906 25848 13912 25860
rect 13964 25848 13970 25900
rect 14936 25888 14964 25919
rect 18690 25916 18696 25928
rect 18748 25916 18754 25968
rect 15749 25891 15807 25897
rect 15749 25888 15761 25891
rect 14936 25860 15761 25888
rect 15749 25857 15761 25860
rect 15795 25888 15807 25891
rect 15838 25888 15844 25900
rect 15795 25860 15844 25888
rect 15795 25857 15807 25860
rect 15749 25851 15807 25857
rect 15838 25848 15844 25860
rect 15896 25848 15902 25900
rect 16853 25891 16911 25897
rect 16853 25857 16865 25891
rect 16899 25888 16911 25891
rect 17129 25891 17187 25897
rect 17129 25888 17141 25891
rect 16899 25860 17141 25888
rect 16899 25857 16911 25860
rect 16853 25851 16911 25857
rect 17129 25857 17141 25860
rect 17175 25857 17187 25891
rect 17129 25851 17187 25857
rect 17589 25891 17647 25897
rect 17589 25857 17601 25891
rect 17635 25888 17647 25891
rect 17678 25888 17684 25900
rect 17635 25860 17684 25888
rect 17635 25857 17647 25860
rect 17589 25851 17647 25857
rect 13280 25820 13308 25848
rect 12176 25792 12756 25820
rect 12820 25792 13308 25820
rect 12728 25752 12756 25792
rect 13998 25780 14004 25832
rect 14056 25820 14062 25832
rect 16868 25820 16896 25851
rect 17678 25848 17684 25860
rect 17736 25848 17742 25900
rect 17865 25891 17923 25897
rect 17865 25857 17877 25891
rect 17911 25857 17923 25891
rect 17865 25851 17923 25857
rect 14056 25792 16896 25820
rect 17880 25820 17908 25851
rect 17954 25848 17960 25900
rect 18012 25888 18018 25900
rect 18800 25897 18828 25996
rect 19334 25984 19340 25996
rect 19392 25984 19398 26036
rect 19981 26027 20039 26033
rect 19444 25996 19748 26024
rect 19444 25956 19472 25996
rect 18984 25928 19472 25956
rect 19613 25959 19671 25965
rect 18984 25897 19012 25928
rect 19613 25925 19625 25959
rect 19659 25925 19671 25959
rect 19720 25956 19748 25996
rect 19981 25993 19993 26027
rect 20027 26024 20039 26027
rect 20438 26024 20444 26036
rect 20027 25996 20444 26024
rect 20027 25993 20039 25996
rect 19981 25987 20039 25993
rect 20438 25984 20444 25996
rect 20496 25984 20502 26036
rect 22002 25984 22008 26036
rect 22060 25984 22066 26036
rect 22278 25984 22284 26036
rect 22336 26024 22342 26036
rect 22373 26027 22431 26033
rect 22373 26024 22385 26027
rect 22336 25996 22385 26024
rect 22336 25984 22342 25996
rect 22373 25993 22385 25996
rect 22419 25993 22431 26027
rect 24026 26024 24032 26036
rect 22373 25987 22431 25993
rect 23492 25996 24032 26024
rect 20898 25956 20904 25968
rect 19720 25928 20904 25956
rect 19613 25919 19671 25925
rect 18785 25891 18843 25897
rect 18012 25860 18057 25888
rect 18012 25848 18018 25860
rect 18785 25857 18797 25891
rect 18831 25857 18843 25891
rect 18785 25851 18843 25857
rect 18969 25891 19027 25897
rect 18969 25857 18981 25891
rect 19015 25857 19027 25891
rect 18969 25851 19027 25857
rect 19242 25848 19248 25900
rect 19300 25888 19306 25900
rect 19429 25892 19487 25897
rect 19352 25891 19487 25892
rect 19352 25888 19441 25891
rect 19300 25864 19441 25888
rect 19300 25860 19380 25864
rect 19300 25848 19306 25860
rect 19429 25857 19441 25864
rect 19475 25857 19487 25891
rect 19429 25851 19487 25857
rect 19628 25832 19656 25919
rect 20898 25916 20904 25928
rect 20956 25956 20962 25968
rect 22020 25956 22048 25984
rect 20956 25928 22048 25956
rect 20956 25916 20962 25928
rect 22094 25916 22100 25968
rect 22152 25956 22158 25968
rect 22738 25956 22744 25968
rect 22152 25928 22744 25956
rect 22152 25916 22158 25928
rect 22738 25916 22744 25928
rect 22796 25916 22802 25968
rect 23492 25965 23520 25996
rect 24026 25984 24032 25996
rect 24084 25984 24090 26036
rect 24578 26024 24584 26036
rect 24539 25996 24584 26024
rect 24578 25984 24584 25996
rect 24636 25984 24642 26036
rect 25409 26027 25467 26033
rect 25409 25993 25421 26027
rect 25455 26024 25467 26027
rect 26418 26024 26424 26036
rect 25455 25996 26424 26024
rect 25455 25993 25467 25996
rect 25409 25987 25467 25993
rect 26418 25984 26424 25996
rect 26476 25984 26482 26036
rect 23477 25959 23535 25965
rect 23477 25925 23489 25959
rect 23523 25925 23535 25959
rect 24118 25956 24124 25968
rect 23477 25919 23535 25925
rect 23584 25928 24124 25956
rect 19705 25891 19763 25897
rect 19705 25857 19717 25891
rect 19751 25857 19763 25891
rect 19705 25851 19763 25857
rect 18138 25820 18144 25832
rect 17880 25792 18144 25820
rect 14056 25780 14062 25792
rect 18138 25780 18144 25792
rect 18196 25820 18202 25832
rect 18598 25820 18604 25832
rect 18196 25792 18604 25820
rect 18196 25780 18202 25792
rect 18598 25780 18604 25792
rect 18656 25780 18662 25832
rect 19610 25780 19616 25832
rect 19668 25780 19674 25832
rect 19720 25820 19748 25851
rect 19794 25848 19800 25900
rect 19852 25888 19858 25900
rect 19852 25860 19897 25888
rect 19852 25848 19858 25860
rect 19978 25848 19984 25900
rect 20036 25888 20042 25900
rect 20622 25888 20628 25900
rect 20036 25860 20628 25888
rect 20036 25848 20042 25860
rect 20622 25848 20628 25860
rect 20680 25848 20686 25900
rect 21082 25888 21088 25900
rect 21043 25860 21088 25888
rect 21082 25848 21088 25860
rect 21140 25848 21146 25900
rect 21174 25848 21180 25900
rect 21232 25888 21238 25900
rect 21269 25891 21327 25897
rect 21269 25888 21281 25891
rect 21232 25860 21281 25888
rect 21232 25848 21238 25860
rect 21269 25857 21281 25860
rect 21315 25857 21327 25891
rect 21818 25888 21824 25900
rect 21779 25860 21824 25888
rect 21269 25851 21327 25857
rect 21818 25848 21824 25860
rect 21876 25848 21882 25900
rect 21910 25848 21916 25900
rect 21968 25888 21974 25900
rect 22005 25891 22063 25897
rect 22005 25888 22017 25891
rect 21968 25860 22017 25888
rect 21968 25848 21974 25860
rect 22005 25857 22017 25860
rect 22051 25857 22063 25891
rect 22005 25851 22063 25857
rect 22189 25891 22247 25897
rect 22189 25857 22201 25891
rect 22235 25857 22247 25891
rect 23198 25888 23204 25900
rect 23159 25860 23204 25888
rect 22189 25851 22247 25857
rect 20806 25820 20812 25832
rect 19720 25792 20812 25820
rect 20806 25780 20812 25792
rect 20864 25780 20870 25832
rect 12989 25755 13047 25761
rect 12989 25752 13001 25755
rect 10060 25724 12664 25752
rect 12728 25724 13001 25752
rect 9953 25715 10011 25721
rect 1302 25644 1308 25696
rect 1360 25684 1366 25696
rect 1578 25684 1584 25696
rect 1360 25656 1584 25684
rect 1360 25644 1366 25656
rect 1578 25644 1584 25656
rect 1636 25644 1642 25696
rect 3237 25687 3295 25693
rect 3237 25653 3249 25687
rect 3283 25684 3295 25687
rect 4798 25684 4804 25696
rect 3283 25656 4804 25684
rect 3283 25653 3295 25656
rect 3237 25647 3295 25653
rect 4798 25644 4804 25656
rect 4856 25644 4862 25696
rect 4890 25644 4896 25696
rect 4948 25684 4954 25696
rect 6270 25684 6276 25696
rect 4948 25656 6276 25684
rect 4948 25644 4954 25656
rect 6270 25644 6276 25656
rect 6328 25644 6334 25696
rect 6454 25684 6460 25696
rect 6415 25656 6460 25684
rect 6454 25644 6460 25656
rect 6512 25644 6518 25696
rect 6917 25687 6975 25693
rect 6917 25653 6929 25687
rect 6963 25684 6975 25687
rect 7282 25684 7288 25696
rect 6963 25656 7288 25684
rect 6963 25653 6975 25656
rect 6917 25647 6975 25653
rect 7282 25644 7288 25656
rect 7340 25644 7346 25696
rect 9769 25687 9827 25693
rect 9769 25653 9781 25687
rect 9815 25684 9827 25687
rect 9858 25684 9864 25696
rect 9815 25656 9864 25684
rect 9815 25653 9827 25656
rect 9769 25647 9827 25653
rect 9858 25644 9864 25656
rect 9916 25644 9922 25696
rect 12250 25644 12256 25696
rect 12308 25684 12314 25696
rect 12437 25687 12495 25693
rect 12437 25684 12449 25687
rect 12308 25656 12449 25684
rect 12308 25644 12314 25656
rect 12437 25653 12449 25656
rect 12483 25653 12495 25687
rect 12636 25684 12664 25724
rect 12989 25721 13001 25724
rect 13035 25721 13047 25755
rect 12989 25715 13047 25721
rect 13722 25712 13728 25764
rect 13780 25752 13786 25764
rect 15289 25755 15347 25761
rect 15289 25752 15301 25755
rect 13780 25724 15301 25752
rect 13780 25712 13786 25724
rect 15289 25721 15301 25724
rect 15335 25721 15347 25755
rect 15289 25715 15347 25721
rect 16669 25755 16727 25761
rect 16669 25721 16681 25755
rect 16715 25752 16727 25755
rect 17402 25752 17408 25764
rect 16715 25724 17408 25752
rect 16715 25721 16727 25724
rect 16669 25715 16727 25721
rect 17402 25712 17408 25724
rect 17460 25712 17466 25764
rect 18506 25712 18512 25764
rect 18564 25752 18570 25764
rect 21085 25755 21143 25761
rect 21085 25752 21097 25755
rect 18564 25724 21097 25752
rect 18564 25712 18570 25724
rect 21085 25721 21097 25724
rect 21131 25721 21143 25755
rect 21085 25715 21143 25721
rect 14826 25684 14832 25696
rect 12636 25656 14832 25684
rect 12437 25647 12495 25653
rect 14826 25644 14832 25656
rect 14884 25644 14890 25696
rect 15102 25684 15108 25696
rect 15063 25656 15108 25684
rect 15102 25644 15108 25656
rect 15160 25644 15166 25696
rect 15930 25684 15936 25696
rect 15843 25656 15936 25684
rect 15930 25644 15936 25656
rect 15988 25684 15994 25696
rect 16482 25684 16488 25696
rect 15988 25656 16488 25684
rect 15988 25644 15994 25656
rect 16482 25644 16488 25656
rect 16540 25644 16546 25696
rect 18785 25687 18843 25693
rect 18785 25653 18797 25687
rect 18831 25684 18843 25687
rect 19794 25684 19800 25696
rect 18831 25656 19800 25684
rect 18831 25653 18843 25656
rect 18785 25647 18843 25653
rect 19794 25644 19800 25656
rect 19852 25644 19858 25696
rect 20441 25687 20499 25693
rect 20441 25653 20453 25687
rect 20487 25684 20499 25687
rect 20530 25684 20536 25696
rect 20487 25656 20536 25684
rect 20487 25653 20499 25656
rect 20441 25647 20499 25653
rect 20530 25644 20536 25656
rect 20588 25644 20594 25696
rect 22204 25684 22232 25851
rect 23198 25848 23204 25860
rect 23256 25848 23262 25900
rect 23290 25848 23296 25900
rect 23348 25888 23354 25900
rect 23584 25897 23612 25928
rect 24118 25916 24124 25928
rect 24176 25916 24182 25968
rect 23385 25891 23443 25897
rect 23385 25888 23397 25891
rect 23348 25860 23397 25888
rect 23348 25848 23354 25860
rect 23385 25857 23397 25860
rect 23431 25857 23443 25891
rect 23385 25851 23443 25857
rect 23569 25891 23627 25897
rect 23569 25857 23581 25891
rect 23615 25857 23627 25891
rect 24397 25891 24455 25897
rect 24397 25888 24409 25891
rect 23569 25851 23627 25857
rect 23768 25860 24409 25888
rect 23768 25761 23796 25860
rect 24397 25857 24409 25860
rect 24443 25857 24455 25891
rect 24397 25851 24455 25857
rect 24946 25848 24952 25900
rect 25004 25888 25010 25900
rect 25225 25891 25283 25897
rect 25225 25888 25237 25891
rect 25004 25860 25237 25888
rect 25004 25848 25010 25860
rect 25225 25857 25237 25860
rect 25271 25857 25283 25891
rect 25225 25851 25283 25857
rect 26329 25891 26387 25897
rect 26329 25857 26341 25891
rect 26375 25888 26387 25891
rect 26418 25888 26424 25900
rect 26375 25860 26424 25888
rect 26375 25857 26387 25860
rect 26329 25851 26387 25857
rect 26418 25848 26424 25860
rect 26476 25848 26482 25900
rect 27154 25888 27160 25900
rect 27115 25860 27160 25888
rect 27154 25848 27160 25860
rect 27212 25848 27218 25900
rect 24210 25820 24216 25832
rect 24123 25792 24216 25820
rect 24210 25780 24216 25792
rect 24268 25820 24274 25832
rect 25041 25823 25099 25829
rect 25041 25820 25053 25823
rect 24268 25792 25053 25820
rect 24268 25780 24274 25792
rect 25041 25789 25053 25792
rect 25087 25820 25099 25823
rect 26142 25820 26148 25832
rect 25087 25792 26148 25820
rect 25087 25789 25099 25792
rect 25041 25783 25099 25789
rect 26142 25780 26148 25792
rect 26200 25780 26206 25832
rect 23753 25755 23811 25761
rect 23753 25721 23765 25755
rect 23799 25721 23811 25755
rect 23753 25715 23811 25721
rect 22278 25684 22284 25696
rect 22204 25656 22284 25684
rect 22278 25644 22284 25656
rect 22336 25644 22342 25696
rect 24854 25644 24860 25696
rect 24912 25684 24918 25696
rect 26145 25687 26203 25693
rect 26145 25684 26157 25687
rect 24912 25656 26157 25684
rect 24912 25644 24918 25656
rect 26145 25653 26157 25656
rect 26191 25653 26203 25687
rect 26145 25647 26203 25653
rect 26786 25644 26792 25696
rect 26844 25684 26850 25696
rect 26973 25687 27031 25693
rect 26973 25684 26985 25687
rect 26844 25656 26985 25684
rect 26844 25644 26850 25656
rect 26973 25653 26985 25656
rect 27019 25653 27031 25687
rect 26973 25647 27031 25653
rect 1104 25594 28060 25616
rect 1104 25542 5442 25594
rect 5494 25542 5506 25594
rect 5558 25542 5570 25594
rect 5622 25542 5634 25594
rect 5686 25542 5698 25594
rect 5750 25542 14428 25594
rect 14480 25542 14492 25594
rect 14544 25542 14556 25594
rect 14608 25542 14620 25594
rect 14672 25542 14684 25594
rect 14736 25542 23413 25594
rect 23465 25542 23477 25594
rect 23529 25542 23541 25594
rect 23593 25542 23605 25594
rect 23657 25542 23669 25594
rect 23721 25542 28060 25594
rect 1104 25520 28060 25542
rect 1765 25483 1823 25489
rect 1765 25449 1777 25483
rect 1811 25480 1823 25483
rect 2958 25480 2964 25492
rect 1811 25452 2964 25480
rect 1811 25449 1823 25452
rect 1765 25443 1823 25449
rect 2958 25440 2964 25452
rect 3016 25440 3022 25492
rect 4062 25480 4068 25492
rect 3068 25452 4068 25480
rect 2409 25415 2467 25421
rect 2409 25381 2421 25415
rect 2455 25412 2467 25415
rect 3068 25412 3096 25452
rect 4062 25440 4068 25452
rect 4120 25440 4126 25492
rect 4249 25483 4307 25489
rect 4249 25449 4261 25483
rect 4295 25480 4307 25483
rect 4614 25480 4620 25492
rect 4295 25452 4620 25480
rect 4295 25449 4307 25452
rect 4249 25443 4307 25449
rect 4614 25440 4620 25452
rect 4672 25440 4678 25492
rect 5166 25440 5172 25492
rect 5224 25480 5230 25492
rect 9401 25483 9459 25489
rect 9401 25480 9413 25483
rect 5224 25452 9413 25480
rect 5224 25440 5230 25452
rect 9401 25449 9413 25452
rect 9447 25449 9459 25483
rect 9401 25443 9459 25449
rect 9582 25440 9588 25492
rect 9640 25480 9646 25492
rect 9861 25483 9919 25489
rect 9861 25480 9873 25483
rect 9640 25452 9873 25480
rect 9640 25440 9646 25452
rect 9861 25449 9873 25452
rect 9907 25449 9919 25483
rect 9861 25443 9919 25449
rect 12434 25440 12440 25492
rect 12492 25480 12498 25492
rect 12986 25480 12992 25492
rect 12492 25452 12537 25480
rect 12636 25452 12992 25480
rect 12492 25440 12498 25452
rect 4154 25412 4160 25424
rect 2455 25384 3096 25412
rect 3160 25384 4160 25412
rect 2455 25381 2467 25384
rect 2409 25375 2467 25381
rect 3160 25344 3188 25384
rect 4154 25372 4160 25384
rect 4212 25372 4218 25424
rect 7009 25415 7067 25421
rect 7009 25381 7021 25415
rect 7055 25412 7067 25415
rect 7466 25412 7472 25424
rect 7055 25384 7472 25412
rect 7055 25381 7067 25384
rect 7009 25375 7067 25381
rect 7466 25372 7472 25384
rect 7524 25372 7530 25424
rect 7929 25415 7987 25421
rect 7929 25381 7941 25415
rect 7975 25412 7987 25415
rect 8018 25412 8024 25424
rect 7975 25384 8024 25412
rect 7975 25381 7987 25384
rect 7929 25375 7987 25381
rect 8018 25372 8024 25384
rect 8076 25372 8082 25424
rect 10318 25372 10324 25424
rect 10376 25372 10382 25424
rect 4617 25347 4675 25353
rect 4617 25344 4629 25347
rect 1964 25316 3188 25344
rect 3252 25316 4629 25344
rect 1964 25285 1992 25316
rect 3252 25288 3280 25316
rect 4617 25313 4629 25316
rect 4663 25313 4675 25347
rect 4798 25344 4804 25356
rect 4759 25316 4804 25344
rect 4617 25307 4675 25313
rect 4798 25304 4804 25316
rect 4856 25304 4862 25356
rect 4909 25316 5764 25344
rect 1949 25279 2007 25285
rect 1949 25245 1961 25279
rect 1995 25245 2007 25279
rect 1949 25239 2007 25245
rect 2593 25279 2651 25285
rect 2593 25245 2605 25279
rect 2639 25276 2651 25279
rect 3234 25276 3240 25288
rect 2639 25248 2774 25276
rect 3147 25248 3240 25276
rect 2639 25245 2651 25248
rect 2593 25239 2651 25245
rect 2746 25208 2774 25248
rect 3234 25236 3240 25248
rect 3292 25236 3298 25288
rect 4157 25279 4215 25285
rect 4157 25245 4169 25279
rect 4203 25245 4215 25279
rect 4157 25239 4215 25245
rect 4341 25279 4399 25285
rect 4341 25245 4353 25279
rect 4387 25276 4399 25279
rect 4909 25276 4937 25316
rect 5736 25288 5764 25316
rect 5902 25304 5908 25356
rect 5960 25344 5966 25356
rect 5997 25347 6055 25353
rect 5997 25344 6009 25347
rect 5960 25316 6009 25344
rect 5960 25304 5966 25316
rect 5997 25313 6009 25316
rect 6043 25313 6055 25347
rect 10336 25344 10364 25372
rect 5997 25307 6055 25313
rect 9692 25316 10364 25344
rect 5074 25276 5080 25288
rect 4387 25248 4937 25276
rect 5035 25248 5080 25276
rect 4387 25245 4399 25248
rect 4341 25239 4399 25245
rect 3326 25208 3332 25220
rect 2746 25180 3332 25208
rect 3326 25168 3332 25180
rect 3384 25208 3390 25220
rect 3973 25211 4031 25217
rect 3973 25208 3985 25211
rect 3384 25180 3985 25208
rect 3384 25168 3390 25180
rect 3973 25177 3985 25180
rect 4019 25177 4031 25211
rect 4172 25208 4200 25239
rect 5074 25236 5080 25248
rect 5132 25236 5138 25288
rect 5718 25276 5724 25288
rect 5679 25248 5724 25276
rect 5718 25236 5724 25248
rect 5776 25236 5782 25288
rect 5813 25279 5871 25285
rect 5813 25245 5825 25279
rect 5859 25276 5871 25279
rect 6086 25276 6092 25288
rect 5859 25248 6092 25276
rect 5859 25245 5871 25248
rect 5813 25239 5871 25245
rect 5828 25208 5856 25239
rect 6086 25236 6092 25248
rect 6144 25236 6150 25288
rect 6822 25276 6828 25288
rect 6783 25248 6828 25276
rect 6822 25236 6828 25248
rect 6880 25236 6886 25288
rect 9398 25276 9404 25288
rect 9359 25248 9404 25276
rect 9398 25236 9404 25248
rect 9456 25236 9462 25288
rect 9692 25285 9720 25316
rect 12434 25304 12440 25356
rect 12492 25344 12498 25356
rect 12636 25353 12664 25452
rect 12986 25440 12992 25452
rect 13044 25440 13050 25492
rect 13078 25440 13084 25492
rect 13136 25480 13142 25492
rect 14369 25483 14427 25489
rect 14369 25480 14381 25483
rect 13136 25452 14381 25480
rect 13136 25440 13142 25452
rect 14369 25449 14381 25452
rect 14415 25480 14427 25483
rect 14415 25452 14780 25480
rect 14415 25449 14427 25452
rect 14369 25443 14427 25449
rect 14274 25372 14280 25424
rect 14332 25412 14338 25424
rect 14553 25415 14611 25421
rect 14553 25412 14565 25415
rect 14332 25384 14565 25412
rect 14332 25372 14338 25384
rect 14553 25381 14565 25384
rect 14599 25381 14611 25415
rect 14553 25375 14611 25381
rect 12621 25347 12679 25353
rect 12621 25344 12633 25347
rect 12492 25316 12633 25344
rect 12492 25304 12498 25316
rect 12621 25313 12633 25316
rect 12667 25313 12679 25347
rect 12802 25344 12808 25356
rect 12763 25316 12808 25344
rect 12621 25307 12679 25313
rect 12802 25304 12808 25316
rect 12860 25304 12866 25356
rect 14752 25344 14780 25452
rect 15102 25440 15108 25492
rect 15160 25480 15166 25492
rect 15841 25483 15899 25489
rect 15841 25480 15853 25483
rect 15160 25452 15853 25480
rect 15160 25440 15166 25452
rect 15841 25449 15853 25452
rect 15887 25480 15899 25483
rect 15887 25452 16804 25480
rect 15887 25449 15899 25452
rect 15841 25443 15899 25449
rect 14826 25372 14832 25424
rect 14884 25412 14890 25424
rect 15286 25412 15292 25424
rect 14884 25384 15292 25412
rect 14884 25372 14890 25384
rect 15286 25372 15292 25384
rect 15344 25372 15350 25424
rect 16298 25412 16304 25424
rect 15396 25384 16304 25412
rect 15396 25344 15424 25384
rect 16298 25372 16304 25384
rect 16356 25372 16362 25424
rect 16776 25421 16804 25452
rect 19610 25440 19616 25492
rect 19668 25480 19674 25492
rect 19705 25483 19763 25489
rect 19705 25480 19717 25483
rect 19668 25452 19717 25480
rect 19668 25440 19674 25452
rect 19705 25449 19717 25452
rect 19751 25449 19763 25483
rect 19705 25443 19763 25449
rect 22373 25483 22431 25489
rect 22373 25449 22385 25483
rect 22419 25480 22431 25483
rect 22462 25480 22468 25492
rect 22419 25452 22468 25480
rect 22419 25449 22431 25452
rect 22373 25443 22431 25449
rect 22462 25440 22468 25452
rect 22520 25440 22526 25492
rect 24946 25480 24952 25492
rect 24907 25452 24952 25480
rect 24946 25440 24952 25452
rect 25004 25440 25010 25492
rect 16761 25415 16819 25421
rect 16761 25381 16773 25415
rect 16807 25381 16819 25415
rect 16761 25375 16819 25381
rect 17862 25372 17868 25424
rect 17920 25372 17926 25424
rect 22738 25412 22744 25424
rect 18432 25384 22744 25412
rect 14752 25316 15424 25344
rect 15657 25347 15715 25353
rect 15657 25313 15669 25347
rect 15703 25344 15715 25347
rect 17880 25344 17908 25372
rect 15703 25316 17908 25344
rect 15703 25313 15715 25316
rect 15657 25307 15715 25313
rect 17954 25304 17960 25356
rect 18012 25344 18018 25356
rect 18141 25347 18199 25353
rect 18141 25344 18153 25347
rect 18012 25316 18153 25344
rect 18012 25304 18018 25316
rect 18141 25313 18153 25316
rect 18187 25313 18199 25347
rect 18141 25307 18199 25313
rect 9585 25279 9643 25285
rect 9585 25245 9597 25279
rect 9631 25245 9643 25279
rect 9585 25239 9643 25245
rect 9677 25279 9735 25285
rect 9677 25245 9689 25279
rect 9723 25245 9735 25279
rect 9677 25239 9735 25245
rect 10321 25279 10379 25285
rect 10321 25245 10333 25279
rect 10367 25276 10379 25279
rect 10962 25276 10968 25288
rect 10367 25248 10968 25276
rect 10367 25245 10379 25248
rect 10321 25239 10379 25245
rect 4172 25180 5856 25208
rect 5997 25211 6055 25217
rect 3973 25171 4031 25177
rect 5997 25177 6009 25211
rect 6043 25208 6055 25211
rect 6362 25208 6368 25220
rect 6043 25180 6368 25208
rect 6043 25177 6055 25180
rect 5997 25171 6055 25177
rect 6362 25168 6368 25180
rect 6420 25168 6426 25220
rect 7558 25168 7564 25220
rect 7616 25208 7622 25220
rect 7745 25211 7803 25217
rect 7745 25208 7757 25211
rect 7616 25180 7757 25208
rect 7616 25168 7622 25180
rect 7745 25177 7757 25180
rect 7791 25177 7803 25211
rect 7745 25171 7803 25177
rect 3050 25140 3056 25152
rect 3011 25112 3056 25140
rect 3050 25100 3056 25112
rect 3108 25100 3114 25152
rect 4246 25100 4252 25152
rect 4304 25140 4310 25152
rect 4706 25140 4712 25152
rect 4304 25112 4712 25140
rect 4304 25100 4310 25112
rect 4706 25100 4712 25112
rect 4764 25140 4770 25152
rect 5350 25140 5356 25152
rect 4764 25112 5356 25140
rect 4764 25100 4770 25112
rect 5350 25100 5356 25112
rect 5408 25100 5414 25152
rect 9600 25140 9628 25239
rect 10962 25236 10968 25248
rect 11020 25276 11026 25288
rect 11790 25276 11796 25288
rect 11020 25248 11796 25276
rect 11020 25236 11026 25248
rect 11790 25236 11796 25248
rect 11848 25236 11854 25288
rect 12713 25279 12771 25285
rect 12713 25245 12725 25279
rect 12759 25245 12771 25279
rect 12894 25276 12900 25288
rect 12855 25248 12900 25276
rect 12713 25239 12771 25245
rect 10588 25211 10646 25217
rect 10588 25177 10600 25211
rect 10634 25208 10646 25211
rect 10870 25208 10876 25220
rect 10634 25180 10876 25208
rect 10634 25177 10646 25180
rect 10588 25171 10646 25177
rect 10870 25168 10876 25180
rect 10928 25168 10934 25220
rect 12728 25208 12756 25239
rect 12894 25236 12900 25248
rect 12952 25236 12958 25288
rect 13262 25276 13268 25288
rect 13096 25248 13268 25276
rect 13096 25208 13124 25248
rect 13262 25236 13268 25248
rect 13320 25276 13326 25288
rect 15565 25279 15623 25285
rect 15565 25276 15577 25279
rect 13320 25248 15577 25276
rect 13320 25236 13326 25248
rect 15565 25245 15577 25248
rect 15611 25276 15623 25279
rect 15838 25276 15844 25288
rect 15611 25248 15844 25276
rect 15611 25245 15623 25248
rect 15565 25239 15623 25245
rect 15838 25236 15844 25248
rect 15896 25236 15902 25288
rect 16390 25236 16396 25288
rect 16448 25276 16454 25288
rect 17865 25279 17923 25285
rect 17865 25276 17877 25279
rect 16448 25248 17877 25276
rect 16448 25236 16454 25248
rect 17865 25245 17877 25248
rect 17911 25276 17923 25279
rect 18432 25276 18460 25384
rect 22738 25372 22744 25384
rect 22796 25372 22802 25424
rect 20346 25344 20352 25356
rect 20307 25316 20352 25344
rect 20346 25304 20352 25316
rect 20404 25304 20410 25356
rect 22278 25344 22284 25356
rect 22191 25316 22284 25344
rect 17911 25248 18460 25276
rect 17911 25245 17923 25248
rect 17865 25239 17923 25245
rect 19886 25236 19892 25288
rect 19944 25276 19950 25288
rect 21082 25276 21088 25288
rect 19944 25248 21088 25276
rect 19944 25236 19950 25248
rect 21082 25236 21088 25248
rect 21140 25236 21146 25288
rect 21358 25276 21364 25288
rect 21319 25248 21364 25276
rect 21358 25236 21364 25248
rect 21416 25236 21422 25288
rect 21818 25276 21824 25288
rect 21779 25248 21824 25276
rect 21818 25236 21824 25248
rect 21876 25236 21882 25288
rect 22204 25285 22232 25316
rect 22278 25304 22284 25316
rect 22336 25344 22342 25356
rect 23293 25347 23351 25353
rect 23293 25344 23305 25347
rect 22336 25316 23305 25344
rect 22336 25304 22342 25316
rect 23293 25313 23305 25316
rect 23339 25344 23351 25347
rect 24118 25344 24124 25356
rect 23339 25316 24124 25344
rect 23339 25313 23351 25316
rect 23293 25307 23351 25313
rect 24118 25304 24124 25316
rect 24176 25344 24182 25356
rect 25406 25344 25412 25356
rect 24176 25316 24808 25344
rect 25367 25316 25412 25344
rect 24176 25304 24182 25316
rect 22189 25279 22247 25285
rect 22189 25245 22201 25279
rect 22235 25245 22247 25279
rect 22189 25239 22247 25245
rect 22738 25236 22744 25288
rect 22796 25276 22802 25288
rect 23017 25279 23075 25285
rect 23017 25276 23029 25279
rect 22796 25248 23029 25276
rect 22796 25236 22802 25248
rect 23017 25245 23029 25248
rect 23063 25245 23075 25279
rect 24394 25276 24400 25288
rect 24355 25248 24400 25276
rect 23017 25239 23075 25245
rect 24394 25236 24400 25248
rect 24452 25236 24458 25288
rect 24578 25276 24584 25288
rect 24539 25248 24584 25276
rect 24578 25236 24584 25248
rect 24636 25236 24642 25288
rect 24780 25285 24808 25316
rect 25406 25304 25412 25316
rect 25464 25304 25470 25356
rect 24765 25279 24823 25285
rect 24765 25245 24777 25279
rect 24811 25276 24823 25279
rect 24946 25276 24952 25288
rect 24811 25248 24952 25276
rect 24811 25245 24823 25248
rect 24765 25239 24823 25245
rect 24946 25236 24952 25248
rect 25004 25236 25010 25288
rect 25676 25279 25734 25285
rect 25676 25245 25688 25279
rect 25722 25276 25734 25279
rect 26234 25276 26240 25288
rect 25722 25248 26240 25276
rect 25722 25245 25734 25248
rect 25676 25239 25734 25245
rect 26234 25236 26240 25248
rect 26292 25236 26298 25288
rect 14182 25208 14188 25220
rect 12728 25180 13124 25208
rect 14143 25180 14188 25208
rect 14182 25168 14188 25180
rect 14240 25168 14246 25220
rect 16485 25211 16543 25217
rect 16485 25177 16497 25211
rect 16531 25208 16543 25211
rect 16850 25208 16856 25220
rect 16531 25180 16856 25208
rect 16531 25177 16543 25180
rect 16485 25171 16543 25177
rect 16850 25168 16856 25180
rect 16908 25168 16914 25220
rect 20073 25211 20131 25217
rect 20073 25177 20085 25211
rect 20119 25208 20131 25211
rect 20806 25208 20812 25220
rect 20119 25180 20812 25208
rect 20119 25177 20131 25180
rect 20073 25171 20131 25177
rect 20806 25168 20812 25180
rect 20864 25168 20870 25220
rect 22002 25208 22008 25220
rect 21963 25180 22008 25208
rect 22002 25168 22008 25180
rect 22060 25168 22066 25220
rect 22097 25211 22155 25217
rect 22097 25177 22109 25211
rect 22143 25208 22155 25211
rect 22462 25208 22468 25220
rect 22143 25180 22468 25208
rect 22143 25177 22155 25180
rect 22097 25171 22155 25177
rect 22462 25168 22468 25180
rect 22520 25208 22526 25220
rect 24670 25217 24676 25220
rect 22520 25180 23060 25208
rect 22520 25168 22526 25180
rect 23032 25152 23060 25180
rect 24669 25171 24676 25217
rect 24728 25208 24734 25220
rect 24728 25180 26832 25208
rect 24670 25168 24676 25171
rect 24728 25168 24734 25180
rect 10962 25140 10968 25152
rect 9600 25112 10968 25140
rect 10962 25100 10968 25112
rect 11020 25140 11026 25152
rect 11701 25143 11759 25149
rect 11701 25140 11713 25143
rect 11020 25112 11713 25140
rect 11020 25100 11026 25112
rect 11701 25109 11713 25112
rect 11747 25109 11759 25143
rect 11701 25103 11759 25109
rect 14395 25143 14453 25149
rect 14395 25109 14407 25143
rect 14441 25140 14453 25143
rect 15194 25140 15200 25152
rect 14441 25112 15200 25140
rect 14441 25109 14453 25112
rect 14395 25103 14453 25109
rect 15194 25100 15200 25112
rect 15252 25100 15258 25152
rect 16942 25140 16948 25152
rect 16903 25112 16948 25140
rect 16942 25100 16948 25112
rect 17000 25100 17006 25152
rect 20162 25140 20168 25152
rect 20123 25112 20168 25140
rect 20162 25100 20168 25112
rect 20220 25100 20226 25152
rect 21177 25143 21235 25149
rect 21177 25109 21189 25143
rect 21223 25140 21235 25143
rect 21726 25140 21732 25152
rect 21223 25112 21732 25140
rect 21223 25109 21235 25112
rect 21177 25103 21235 25109
rect 21726 25100 21732 25112
rect 21784 25100 21790 25152
rect 23014 25100 23020 25152
rect 23072 25100 23078 25152
rect 26804 25149 26832 25180
rect 26789 25143 26847 25149
rect 26789 25109 26801 25143
rect 26835 25109 26847 25143
rect 26789 25103 26847 25109
rect 1104 25050 28060 25072
rect 1104 24998 9935 25050
rect 9987 24998 9999 25050
rect 10051 24998 10063 25050
rect 10115 24998 10127 25050
rect 10179 24998 10191 25050
rect 10243 24998 18920 25050
rect 18972 24998 18984 25050
rect 19036 24998 19048 25050
rect 19100 24998 19112 25050
rect 19164 24998 19176 25050
rect 19228 24998 28060 25050
rect 1104 24976 28060 24998
rect 3145 24939 3203 24945
rect 3145 24905 3157 24939
rect 3191 24936 3203 24939
rect 5635 24939 5693 24945
rect 3191 24908 4568 24936
rect 3191 24905 3203 24908
rect 3145 24899 3203 24905
rect 2240 24840 2544 24868
rect 1765 24803 1823 24809
rect 1765 24769 1777 24803
rect 1811 24800 1823 24803
rect 2240 24800 2268 24840
rect 2406 24800 2412 24812
rect 1811 24772 2268 24800
rect 2367 24772 2412 24800
rect 1811 24769 1823 24772
rect 1765 24763 1823 24769
rect 2406 24760 2412 24772
rect 2464 24760 2470 24812
rect 2516 24800 2544 24840
rect 3160 24800 3188 24899
rect 3510 24868 3516 24880
rect 3252 24840 3516 24868
rect 3252 24809 3280 24840
rect 3510 24828 3516 24840
rect 3568 24868 3574 24880
rect 3970 24868 3976 24880
rect 3568 24840 3976 24868
rect 3568 24828 3574 24840
rect 3970 24828 3976 24840
rect 4028 24828 4034 24880
rect 2516 24772 3188 24800
rect 3237 24803 3295 24809
rect 3237 24769 3249 24803
rect 3283 24769 3295 24803
rect 3789 24803 3847 24809
rect 3789 24800 3801 24803
rect 3237 24763 3295 24769
rect 3344 24772 3801 24800
rect 1302 24692 1308 24744
rect 1360 24732 1366 24744
rect 3344 24732 3372 24772
rect 3789 24769 3801 24772
rect 3835 24769 3847 24803
rect 3789 24763 3847 24769
rect 4062 24760 4068 24812
rect 4120 24800 4126 24812
rect 4433 24803 4491 24809
rect 4433 24800 4445 24803
rect 4120 24772 4445 24800
rect 4120 24760 4126 24772
rect 4433 24769 4445 24772
rect 4479 24769 4491 24803
rect 4540 24800 4568 24908
rect 5635 24905 5647 24939
rect 5681 24936 5693 24939
rect 5810 24936 5816 24948
rect 5681 24908 5816 24936
rect 5681 24905 5693 24908
rect 5635 24899 5693 24905
rect 5810 24896 5816 24908
rect 5868 24896 5874 24948
rect 6454 24896 6460 24948
rect 6512 24936 6518 24948
rect 6733 24939 6791 24945
rect 6733 24936 6745 24939
rect 6512 24908 6745 24936
rect 6512 24896 6518 24908
rect 6733 24905 6745 24908
rect 6779 24905 6791 24939
rect 6733 24899 6791 24905
rect 9217 24939 9275 24945
rect 9217 24905 9229 24939
rect 9263 24936 9275 24939
rect 9306 24936 9312 24948
rect 9263 24908 9312 24936
rect 9263 24905 9275 24908
rect 9217 24899 9275 24905
rect 9306 24896 9312 24908
rect 9364 24896 9370 24948
rect 9766 24896 9772 24948
rect 9824 24936 9830 24948
rect 10229 24939 10287 24945
rect 10229 24936 10241 24939
rect 9824 24908 10241 24936
rect 9824 24896 9830 24908
rect 10229 24905 10241 24908
rect 10275 24905 10287 24939
rect 10870 24936 10876 24948
rect 10831 24908 10876 24936
rect 10229 24899 10287 24905
rect 10870 24896 10876 24908
rect 10928 24896 10934 24948
rect 11701 24939 11759 24945
rect 11701 24905 11713 24939
rect 11747 24936 11759 24939
rect 12434 24936 12440 24948
rect 11747 24908 12440 24936
rect 11747 24905 11759 24908
rect 11701 24899 11759 24905
rect 12434 24896 12440 24908
rect 12492 24896 12498 24948
rect 13078 24936 13084 24948
rect 12820 24908 13084 24936
rect 4617 24871 4675 24877
rect 4617 24837 4629 24871
rect 4663 24868 4675 24871
rect 4798 24868 4804 24880
rect 4663 24840 4804 24868
rect 4663 24837 4675 24840
rect 4617 24831 4675 24837
rect 4798 24828 4804 24840
rect 4856 24828 4862 24880
rect 7466 24868 7472 24880
rect 5828 24840 6500 24868
rect 7427 24840 7472 24868
rect 4890 24800 4896 24812
rect 4540 24772 4896 24800
rect 4433 24763 4491 24769
rect 4890 24760 4896 24772
rect 4948 24760 4954 24812
rect 5534 24800 5540 24812
rect 5495 24772 5540 24800
rect 5534 24760 5540 24772
rect 5592 24760 5598 24812
rect 5718 24800 5724 24812
rect 5631 24772 5724 24800
rect 5718 24760 5724 24772
rect 5776 24760 5782 24812
rect 5828 24809 5856 24840
rect 5813 24803 5871 24809
rect 5813 24769 5825 24803
rect 5859 24769 5871 24803
rect 5813 24763 5871 24769
rect 5902 24760 5908 24812
rect 5960 24800 5966 24812
rect 6365 24803 6423 24809
rect 6365 24800 6377 24803
rect 5960 24772 6377 24800
rect 5960 24760 5966 24772
rect 6365 24769 6377 24772
rect 6411 24769 6423 24803
rect 6472 24800 6500 24840
rect 7466 24828 7472 24840
rect 7524 24828 7530 24880
rect 12618 24868 12624 24880
rect 9324 24840 9720 24868
rect 7650 24800 7656 24812
rect 6472 24772 6664 24800
rect 7611 24772 7656 24800
rect 6365 24763 6423 24769
rect 1360 24704 3372 24732
rect 1360 24692 1366 24704
rect 3418 24692 3424 24744
rect 3476 24692 3482 24744
rect 3513 24735 3571 24741
rect 3513 24701 3525 24735
rect 3559 24701 3571 24735
rect 3513 24695 3571 24701
rect 2406 24624 2412 24676
rect 2464 24664 2470 24676
rect 2777 24667 2835 24673
rect 2777 24664 2789 24667
rect 2464 24636 2789 24664
rect 2464 24624 2470 24636
rect 2777 24633 2789 24636
rect 2823 24664 2835 24667
rect 3142 24664 3148 24676
rect 2823 24636 3148 24664
rect 2823 24633 2835 24636
rect 2777 24627 2835 24633
rect 3142 24624 3148 24636
rect 3200 24624 3206 24676
rect 3329 24667 3387 24673
rect 3329 24633 3341 24667
rect 3375 24664 3387 24667
rect 3436 24664 3464 24692
rect 3375 24636 3464 24664
rect 3528 24664 3556 24695
rect 3694 24692 3700 24744
rect 3752 24732 3758 24744
rect 5626 24732 5632 24744
rect 3752 24704 5632 24732
rect 3752 24692 3758 24704
rect 5626 24692 5632 24704
rect 5684 24692 5690 24744
rect 5736 24732 5764 24760
rect 6178 24732 6184 24744
rect 5736 24704 6184 24732
rect 6178 24692 6184 24704
rect 6236 24732 6242 24744
rect 6454 24732 6460 24744
rect 6236 24704 6460 24732
rect 6236 24692 6242 24704
rect 6454 24692 6460 24704
rect 6512 24692 6518 24744
rect 3786 24664 3792 24676
rect 3528 24636 3792 24664
rect 3375 24633 3387 24636
rect 3329 24627 3387 24633
rect 3786 24624 3792 24636
rect 3844 24624 3850 24676
rect 6086 24624 6092 24676
rect 6144 24664 6150 24676
rect 6636 24664 6664 24772
rect 7650 24760 7656 24772
rect 7708 24760 7714 24812
rect 7742 24760 7748 24812
rect 7800 24800 7806 24812
rect 8205 24803 8263 24809
rect 7800 24772 7845 24800
rect 7800 24760 7806 24772
rect 8205 24769 8217 24803
rect 8251 24800 8263 24803
rect 8754 24800 8760 24812
rect 8251 24772 8760 24800
rect 8251 24769 8263 24772
rect 8205 24763 8263 24769
rect 8754 24760 8760 24772
rect 8812 24760 8818 24812
rect 9033 24803 9091 24809
rect 9033 24769 9045 24803
rect 9079 24800 9091 24803
rect 9324 24800 9352 24840
rect 9079 24772 9352 24800
rect 9401 24803 9459 24809
rect 9079 24769 9091 24772
rect 9033 24763 9091 24769
rect 9401 24769 9413 24803
rect 9447 24769 9459 24803
rect 9582 24800 9588 24812
rect 9543 24772 9588 24800
rect 9401 24763 9459 24769
rect 6914 24692 6920 24744
rect 6972 24732 6978 24744
rect 6972 24704 8432 24732
rect 6972 24692 6978 24704
rect 7469 24667 7527 24673
rect 7469 24664 7481 24667
rect 6144 24636 6408 24664
rect 6636 24636 7481 24664
rect 6144 24624 6150 24636
rect 1581 24599 1639 24605
rect 1581 24565 1593 24599
rect 1627 24596 1639 24599
rect 1946 24596 1952 24608
rect 1627 24568 1952 24596
rect 1627 24565 1639 24568
rect 1581 24559 1639 24565
rect 1946 24556 1952 24568
rect 2004 24556 2010 24608
rect 2225 24599 2283 24605
rect 2225 24565 2237 24599
rect 2271 24596 2283 24599
rect 2958 24596 2964 24608
rect 2271 24568 2964 24596
rect 2271 24565 2283 24568
rect 2225 24559 2283 24565
rect 2958 24556 2964 24568
rect 3016 24556 3022 24608
rect 3418 24556 3424 24608
rect 3476 24596 3482 24608
rect 3605 24599 3663 24605
rect 3476 24568 3521 24596
rect 3476 24556 3482 24568
rect 3605 24565 3617 24599
rect 3651 24596 3663 24599
rect 3694 24596 3700 24608
rect 3651 24568 3700 24596
rect 3651 24565 3663 24568
rect 3605 24559 3663 24565
rect 3694 24556 3700 24568
rect 3752 24556 3758 24608
rect 4154 24556 4160 24608
rect 4212 24596 4218 24608
rect 4249 24599 4307 24605
rect 4249 24596 4261 24599
rect 4212 24568 4261 24596
rect 4212 24556 4218 24568
rect 4249 24565 4261 24568
rect 4295 24565 4307 24599
rect 4249 24559 4307 24565
rect 4801 24599 4859 24605
rect 4801 24565 4813 24599
rect 4847 24596 4859 24599
rect 6178 24596 6184 24608
rect 4847 24568 6184 24596
rect 4847 24565 4859 24568
rect 4801 24559 4859 24565
rect 6178 24556 6184 24568
rect 6236 24556 6242 24608
rect 6380 24605 6408 24636
rect 7469 24633 7481 24636
rect 7515 24633 7527 24667
rect 7469 24627 7527 24633
rect 7834 24624 7840 24676
rect 7892 24664 7898 24676
rect 8404 24673 8432 24704
rect 8478 24692 8484 24744
rect 8536 24732 8542 24744
rect 9416 24732 9444 24763
rect 9582 24760 9588 24772
rect 9640 24760 9646 24812
rect 9692 24800 9720 24840
rect 11624 24840 12624 24868
rect 10137 24803 10195 24809
rect 9692 24772 10088 24800
rect 9674 24732 9680 24744
rect 8536 24704 8581 24732
rect 9416 24704 9680 24732
rect 8536 24692 8542 24704
rect 9674 24692 9680 24704
rect 9732 24692 9738 24744
rect 10060 24732 10088 24772
rect 10137 24769 10149 24803
rect 10183 24800 10195 24803
rect 10318 24800 10324 24812
rect 10183 24772 10324 24800
rect 10183 24769 10195 24772
rect 10137 24763 10195 24769
rect 10318 24760 10324 24772
rect 10376 24760 10382 24812
rect 10778 24800 10784 24812
rect 10739 24772 10784 24800
rect 10778 24760 10784 24772
rect 10836 24760 10842 24812
rect 10870 24760 10876 24812
rect 10928 24800 10934 24812
rect 10965 24803 11023 24809
rect 10965 24800 10977 24803
rect 10928 24772 10977 24800
rect 10928 24760 10934 24772
rect 10965 24769 10977 24772
rect 11011 24800 11023 24803
rect 11146 24800 11152 24812
rect 11011 24772 11152 24800
rect 11011 24769 11023 24772
rect 10965 24763 11023 24769
rect 11146 24760 11152 24772
rect 11204 24760 11210 24812
rect 11517 24803 11575 24809
rect 11517 24769 11529 24803
rect 11563 24800 11575 24803
rect 11624 24800 11652 24840
rect 12618 24828 12624 24840
rect 12676 24828 12682 24880
rect 12820 24877 12848 24908
rect 13078 24896 13084 24908
rect 13136 24896 13142 24948
rect 18690 24936 18696 24948
rect 18651 24908 18696 24936
rect 18690 24896 18696 24908
rect 18748 24896 18754 24948
rect 19153 24939 19211 24945
rect 19153 24936 19165 24939
rect 18800 24908 19165 24936
rect 12805 24871 12863 24877
rect 12805 24837 12817 24871
rect 12851 24837 12863 24871
rect 16761 24871 16819 24877
rect 12805 24831 12863 24837
rect 13035 24837 13093 24843
rect 11563 24772 11652 24800
rect 11701 24803 11759 24809
rect 11563 24769 11575 24772
rect 11517 24763 11575 24769
rect 11701 24769 11713 24803
rect 11747 24800 11759 24803
rect 12066 24800 12072 24812
rect 11747 24772 12072 24800
rect 11747 24769 11759 24772
rect 11701 24763 11759 24769
rect 12066 24760 12072 24772
rect 12124 24760 12130 24812
rect 12161 24803 12219 24809
rect 12161 24769 12173 24803
rect 12207 24769 12219 24803
rect 12342 24800 12348 24812
rect 12303 24772 12348 24800
rect 12161 24763 12219 24769
rect 10686 24732 10692 24744
rect 10060 24704 10692 24732
rect 10686 24692 10692 24704
rect 10744 24692 10750 24744
rect 12176 24732 12204 24763
rect 12342 24760 12348 24772
rect 12400 24760 12406 24812
rect 13035 24803 13047 24837
rect 13081 24803 13093 24837
rect 16761 24837 16773 24871
rect 16807 24868 16819 24871
rect 16807 24840 18000 24868
rect 16807 24837 16819 24840
rect 16761 24831 16819 24837
rect 13035 24800 13093 24803
rect 12535 24797 13093 24800
rect 12535 24772 13078 24797
rect 12535 24732 12563 24772
rect 13538 24760 13544 24812
rect 13596 24800 13602 24812
rect 13633 24803 13691 24809
rect 13633 24800 13645 24803
rect 13596 24772 13645 24800
rect 13596 24760 13602 24772
rect 13633 24769 13645 24772
rect 13679 24800 13691 24803
rect 14182 24800 14188 24812
rect 13679 24772 14188 24800
rect 13679 24769 13691 24772
rect 13633 24763 13691 24769
rect 14182 24760 14188 24772
rect 14240 24800 14246 24812
rect 14369 24803 14427 24809
rect 14369 24800 14381 24803
rect 14240 24772 14381 24800
rect 14240 24760 14246 24772
rect 14369 24769 14381 24772
rect 14415 24769 14427 24803
rect 15194 24800 15200 24812
rect 15155 24772 15200 24800
rect 14369 24763 14427 24769
rect 15194 24760 15200 24772
rect 15252 24760 15258 24812
rect 16669 24803 16727 24809
rect 16669 24769 16681 24803
rect 16715 24769 16727 24803
rect 16669 24763 16727 24769
rect 16853 24803 16911 24809
rect 16853 24769 16865 24803
rect 16899 24800 16911 24803
rect 17494 24800 17500 24812
rect 16899 24772 17500 24800
rect 16899 24769 16911 24772
rect 16853 24763 16911 24769
rect 12084 24704 12563 24732
rect 12084 24676 12112 24704
rect 12618 24692 12624 24744
rect 12676 24732 12682 24744
rect 12802 24732 12808 24744
rect 12676 24704 12808 24732
rect 12676 24692 12682 24704
rect 12802 24692 12808 24704
rect 12860 24732 12866 24744
rect 15289 24735 15347 24741
rect 12860 24704 14596 24732
rect 12860 24692 12866 24704
rect 8297 24667 8355 24673
rect 8297 24664 8309 24667
rect 7892 24636 8309 24664
rect 7892 24624 7898 24636
rect 8297 24633 8309 24636
rect 8343 24633 8355 24667
rect 8297 24627 8355 24633
rect 8389 24667 8447 24673
rect 8389 24633 8401 24667
rect 8435 24633 8447 24667
rect 9858 24664 9864 24676
rect 8389 24627 8447 24633
rect 9416 24636 9864 24664
rect 6365 24599 6423 24605
rect 6365 24565 6377 24599
rect 6411 24565 6423 24599
rect 6365 24559 6423 24565
rect 6914 24556 6920 24608
rect 6972 24596 6978 24608
rect 9416 24605 9444 24636
rect 9858 24624 9864 24636
rect 9916 24624 9922 24676
rect 12066 24624 12072 24676
rect 12124 24624 12130 24676
rect 12250 24664 12256 24676
rect 12211 24636 12256 24664
rect 12250 24624 12256 24636
rect 12308 24624 12314 24676
rect 13170 24664 13176 24676
rect 13131 24636 13176 24664
rect 13170 24624 13176 24636
rect 13228 24624 13234 24676
rect 14568 24673 14596 24704
rect 15289 24701 15301 24735
rect 15335 24732 15347 24735
rect 16684 24732 16712 24763
rect 17494 24760 17500 24772
rect 17552 24760 17558 24812
rect 17678 24800 17684 24812
rect 17639 24772 17684 24800
rect 17678 24760 17684 24772
rect 17736 24760 17742 24812
rect 15335 24704 16252 24732
rect 16684 24704 17172 24732
rect 15335 24701 15347 24704
rect 15289 24695 15347 24701
rect 14553 24667 14611 24673
rect 14553 24633 14565 24667
rect 14599 24664 14611 24667
rect 15378 24664 15384 24676
rect 14599 24636 15384 24664
rect 14599 24633 14611 24636
rect 14553 24627 14611 24633
rect 15378 24624 15384 24636
rect 15436 24624 15442 24676
rect 9401 24599 9459 24605
rect 9401 24596 9413 24599
rect 6972 24568 9413 24596
rect 6972 24556 6978 24568
rect 9401 24565 9413 24568
rect 9447 24565 9459 24599
rect 9401 24559 9459 24565
rect 11514 24556 11520 24608
rect 11572 24596 11578 24608
rect 12342 24596 12348 24608
rect 11572 24568 12348 24596
rect 11572 24556 11578 24568
rect 12342 24556 12348 24568
rect 12400 24596 12406 24608
rect 12894 24596 12900 24608
rect 12400 24568 12900 24596
rect 12400 24556 12406 24568
rect 12894 24556 12900 24568
rect 12952 24596 12958 24608
rect 12989 24599 13047 24605
rect 12989 24596 13001 24599
rect 12952 24568 13001 24596
rect 12952 24556 12958 24568
rect 12989 24565 13001 24568
rect 13035 24565 13047 24599
rect 12989 24559 13047 24565
rect 13630 24556 13636 24608
rect 13688 24596 13694 24608
rect 13725 24599 13783 24605
rect 13725 24596 13737 24599
rect 13688 24568 13737 24596
rect 13688 24556 13694 24568
rect 13725 24565 13737 24568
rect 13771 24596 13783 24599
rect 13906 24596 13912 24608
rect 13771 24568 13912 24596
rect 13771 24565 13783 24568
rect 13725 24559 13783 24565
rect 13906 24556 13912 24568
rect 13964 24556 13970 24608
rect 15473 24599 15531 24605
rect 15473 24565 15485 24599
rect 15519 24596 15531 24599
rect 15654 24596 15660 24608
rect 15519 24568 15660 24596
rect 15519 24565 15531 24568
rect 15473 24559 15531 24565
rect 15654 24556 15660 24568
rect 15712 24556 15718 24608
rect 16224 24596 16252 24704
rect 16850 24596 16856 24608
rect 16224 24568 16856 24596
rect 16850 24556 16856 24568
rect 16908 24556 16914 24608
rect 17144 24596 17172 24704
rect 17218 24692 17224 24744
rect 17276 24732 17282 24744
rect 17405 24735 17463 24741
rect 17405 24732 17417 24735
rect 17276 24704 17417 24732
rect 17276 24692 17282 24704
rect 17405 24701 17417 24704
rect 17451 24701 17463 24735
rect 17405 24695 17463 24701
rect 17972 24664 18000 24840
rect 18598 24828 18604 24880
rect 18656 24868 18662 24880
rect 18800 24868 18828 24908
rect 19153 24905 19165 24908
rect 19199 24905 19211 24939
rect 19153 24899 19211 24905
rect 19518 24896 19524 24948
rect 19576 24936 19582 24948
rect 19889 24939 19947 24945
rect 19889 24936 19901 24939
rect 19576 24908 19901 24936
rect 19576 24896 19582 24908
rect 19889 24905 19901 24908
rect 19935 24905 19947 24939
rect 19889 24899 19947 24905
rect 20346 24896 20352 24948
rect 20404 24936 20410 24948
rect 21174 24936 21180 24948
rect 20404 24908 21180 24936
rect 20404 24896 20410 24908
rect 21174 24896 21180 24908
rect 21232 24896 21238 24948
rect 22002 24936 22008 24948
rect 21963 24908 22008 24936
rect 22002 24896 22008 24908
rect 22060 24896 22066 24948
rect 20257 24871 20315 24877
rect 20257 24868 20269 24871
rect 18656 24840 18828 24868
rect 19168 24840 20269 24868
rect 18656 24828 18662 24840
rect 18230 24760 18236 24812
rect 18288 24800 18294 24812
rect 19061 24803 19119 24809
rect 19061 24800 19073 24803
rect 18288 24772 19073 24800
rect 18288 24760 18294 24772
rect 19061 24769 19073 24772
rect 19107 24800 19119 24803
rect 19168 24800 19196 24840
rect 20257 24837 20269 24840
rect 20303 24868 20315 24871
rect 22462 24868 22468 24880
rect 20303 24840 21956 24868
rect 22423 24840 22468 24868
rect 20303 24837 20315 24840
rect 20257 24831 20315 24837
rect 19107 24772 19196 24800
rect 19107 24769 19119 24772
rect 19061 24763 19119 24769
rect 20070 24760 20076 24812
rect 20128 24798 20134 24812
rect 20180 24798 20392 24800
rect 20128 24772 20392 24798
rect 20128 24770 20208 24772
rect 20128 24760 20134 24770
rect 19242 24732 19248 24744
rect 19203 24704 19248 24732
rect 19242 24692 19248 24704
rect 19300 24692 19306 24744
rect 20364 24741 20392 24772
rect 21174 24760 21180 24812
rect 21232 24800 21238 24812
rect 21269 24803 21327 24809
rect 21269 24800 21281 24803
rect 21232 24772 21281 24800
rect 21232 24760 21238 24772
rect 21269 24769 21281 24772
rect 21315 24769 21327 24803
rect 21928 24800 21956 24840
rect 22462 24828 22468 24840
rect 22520 24828 22526 24880
rect 23198 24828 23204 24880
rect 23256 24868 23262 24880
rect 23256 24840 23612 24868
rect 23256 24828 23262 24840
rect 22370 24800 22376 24812
rect 21928 24772 22376 24800
rect 21269 24763 21327 24769
rect 22370 24760 22376 24772
rect 22428 24760 22434 24812
rect 22554 24760 22560 24812
rect 22612 24800 22618 24812
rect 23584 24809 23612 24840
rect 27264 24840 27476 24868
rect 23293 24803 23351 24809
rect 23293 24800 23305 24803
rect 22612 24772 23305 24800
rect 22612 24760 22618 24772
rect 23293 24769 23305 24772
rect 23339 24769 23351 24803
rect 23293 24763 23351 24769
rect 23569 24803 23627 24809
rect 23569 24769 23581 24803
rect 23615 24800 23627 24803
rect 24394 24800 24400 24812
rect 23615 24772 24400 24800
rect 23615 24769 23627 24772
rect 23569 24763 23627 24769
rect 20349 24735 20407 24741
rect 19352 24704 19555 24732
rect 19352 24664 19380 24704
rect 17972 24636 19380 24664
rect 19527 24664 19555 24704
rect 20349 24701 20361 24735
rect 20395 24701 20407 24735
rect 20530 24732 20536 24744
rect 20491 24704 20536 24732
rect 20349 24695 20407 24701
rect 20530 24692 20536 24704
rect 20588 24692 20594 24744
rect 22649 24735 22707 24741
rect 22649 24701 22661 24735
rect 22695 24732 22707 24735
rect 23198 24732 23204 24744
rect 22695 24704 23204 24732
rect 22695 24701 22707 24704
rect 22649 24695 22707 24701
rect 23198 24692 23204 24704
rect 23256 24692 23262 24744
rect 23308 24732 23336 24763
rect 24394 24760 24400 24772
rect 24452 24800 24458 24812
rect 24581 24803 24639 24809
rect 24581 24800 24593 24803
rect 24452 24772 24593 24800
rect 24452 24760 24458 24772
rect 24581 24769 24593 24772
rect 24627 24769 24639 24803
rect 24762 24800 24768 24812
rect 24723 24772 24768 24800
rect 24581 24763 24639 24769
rect 24762 24760 24768 24772
rect 24820 24760 24826 24812
rect 24857 24803 24915 24809
rect 24857 24769 24869 24803
rect 24903 24769 24915 24803
rect 24857 24763 24915 24769
rect 23842 24732 23848 24744
rect 23308 24704 23848 24732
rect 23842 24692 23848 24704
rect 23900 24692 23906 24744
rect 24872 24732 24900 24763
rect 24946 24760 24952 24812
rect 25004 24800 25010 24812
rect 25777 24803 25835 24809
rect 25004 24772 25049 24800
rect 25004 24760 25010 24772
rect 25777 24769 25789 24803
rect 25823 24769 25835 24803
rect 25777 24763 25835 24769
rect 25038 24732 25044 24744
rect 24872 24704 25044 24732
rect 25038 24692 25044 24704
rect 25096 24692 25102 24744
rect 25792 24732 25820 24763
rect 26234 24760 26240 24812
rect 26292 24800 26298 24812
rect 26421 24803 26479 24809
rect 26421 24800 26433 24803
rect 26292 24772 26433 24800
rect 26292 24760 26298 24772
rect 26421 24769 26433 24772
rect 26467 24769 26479 24803
rect 26421 24763 26479 24769
rect 27264 24732 27292 24840
rect 27341 24803 27399 24809
rect 27341 24769 27353 24803
rect 27387 24769 27399 24803
rect 27448 24800 27476 24840
rect 27982 24800 27988 24812
rect 27448 24772 27988 24800
rect 27341 24763 27399 24769
rect 25792 24704 27292 24732
rect 19527 24636 21220 24664
rect 19426 24596 19432 24608
rect 17144 24568 19432 24596
rect 19426 24556 19432 24568
rect 19484 24556 19490 24608
rect 21082 24596 21088 24608
rect 21043 24568 21088 24596
rect 21082 24556 21088 24568
rect 21140 24556 21146 24608
rect 21192 24596 21220 24636
rect 21266 24624 21272 24676
rect 21324 24664 21330 24676
rect 27356 24664 27384 24763
rect 27982 24760 27988 24772
rect 28040 24760 28046 24812
rect 21324 24636 27384 24664
rect 21324 24624 21330 24636
rect 24946 24596 24952 24608
rect 21192 24568 24952 24596
rect 24946 24556 24952 24568
rect 25004 24556 25010 24608
rect 25133 24599 25191 24605
rect 25133 24565 25145 24599
rect 25179 24596 25191 24599
rect 25314 24596 25320 24608
rect 25179 24568 25320 24596
rect 25179 24565 25191 24568
rect 25133 24559 25191 24565
rect 25314 24556 25320 24568
rect 25372 24556 25378 24608
rect 25590 24596 25596 24608
rect 25551 24568 25596 24596
rect 25590 24556 25596 24568
rect 25648 24556 25654 24608
rect 26237 24599 26295 24605
rect 26237 24565 26249 24599
rect 26283 24596 26295 24599
rect 27062 24596 27068 24608
rect 26283 24568 27068 24596
rect 26283 24565 26295 24568
rect 26237 24559 26295 24565
rect 27062 24556 27068 24568
rect 27120 24556 27126 24608
rect 27157 24599 27215 24605
rect 27157 24565 27169 24599
rect 27203 24596 27215 24599
rect 27522 24596 27528 24608
rect 27203 24568 27528 24596
rect 27203 24565 27215 24568
rect 27157 24559 27215 24565
rect 27522 24556 27528 24568
rect 27580 24556 27586 24608
rect 1104 24506 28060 24528
rect 1104 24454 5442 24506
rect 5494 24454 5506 24506
rect 5558 24454 5570 24506
rect 5622 24454 5634 24506
rect 5686 24454 5698 24506
rect 5750 24454 14428 24506
rect 14480 24454 14492 24506
rect 14544 24454 14556 24506
rect 14608 24454 14620 24506
rect 14672 24454 14684 24506
rect 14736 24454 23413 24506
rect 23465 24454 23477 24506
rect 23529 24454 23541 24506
rect 23593 24454 23605 24506
rect 23657 24454 23669 24506
rect 23721 24454 28060 24506
rect 1104 24432 28060 24454
rect 198 24352 204 24404
rect 256 24392 262 24404
rect 3234 24392 3240 24404
rect 256 24364 3240 24392
rect 256 24352 262 24364
rect 3234 24352 3240 24364
rect 3292 24352 3298 24404
rect 3510 24352 3516 24404
rect 3568 24392 3574 24404
rect 3789 24395 3847 24401
rect 3789 24392 3801 24395
rect 3568 24364 3801 24392
rect 3568 24352 3574 24364
rect 3789 24361 3801 24364
rect 3835 24361 3847 24395
rect 3789 24355 3847 24361
rect 4709 24395 4767 24401
rect 4709 24361 4721 24395
rect 4755 24392 4767 24395
rect 5258 24392 5264 24404
rect 4755 24364 5264 24392
rect 4755 24361 4767 24364
rect 4709 24355 4767 24361
rect 5258 24352 5264 24364
rect 5316 24352 5322 24404
rect 5902 24392 5908 24404
rect 5863 24364 5908 24392
rect 5902 24352 5908 24364
rect 5960 24352 5966 24404
rect 7561 24395 7619 24401
rect 7561 24361 7573 24395
rect 7607 24392 7619 24395
rect 7742 24392 7748 24404
rect 7607 24364 7748 24392
rect 7607 24361 7619 24364
rect 7561 24355 7619 24361
rect 7742 24352 7748 24364
rect 7800 24352 7806 24404
rect 8294 24352 8300 24404
rect 8352 24392 8358 24404
rect 9033 24395 9091 24401
rect 9033 24392 9045 24395
rect 8352 24364 9045 24392
rect 8352 24352 8358 24364
rect 9033 24361 9045 24364
rect 9079 24361 9091 24395
rect 9033 24355 9091 24361
rect 9861 24395 9919 24401
rect 9861 24361 9873 24395
rect 9907 24392 9919 24395
rect 10778 24392 10784 24404
rect 9907 24364 10784 24392
rect 9907 24361 9919 24364
rect 9861 24355 9919 24361
rect 10778 24352 10784 24364
rect 10836 24352 10842 24404
rect 12526 24352 12532 24404
rect 12584 24392 12590 24404
rect 12621 24395 12679 24401
rect 12621 24392 12633 24395
rect 12584 24364 12633 24392
rect 12584 24352 12590 24364
rect 12621 24361 12633 24364
rect 12667 24361 12679 24395
rect 14826 24392 14832 24404
rect 14787 24364 14832 24392
rect 12621 24355 12679 24361
rect 14826 24352 14832 24364
rect 14884 24352 14890 24404
rect 17218 24352 17224 24404
rect 17276 24352 17282 24404
rect 17770 24352 17776 24404
rect 17828 24392 17834 24404
rect 17865 24395 17923 24401
rect 17865 24392 17877 24395
rect 17828 24364 17877 24392
rect 17828 24352 17834 24364
rect 17865 24361 17877 24364
rect 17911 24361 17923 24395
rect 17865 24355 17923 24361
rect 18782 24352 18788 24404
rect 18840 24392 18846 24404
rect 19245 24395 19303 24401
rect 19245 24392 19257 24395
rect 18840 24364 19257 24392
rect 18840 24352 18846 24364
rect 19245 24361 19257 24364
rect 19291 24361 19303 24395
rect 19245 24355 19303 24361
rect 19426 24352 19432 24404
rect 19484 24392 19490 24404
rect 20714 24392 20720 24404
rect 19484 24364 20720 24392
rect 19484 24352 19490 24364
rect 20714 24352 20720 24364
rect 20772 24352 20778 24404
rect 21085 24395 21143 24401
rect 21085 24361 21097 24395
rect 21131 24392 21143 24395
rect 21910 24392 21916 24404
rect 21131 24364 21916 24392
rect 21131 24361 21143 24364
rect 21085 24355 21143 24361
rect 21910 24352 21916 24364
rect 21968 24352 21974 24404
rect 22554 24352 22560 24404
rect 22612 24352 22618 24404
rect 22738 24352 22744 24404
rect 22796 24392 22802 24404
rect 23017 24395 23075 24401
rect 22796 24364 22968 24392
rect 22796 24352 22802 24364
rect 2958 24284 2964 24336
rect 3016 24324 3022 24336
rect 4522 24324 4528 24336
rect 3016 24296 4528 24324
rect 3016 24284 3022 24296
rect 4522 24284 4528 24296
rect 4580 24284 4586 24336
rect 5810 24284 5816 24336
rect 5868 24324 5874 24336
rect 6178 24324 6184 24336
rect 5868 24296 6184 24324
rect 5868 24284 5874 24296
rect 6178 24284 6184 24296
rect 6236 24284 6242 24336
rect 7650 24284 7656 24336
rect 7708 24324 7714 24336
rect 10321 24327 10379 24333
rect 10321 24324 10333 24327
rect 7708 24296 10333 24324
rect 7708 24284 7714 24296
rect 10321 24293 10333 24296
rect 10367 24293 10379 24327
rect 10321 24287 10379 24293
rect 16209 24327 16267 24333
rect 16209 24293 16221 24327
rect 16255 24324 16267 24327
rect 16850 24324 16856 24336
rect 16255 24296 16856 24324
rect 16255 24293 16267 24296
rect 16209 24287 16267 24293
rect 16850 24284 16856 24296
rect 16908 24284 16914 24336
rect 17236 24324 17264 24352
rect 17678 24324 17684 24336
rect 17236 24296 17684 24324
rect 17678 24284 17684 24296
rect 17736 24324 17742 24336
rect 22572 24324 22600 24352
rect 17736 24296 22600 24324
rect 22940 24324 22968 24364
rect 23017 24361 23029 24395
rect 23063 24392 23075 24395
rect 23290 24392 23296 24404
rect 23063 24364 23296 24392
rect 23063 24361 23075 24364
rect 23017 24355 23075 24361
rect 23290 24352 23296 24364
rect 23348 24352 23354 24404
rect 25498 24392 25504 24404
rect 25459 24364 25504 24392
rect 25498 24352 25504 24364
rect 25556 24352 25562 24404
rect 25958 24352 25964 24404
rect 26016 24392 26022 24404
rect 27154 24392 27160 24404
rect 26016 24364 27160 24392
rect 26016 24352 26022 24364
rect 27154 24352 27160 24364
rect 27212 24352 27218 24404
rect 23382 24324 23388 24336
rect 22940 24296 23388 24324
rect 17736 24284 17742 24296
rect 23382 24284 23388 24296
rect 23440 24284 23446 24336
rect 1394 24256 1400 24268
rect 1355 24228 1400 24256
rect 1394 24216 1400 24228
rect 1452 24216 1458 24268
rect 3142 24216 3148 24268
rect 3200 24256 3206 24268
rect 4706 24256 4712 24268
rect 3200 24228 4712 24256
rect 3200 24216 3206 24228
rect 4706 24216 4712 24228
rect 4764 24216 4770 24268
rect 5350 24256 5356 24268
rect 5311 24228 5356 24256
rect 5350 24216 5356 24228
rect 5408 24216 5414 24268
rect 6549 24259 6607 24265
rect 6549 24225 6561 24259
rect 6595 24256 6607 24259
rect 6914 24256 6920 24268
rect 6595 24228 6920 24256
rect 6595 24225 6607 24228
rect 6549 24219 6607 24225
rect 6914 24216 6920 24228
rect 6972 24216 6978 24268
rect 7745 24259 7803 24265
rect 7745 24225 7757 24259
rect 7791 24256 7803 24259
rect 8110 24256 8116 24268
rect 7791 24228 8116 24256
rect 7791 24225 7803 24228
rect 7745 24219 7803 24225
rect 8110 24216 8116 24228
rect 8168 24216 8174 24268
rect 8478 24216 8484 24268
rect 8536 24256 8542 24268
rect 9858 24256 9864 24268
rect 8536 24228 9864 24256
rect 8536 24216 8542 24228
rect 9858 24216 9864 24228
rect 9916 24216 9922 24268
rect 10873 24259 10931 24265
rect 10873 24225 10885 24259
rect 10919 24256 10931 24259
rect 10962 24256 10968 24268
rect 10919 24228 10968 24256
rect 10919 24225 10931 24228
rect 10873 24219 10931 24225
rect 10962 24216 10968 24228
rect 11020 24216 11026 24268
rect 15838 24256 15844 24268
rect 15799 24228 15844 24256
rect 15838 24216 15844 24228
rect 15896 24216 15902 24268
rect 16301 24259 16359 24265
rect 16301 24225 16313 24259
rect 16347 24256 16359 24259
rect 17218 24256 17224 24268
rect 16347 24228 17224 24256
rect 16347 24225 16359 24228
rect 16301 24219 16359 24225
rect 17218 24216 17224 24228
rect 17276 24216 17282 24268
rect 18509 24259 18567 24265
rect 17926 24228 18368 24256
rect 3786 24188 3792 24200
rect 3747 24160 3792 24188
rect 3786 24148 3792 24160
rect 3844 24148 3850 24200
rect 3970 24148 3976 24200
rect 4028 24188 4034 24200
rect 6362 24188 6368 24200
rect 4028 24160 6368 24188
rect 4028 24148 4034 24160
rect 6362 24148 6368 24160
rect 6420 24148 6426 24200
rect 7837 24191 7895 24197
rect 7837 24157 7849 24191
rect 7883 24188 7895 24191
rect 7926 24188 7932 24200
rect 7883 24160 7932 24188
rect 7883 24157 7895 24160
rect 7837 24151 7895 24157
rect 7926 24148 7932 24160
rect 7984 24148 7990 24200
rect 8018 24148 8024 24200
rect 8076 24188 8082 24200
rect 8205 24191 8263 24197
rect 8205 24188 8217 24191
rect 8076 24160 8217 24188
rect 8076 24148 8082 24160
rect 8205 24157 8217 24160
rect 8251 24188 8263 24191
rect 8941 24191 8999 24197
rect 8941 24188 8953 24191
rect 8251 24160 8953 24188
rect 8251 24157 8263 24160
rect 8205 24151 8263 24157
rect 1664 24123 1722 24129
rect 1664 24089 1676 24123
rect 1710 24120 1722 24123
rect 3234 24120 3240 24132
rect 1710 24092 3240 24120
rect 1710 24089 1722 24092
rect 1664 24083 1722 24089
rect 3234 24080 3240 24092
rect 3292 24080 3298 24132
rect 4614 24080 4620 24132
rect 4672 24120 4678 24132
rect 5074 24120 5080 24132
rect 4672 24092 5080 24120
rect 4672 24080 4678 24092
rect 5074 24080 5080 24092
rect 5132 24080 5138 24132
rect 6273 24123 6331 24129
rect 6273 24089 6285 24123
rect 6319 24120 6331 24123
rect 6638 24120 6644 24132
rect 6319 24092 6644 24120
rect 6319 24089 6331 24092
rect 6273 24083 6331 24089
rect 6638 24080 6644 24092
rect 6696 24080 6702 24132
rect 2777 24055 2835 24061
rect 2777 24021 2789 24055
rect 2823 24052 2835 24055
rect 2958 24052 2964 24064
rect 2823 24024 2964 24052
rect 2823 24021 2835 24024
rect 2777 24015 2835 24021
rect 2958 24012 2964 24024
rect 3016 24052 3022 24064
rect 4062 24052 4068 24064
rect 3016 24024 4068 24052
rect 3016 24012 3022 24024
rect 4062 24012 4068 24024
rect 4120 24012 4126 24064
rect 4157 24055 4215 24061
rect 4157 24021 4169 24055
rect 4203 24052 4215 24055
rect 4246 24052 4252 24064
rect 4203 24024 4252 24052
rect 4203 24021 4215 24024
rect 4157 24015 4215 24021
rect 4246 24012 4252 24024
rect 4304 24012 4310 24064
rect 5169 24055 5227 24061
rect 5169 24021 5181 24055
rect 5215 24052 5227 24055
rect 5902 24052 5908 24064
rect 5215 24024 5908 24052
rect 5215 24021 5227 24024
rect 5169 24015 5227 24021
rect 5902 24012 5908 24024
rect 5960 24012 5966 24064
rect 6362 24012 6368 24064
rect 6420 24052 6426 24064
rect 6420 24024 6465 24052
rect 6420 24012 6426 24024
rect 7834 24012 7840 24064
rect 7892 24052 7898 24064
rect 7929 24055 7987 24061
rect 7929 24052 7941 24055
rect 7892 24024 7941 24052
rect 7892 24012 7898 24024
rect 7929 24021 7941 24024
rect 7975 24021 7987 24055
rect 7929 24015 7987 24021
rect 8113 24055 8171 24061
rect 8113 24021 8125 24055
rect 8159 24052 8171 24055
rect 8294 24052 8300 24064
rect 8159 24024 8300 24052
rect 8159 24021 8171 24024
rect 8113 24015 8171 24021
rect 8294 24012 8300 24024
rect 8352 24012 8358 24064
rect 8864 24052 8892 24160
rect 8941 24157 8953 24160
rect 8987 24157 8999 24191
rect 8941 24151 8999 24157
rect 9030 24148 9036 24200
rect 9088 24188 9094 24200
rect 9125 24191 9183 24197
rect 9125 24188 9137 24191
rect 9088 24160 9137 24188
rect 9088 24148 9094 24160
rect 9125 24157 9137 24160
rect 9171 24157 9183 24191
rect 9950 24188 9956 24200
rect 9125 24151 9183 24157
rect 9232 24160 9956 24188
rect 9232 24052 9260 24160
rect 9950 24148 9956 24160
rect 10008 24148 10014 24200
rect 10045 24191 10103 24197
rect 10045 24157 10057 24191
rect 10091 24157 10103 24191
rect 10045 24151 10103 24157
rect 10061 24120 10089 24151
rect 10134 24148 10140 24200
rect 10192 24188 10198 24200
rect 10410 24188 10416 24200
rect 10192 24160 10237 24188
rect 10371 24160 10416 24188
rect 10192 24148 10198 24160
rect 10410 24148 10416 24160
rect 10468 24148 10474 24200
rect 11146 24188 11152 24200
rect 11059 24160 11152 24188
rect 11146 24148 11152 24160
rect 11204 24188 11210 24200
rect 11698 24188 11704 24200
rect 11204 24160 11704 24188
rect 11204 24148 11210 24160
rect 11698 24148 11704 24160
rect 11756 24148 11762 24200
rect 13170 24188 13176 24200
rect 12406 24160 13032 24188
rect 13131 24160 13176 24188
rect 11606 24120 11612 24132
rect 10061 24092 11612 24120
rect 11606 24080 11612 24092
rect 11664 24080 11670 24132
rect 8864 24024 9260 24052
rect 9582 24012 9588 24064
rect 9640 24052 9646 24064
rect 12406 24052 12434 24160
rect 12529 24123 12587 24129
rect 12529 24089 12541 24123
rect 12575 24120 12587 24123
rect 12618 24120 12624 24132
rect 12575 24092 12624 24120
rect 12575 24089 12587 24092
rect 12529 24083 12587 24089
rect 12618 24080 12624 24092
rect 12676 24080 12682 24132
rect 13004 24120 13032 24160
rect 13170 24148 13176 24160
rect 13228 24148 13234 24200
rect 14182 24148 14188 24200
rect 14240 24188 14246 24200
rect 14369 24191 14427 24197
rect 14369 24188 14381 24191
rect 14240 24160 14381 24188
rect 14240 24148 14246 24160
rect 14369 24157 14381 24160
rect 14415 24157 14427 24191
rect 14734 24188 14740 24200
rect 14695 24160 14740 24188
rect 14369 24151 14427 24157
rect 14734 24148 14740 24160
rect 14792 24148 14798 24200
rect 15194 24148 15200 24200
rect 15252 24188 15258 24200
rect 16666 24188 16672 24200
rect 15252 24160 16672 24188
rect 15252 24148 15258 24160
rect 16666 24148 16672 24160
rect 16724 24188 16730 24200
rect 16761 24191 16819 24197
rect 16761 24188 16773 24191
rect 16724 24160 16773 24188
rect 16724 24148 16730 24160
rect 16761 24157 16773 24160
rect 16807 24157 16819 24191
rect 16761 24151 16819 24157
rect 16942 24148 16948 24200
rect 17000 24188 17006 24200
rect 17037 24191 17095 24197
rect 17037 24188 17049 24191
rect 17000 24160 17049 24188
rect 17000 24148 17006 24160
rect 17037 24157 17049 24160
rect 17083 24157 17095 24191
rect 17926 24188 17954 24228
rect 18230 24188 18236 24200
rect 17037 24151 17095 24157
rect 17144 24160 17954 24188
rect 18191 24160 18236 24188
rect 13004 24092 14596 24120
rect 13262 24052 13268 24064
rect 9640 24024 12434 24052
rect 13223 24024 13268 24052
rect 9640 24012 9646 24024
rect 13262 24012 13268 24024
rect 13320 24012 13326 24064
rect 14568 24061 14596 24092
rect 15930 24080 15936 24132
rect 15988 24120 15994 24132
rect 17144 24120 17172 24160
rect 18230 24148 18236 24160
rect 18288 24148 18294 24200
rect 18340 24188 18368 24228
rect 18509 24225 18521 24259
rect 18555 24256 18567 24259
rect 19610 24256 19616 24268
rect 18555 24228 19616 24256
rect 18555 24225 18567 24228
rect 18509 24219 18567 24225
rect 19610 24216 19616 24228
rect 19668 24216 19674 24268
rect 19794 24256 19800 24268
rect 19755 24228 19800 24256
rect 19794 24216 19800 24228
rect 19852 24216 19858 24268
rect 20162 24216 20168 24268
rect 20220 24256 20226 24268
rect 21634 24256 21640 24268
rect 20220 24228 20944 24256
rect 21595 24228 21640 24256
rect 20220 24216 20226 24228
rect 19518 24188 19524 24200
rect 18340 24160 19524 24188
rect 19518 24148 19524 24160
rect 19576 24148 19582 24200
rect 19705 24191 19763 24197
rect 19705 24157 19717 24191
rect 19751 24188 19763 24191
rect 20180 24188 20208 24216
rect 19751 24160 20208 24188
rect 19751 24157 19763 24160
rect 19705 24151 19763 24157
rect 20438 24148 20444 24200
rect 20496 24188 20502 24200
rect 20625 24191 20683 24197
rect 20625 24188 20637 24191
rect 20496 24160 20637 24188
rect 20496 24148 20502 24160
rect 20625 24157 20637 24160
rect 20671 24157 20683 24191
rect 20916 24188 20944 24228
rect 21634 24216 21640 24228
rect 21692 24216 21698 24268
rect 22554 24256 22560 24268
rect 21744 24228 22560 24256
rect 21545 24191 21603 24197
rect 21545 24188 21557 24191
rect 20916 24160 21557 24188
rect 20625 24151 20683 24157
rect 21545 24157 21557 24160
rect 21591 24188 21603 24191
rect 21744 24188 21772 24228
rect 22554 24216 22560 24228
rect 22612 24216 22618 24268
rect 22738 24216 22744 24268
rect 22796 24256 22802 24268
rect 23569 24259 23627 24265
rect 23569 24256 23581 24259
rect 22796 24228 23581 24256
rect 22796 24216 22802 24228
rect 23569 24225 23581 24228
rect 23615 24225 23627 24259
rect 23569 24219 23627 24225
rect 25406 24216 25412 24268
rect 25464 24256 25470 24268
rect 25958 24256 25964 24268
rect 25464 24228 25964 24256
rect 25464 24216 25470 24228
rect 25958 24216 25964 24228
rect 26016 24216 26022 24268
rect 21591 24160 21772 24188
rect 21591 24157 21603 24160
rect 21545 24151 21603 24157
rect 21910 24148 21916 24200
rect 21968 24188 21974 24200
rect 22465 24191 22523 24197
rect 22465 24188 22477 24191
rect 21968 24160 22477 24188
rect 21968 24148 21974 24160
rect 22465 24157 22477 24160
rect 22511 24157 22523 24191
rect 22465 24151 22523 24157
rect 24486 24148 24492 24200
rect 24544 24188 24550 24200
rect 24581 24191 24639 24197
rect 24581 24188 24593 24191
rect 24544 24160 24593 24188
rect 24544 24148 24550 24160
rect 24581 24157 24593 24160
rect 24627 24157 24639 24191
rect 24581 24151 24639 24157
rect 25133 24191 25191 24197
rect 25133 24157 25145 24191
rect 25179 24157 25191 24191
rect 25314 24188 25320 24200
rect 25275 24160 25320 24188
rect 25133 24151 25191 24157
rect 15988 24092 17172 24120
rect 15988 24080 15994 24092
rect 17494 24080 17500 24132
rect 17552 24120 17558 24132
rect 21266 24120 21272 24132
rect 17552 24092 21272 24120
rect 17552 24080 17558 24092
rect 21266 24080 21272 24092
rect 21324 24080 21330 24132
rect 21450 24120 21456 24132
rect 21411 24092 21456 24120
rect 21450 24080 21456 24092
rect 21508 24080 21514 24132
rect 21818 24080 21824 24132
rect 21876 24120 21882 24132
rect 22830 24120 22836 24132
rect 21876 24092 22836 24120
rect 21876 24080 21882 24092
rect 22830 24080 22836 24092
rect 22888 24080 22894 24132
rect 23477 24123 23535 24129
rect 23477 24089 23489 24123
rect 23523 24120 23535 24123
rect 24118 24120 24124 24132
rect 23523 24092 24124 24120
rect 23523 24089 23535 24092
rect 23477 24083 23535 24089
rect 24118 24080 24124 24092
rect 24176 24080 24182 24132
rect 25148 24120 25176 24151
rect 25314 24148 25320 24160
rect 25372 24148 25378 24200
rect 26228 24191 26286 24197
rect 26228 24157 26240 24191
rect 26274 24188 26286 24191
rect 26510 24188 26516 24200
rect 26274 24160 26516 24188
rect 26274 24157 26286 24160
rect 26228 24151 26286 24157
rect 26510 24148 26516 24160
rect 26568 24148 26574 24200
rect 26142 24120 26148 24132
rect 25148 24092 26148 24120
rect 26142 24080 26148 24092
rect 26200 24080 26206 24132
rect 14553 24055 14611 24061
rect 14553 24021 14565 24055
rect 14599 24052 14611 24055
rect 15102 24052 15108 24064
rect 14599 24024 15108 24052
rect 14599 24021 14611 24024
rect 14553 24015 14611 24021
rect 15102 24012 15108 24024
rect 15160 24012 15166 24064
rect 17313 24055 17371 24061
rect 17313 24021 17325 24055
rect 17359 24052 17371 24055
rect 18230 24052 18236 24064
rect 17359 24024 18236 24052
rect 17359 24021 17371 24024
rect 17313 24015 17371 24021
rect 18230 24012 18236 24024
rect 18288 24012 18294 24064
rect 18325 24055 18383 24061
rect 18325 24021 18337 24055
rect 18371 24052 18383 24055
rect 18414 24052 18420 24064
rect 18371 24024 18420 24052
rect 18371 24021 18383 24024
rect 18325 24015 18383 24021
rect 18414 24012 18420 24024
rect 18472 24012 18478 24064
rect 19334 24012 19340 24064
rect 19392 24052 19398 24064
rect 19613 24055 19671 24061
rect 19613 24052 19625 24055
rect 19392 24024 19625 24052
rect 19392 24012 19398 24024
rect 19613 24021 19625 24024
rect 19659 24021 19671 24055
rect 19613 24015 19671 24021
rect 20254 24012 20260 24064
rect 20312 24052 20318 24064
rect 20441 24055 20499 24061
rect 20441 24052 20453 24055
rect 20312 24024 20453 24052
rect 20312 24012 20318 24024
rect 20441 24021 20453 24024
rect 20487 24021 20499 24055
rect 20441 24015 20499 24021
rect 20714 24012 20720 24064
rect 20772 24052 20778 24064
rect 21910 24052 21916 24064
rect 20772 24024 21916 24052
rect 20772 24012 20778 24024
rect 21910 24012 21916 24024
rect 21968 24012 21974 24064
rect 22278 24052 22284 24064
rect 22239 24024 22284 24052
rect 22278 24012 22284 24024
rect 22336 24012 22342 24064
rect 22370 24012 22376 24064
rect 22428 24052 22434 24064
rect 23382 24052 23388 24064
rect 22428 24024 23388 24052
rect 22428 24012 22434 24024
rect 23382 24012 23388 24024
rect 23440 24012 23446 24064
rect 24026 24012 24032 24064
rect 24084 24052 24090 24064
rect 24397 24055 24455 24061
rect 24397 24052 24409 24055
rect 24084 24024 24409 24052
rect 24084 24012 24090 24024
rect 24397 24021 24409 24024
rect 24443 24021 24455 24055
rect 24397 24015 24455 24021
rect 25038 24012 25044 24064
rect 25096 24052 25102 24064
rect 25498 24052 25504 24064
rect 25096 24024 25504 24052
rect 25096 24012 25102 24024
rect 25498 24012 25504 24024
rect 25556 24052 25562 24064
rect 27341 24055 27399 24061
rect 27341 24052 27353 24055
rect 25556 24024 27353 24052
rect 25556 24012 25562 24024
rect 27341 24021 27353 24024
rect 27387 24021 27399 24055
rect 27341 24015 27399 24021
rect 1104 23962 28060 23984
rect 1104 23910 9935 23962
rect 9987 23910 9999 23962
rect 10051 23910 10063 23962
rect 10115 23910 10127 23962
rect 10179 23910 10191 23962
rect 10243 23910 18920 23962
rect 18972 23910 18984 23962
rect 19036 23910 19048 23962
rect 19100 23910 19112 23962
rect 19164 23910 19176 23962
rect 19228 23910 28060 23962
rect 1104 23888 28060 23910
rect 1949 23851 2007 23857
rect 1949 23817 1961 23851
rect 1995 23817 2007 23851
rect 1949 23811 2007 23817
rect 3513 23851 3571 23857
rect 3513 23817 3525 23851
rect 3559 23848 3571 23851
rect 4246 23848 4252 23860
rect 3559 23820 4252 23848
rect 3559 23817 3571 23820
rect 3513 23811 3571 23817
rect 1964 23780 1992 23811
rect 4246 23808 4252 23820
rect 4304 23808 4310 23860
rect 5350 23808 5356 23860
rect 5408 23848 5414 23860
rect 5721 23851 5779 23857
rect 5721 23848 5733 23851
rect 5408 23820 5733 23848
rect 5408 23808 5414 23820
rect 5721 23817 5733 23820
rect 5767 23817 5779 23851
rect 5721 23811 5779 23817
rect 4525 23783 4583 23789
rect 4525 23780 4537 23783
rect 1964 23752 3740 23780
rect 1673 23715 1731 23721
rect 1673 23681 1685 23715
rect 1719 23712 1731 23715
rect 2130 23712 2136 23724
rect 1719 23684 2136 23712
rect 1719 23681 1731 23684
rect 1673 23675 1731 23681
rect 2130 23672 2136 23684
rect 2188 23672 2194 23724
rect 3418 23712 3424 23724
rect 3379 23684 3424 23712
rect 3418 23672 3424 23684
rect 3476 23672 3482 23724
rect 3602 23644 3608 23656
rect 3563 23616 3608 23644
rect 3602 23604 3608 23616
rect 3660 23604 3666 23656
rect 3712 23644 3740 23752
rect 3804 23752 4537 23780
rect 3804 23721 3832 23752
rect 4525 23749 4537 23752
rect 4571 23749 4583 23783
rect 5736 23780 5764 23811
rect 6086 23808 6092 23860
rect 6144 23848 6150 23860
rect 6365 23851 6423 23857
rect 6365 23848 6377 23851
rect 6144 23820 6377 23848
rect 6144 23808 6150 23820
rect 6365 23817 6377 23820
rect 6411 23817 6423 23851
rect 6365 23811 6423 23817
rect 6733 23851 6791 23857
rect 6733 23817 6745 23851
rect 6779 23848 6791 23851
rect 7006 23848 7012 23860
rect 6779 23820 7012 23848
rect 6779 23817 6791 23820
rect 6733 23811 6791 23817
rect 7006 23808 7012 23820
rect 7064 23808 7070 23860
rect 7561 23851 7619 23857
rect 7561 23817 7573 23851
rect 7607 23848 7619 23851
rect 7650 23848 7656 23860
rect 7607 23820 7656 23848
rect 7607 23817 7619 23820
rect 7561 23811 7619 23817
rect 7650 23808 7656 23820
rect 7708 23808 7714 23860
rect 7834 23808 7840 23860
rect 7892 23848 7898 23860
rect 7929 23851 7987 23857
rect 7929 23848 7941 23851
rect 7892 23820 7941 23848
rect 7892 23808 7898 23820
rect 7929 23817 7941 23820
rect 7975 23817 7987 23851
rect 7929 23811 7987 23817
rect 8938 23808 8944 23860
rect 8996 23848 9002 23860
rect 9214 23848 9220 23860
rect 8996 23820 9220 23848
rect 8996 23808 9002 23820
rect 9214 23808 9220 23820
rect 9272 23848 9278 23860
rect 9272 23820 11560 23848
rect 9272 23808 9278 23820
rect 8113 23783 8171 23789
rect 5736 23752 7420 23780
rect 4525 23743 4583 23749
rect 3789 23715 3847 23721
rect 3789 23681 3801 23715
rect 3835 23681 3847 23715
rect 3789 23675 3847 23681
rect 4062 23672 4068 23724
rect 4120 23712 4126 23724
rect 4249 23715 4307 23721
rect 4249 23712 4261 23715
rect 4120 23684 4261 23712
rect 4120 23672 4126 23684
rect 4249 23681 4261 23684
rect 4295 23681 4307 23715
rect 5258 23712 5264 23724
rect 4249 23675 4307 23681
rect 4356 23684 5264 23712
rect 4356 23644 4384 23684
rect 5258 23672 5264 23684
rect 5316 23672 5322 23724
rect 5629 23715 5687 23721
rect 5629 23681 5641 23715
rect 5675 23681 5687 23715
rect 5629 23675 5687 23681
rect 6825 23715 6883 23721
rect 6825 23681 6837 23715
rect 6871 23712 6883 23715
rect 7282 23712 7288 23724
rect 6871 23684 7288 23712
rect 6871 23681 6883 23684
rect 6825 23675 6883 23681
rect 3712 23616 4384 23644
rect 4525 23647 4583 23653
rect 4525 23613 4537 23647
rect 4571 23613 4583 23647
rect 4525 23607 4583 23613
rect 3234 23536 3240 23588
rect 3292 23576 3298 23588
rect 3789 23579 3847 23585
rect 3789 23576 3801 23579
rect 3292 23548 3801 23576
rect 3292 23536 3298 23548
rect 3789 23545 3801 23548
rect 3835 23545 3847 23579
rect 3789 23539 3847 23545
rect 2774 23468 2780 23520
rect 2832 23508 2838 23520
rect 2832 23480 2877 23508
rect 2832 23468 2838 23480
rect 3602 23468 3608 23520
rect 3660 23508 3666 23520
rect 4341 23511 4399 23517
rect 4341 23508 4353 23511
rect 3660 23480 4353 23508
rect 3660 23468 3666 23480
rect 4341 23477 4353 23480
rect 4387 23508 4399 23511
rect 4430 23508 4436 23520
rect 4387 23480 4436 23508
rect 4387 23477 4399 23480
rect 4341 23471 4399 23477
rect 4430 23468 4436 23480
rect 4488 23468 4494 23520
rect 4540 23508 4568 23607
rect 5350 23604 5356 23656
rect 5408 23644 5414 23656
rect 5644 23644 5672 23675
rect 7282 23672 7288 23684
rect 7340 23672 7346 23724
rect 7392 23712 7420 23752
rect 8113 23749 8125 23783
rect 8159 23780 8171 23783
rect 8202 23780 8208 23792
rect 8159 23752 8208 23780
rect 8159 23749 8171 23752
rect 8113 23743 8171 23749
rect 8202 23740 8208 23752
rect 8260 23740 8266 23792
rect 8386 23740 8392 23792
rect 8444 23780 8450 23792
rect 9030 23780 9036 23792
rect 8444 23752 9036 23780
rect 8444 23740 8450 23752
rect 9030 23740 9036 23752
rect 9088 23740 9094 23792
rect 9122 23740 9128 23792
rect 9180 23780 9186 23792
rect 9180 23752 9628 23780
rect 9180 23740 9186 23752
rect 9600 23724 9628 23752
rect 7558 23712 7564 23724
rect 7392 23684 7564 23712
rect 7558 23672 7564 23684
rect 7616 23712 7622 23724
rect 8849 23715 8907 23721
rect 7616 23684 8248 23712
rect 7616 23672 7622 23684
rect 6914 23644 6920 23656
rect 5408 23616 6920 23644
rect 5408 23604 5414 23616
rect 6914 23604 6920 23616
rect 6972 23604 6978 23656
rect 7009 23647 7067 23653
rect 7009 23613 7021 23647
rect 7055 23644 7067 23647
rect 7650 23644 7656 23656
rect 7055 23616 7656 23644
rect 7055 23613 7067 23616
rect 7009 23607 7067 23613
rect 7650 23604 7656 23616
rect 7708 23604 7714 23656
rect 7745 23647 7803 23653
rect 7745 23613 7757 23647
rect 7791 23613 7803 23647
rect 7745 23607 7803 23613
rect 7837 23647 7895 23653
rect 7837 23613 7849 23647
rect 7883 23644 7895 23647
rect 7926 23644 7932 23656
rect 7883 23616 7932 23644
rect 7883 23613 7895 23616
rect 7837 23607 7895 23613
rect 7760 23576 7788 23607
rect 7926 23604 7932 23616
rect 7984 23604 7990 23656
rect 8220 23653 8248 23684
rect 8849 23681 8861 23715
rect 8895 23712 8907 23715
rect 9582 23712 9588 23724
rect 8895 23684 9352 23712
rect 9543 23684 9588 23712
rect 8895 23681 8907 23684
rect 8849 23675 8907 23681
rect 9324 23656 9352 23684
rect 9582 23672 9588 23684
rect 9640 23672 9646 23724
rect 9876 23721 9904 23820
rect 10410 23780 10416 23792
rect 10152 23752 10416 23780
rect 10152 23721 10180 23752
rect 10410 23740 10416 23752
rect 10468 23780 10474 23792
rect 11146 23780 11152 23792
rect 10468 23752 11152 23780
rect 10468 23740 10474 23752
rect 11146 23740 11152 23752
rect 11204 23740 11210 23792
rect 11532 23780 11560 23820
rect 11606 23808 11612 23860
rect 11664 23848 11670 23860
rect 11793 23851 11851 23857
rect 11793 23848 11805 23851
rect 11664 23820 11805 23848
rect 11664 23808 11670 23820
rect 11793 23817 11805 23820
rect 11839 23817 11851 23851
rect 13722 23848 13728 23860
rect 11793 23811 11851 23817
rect 12406 23820 13728 23848
rect 11532 23752 11652 23780
rect 9769 23715 9827 23721
rect 9769 23681 9781 23715
rect 9815 23681 9827 23715
rect 9769 23675 9827 23681
rect 9861 23715 9919 23721
rect 9861 23681 9873 23715
rect 9907 23681 9919 23715
rect 9861 23675 9919 23681
rect 10137 23715 10195 23721
rect 10137 23681 10149 23715
rect 10183 23681 10195 23715
rect 10778 23712 10784 23724
rect 10739 23684 10784 23712
rect 10137 23675 10195 23681
rect 8205 23647 8263 23653
rect 8205 23613 8217 23647
rect 8251 23613 8263 23647
rect 8938 23644 8944 23656
rect 8899 23616 8944 23644
rect 8205 23607 8263 23613
rect 8938 23604 8944 23616
rect 8996 23604 9002 23656
rect 9122 23644 9128 23656
rect 9083 23616 9128 23644
rect 9122 23604 9128 23616
rect 9180 23604 9186 23656
rect 9306 23604 9312 23656
rect 9364 23644 9370 23656
rect 9784 23644 9812 23675
rect 10778 23672 10784 23684
rect 10836 23672 10842 23724
rect 11517 23715 11575 23721
rect 11517 23681 11529 23715
rect 11563 23681 11575 23715
rect 11624 23712 11652 23752
rect 12406 23712 12434 23820
rect 13722 23808 13728 23820
rect 13780 23808 13786 23860
rect 15654 23808 15660 23860
rect 15712 23857 15718 23860
rect 15712 23851 15731 23857
rect 15719 23848 15731 23851
rect 17862 23848 17868 23860
rect 15719 23820 17868 23848
rect 15719 23817 15731 23820
rect 15712 23811 15731 23817
rect 15712 23808 15718 23811
rect 17862 23808 17868 23820
rect 17920 23808 17926 23860
rect 18969 23851 19027 23857
rect 18969 23817 18981 23851
rect 19015 23848 19027 23851
rect 19242 23848 19248 23860
rect 19015 23820 19248 23848
rect 19015 23817 19027 23820
rect 18969 23811 19027 23817
rect 19242 23808 19248 23820
rect 19300 23808 19306 23860
rect 20530 23808 20536 23860
rect 20588 23848 20594 23860
rect 22281 23851 22339 23857
rect 22281 23848 22293 23851
rect 20588 23820 22293 23848
rect 20588 23808 20594 23820
rect 22281 23817 22293 23820
rect 22327 23817 22339 23851
rect 22281 23811 22339 23817
rect 22554 23808 22560 23860
rect 22612 23848 22618 23860
rect 23198 23848 23204 23860
rect 22612 23820 23060 23848
rect 23159 23820 23204 23848
rect 22612 23808 22618 23820
rect 15378 23740 15384 23792
rect 15436 23780 15442 23792
rect 15473 23783 15531 23789
rect 15473 23780 15485 23783
rect 15436 23752 15485 23780
rect 15436 23740 15442 23752
rect 15473 23749 15485 23752
rect 15519 23749 15531 23783
rect 18506 23780 18512 23792
rect 18467 23752 18512 23780
rect 15473 23743 15531 23749
rect 18506 23740 18512 23752
rect 18564 23780 18570 23792
rect 19150 23780 19156 23792
rect 18564 23752 19156 23780
rect 18564 23740 18570 23752
rect 19150 23740 19156 23752
rect 19208 23740 19214 23792
rect 19797 23783 19855 23789
rect 19797 23749 19809 23783
rect 19843 23780 19855 23783
rect 23032 23780 23060 23820
rect 23198 23808 23204 23820
rect 23256 23808 23262 23860
rect 24762 23808 24768 23860
rect 24820 23848 24826 23860
rect 25041 23851 25099 23857
rect 25041 23848 25053 23851
rect 24820 23820 25053 23848
rect 24820 23808 24826 23820
rect 25041 23817 25053 23820
rect 25087 23817 25099 23851
rect 25041 23811 25099 23817
rect 25409 23851 25467 23857
rect 25409 23817 25421 23851
rect 25455 23848 25467 23851
rect 25682 23848 25688 23860
rect 25455 23820 25688 23848
rect 25455 23817 25467 23820
rect 25409 23811 25467 23817
rect 25314 23780 25320 23792
rect 19843 23752 22256 23780
rect 23032 23752 25320 23780
rect 19843 23749 19855 23752
rect 19797 23743 19855 23749
rect 12526 23721 12532 23724
rect 11624 23684 12434 23712
rect 11517 23675 11575 23681
rect 12520 23675 12532 23721
rect 12584 23712 12590 23724
rect 12584 23684 12620 23712
rect 9364 23616 9812 23644
rect 9953 23647 10011 23653
rect 9364 23604 9370 23616
rect 9953 23613 9965 23647
rect 9999 23644 10011 23647
rect 10226 23644 10232 23656
rect 9999 23616 10232 23644
rect 9999 23613 10011 23616
rect 9953 23607 10011 23613
rect 10226 23604 10232 23616
rect 10284 23644 10290 23656
rect 10594 23644 10600 23656
rect 10284 23616 10600 23644
rect 10284 23604 10290 23616
rect 10594 23604 10600 23616
rect 10652 23644 10658 23656
rect 11532 23644 11560 23675
rect 12526 23672 12532 23675
rect 12584 23672 12590 23684
rect 13538 23672 13544 23724
rect 13596 23712 13602 23724
rect 14369 23715 14427 23721
rect 14369 23712 14381 23715
rect 13596 23684 14381 23712
rect 13596 23672 13602 23684
rect 14369 23681 14381 23684
rect 14415 23712 14427 23715
rect 14734 23712 14740 23724
rect 14415 23684 14740 23712
rect 14415 23681 14427 23684
rect 14369 23675 14427 23681
rect 14734 23672 14740 23684
rect 14792 23672 14798 23724
rect 17218 23712 17224 23724
rect 17179 23684 17224 23712
rect 17218 23672 17224 23684
rect 17276 23672 17282 23724
rect 18785 23715 18843 23721
rect 18785 23681 18797 23715
rect 18831 23681 18843 23715
rect 19518 23712 19524 23724
rect 18785 23675 18843 23681
rect 19306 23684 19524 23712
rect 10652 23616 11560 23644
rect 10652 23604 10658 23616
rect 11698 23604 11704 23656
rect 11756 23644 11762 23656
rect 11793 23647 11851 23653
rect 11793 23644 11805 23647
rect 11756 23616 11805 23644
rect 11756 23604 11762 23616
rect 11793 23613 11805 23616
rect 11839 23613 11851 23647
rect 11793 23607 11851 23613
rect 11882 23604 11888 23656
rect 11940 23644 11946 23656
rect 12253 23647 12311 23653
rect 12253 23644 12265 23647
rect 11940 23616 12265 23644
rect 11940 23604 11946 23616
rect 12253 23613 12265 23616
rect 12299 23613 12311 23647
rect 12253 23607 12311 23613
rect 14093 23647 14151 23653
rect 14093 23613 14105 23647
rect 14139 23613 14151 23647
rect 14093 23607 14151 23613
rect 8018 23576 8024 23588
rect 7760 23548 8024 23576
rect 8018 23536 8024 23548
rect 8076 23576 8082 23588
rect 10321 23579 10379 23585
rect 10321 23576 10333 23579
rect 8076 23548 10333 23576
rect 8076 23536 8082 23548
rect 10321 23545 10333 23548
rect 10367 23545 10379 23579
rect 10321 23539 10379 23545
rect 11609 23579 11667 23585
rect 11609 23545 11621 23579
rect 11655 23576 11667 23579
rect 13633 23579 13691 23585
rect 11655 23548 12020 23576
rect 11655 23545 11667 23548
rect 11609 23539 11667 23545
rect 8478 23508 8484 23520
rect 4540 23480 8484 23508
rect 8478 23468 8484 23480
rect 8536 23468 8542 23520
rect 9030 23468 9036 23520
rect 9088 23508 9094 23520
rect 10873 23511 10931 23517
rect 9088 23480 9133 23508
rect 9088 23468 9094 23480
rect 10873 23477 10885 23511
rect 10919 23508 10931 23511
rect 11514 23508 11520 23520
rect 10919 23480 11520 23508
rect 10919 23477 10931 23480
rect 10873 23471 10931 23477
rect 11514 23468 11520 23480
rect 11572 23468 11578 23520
rect 11992 23508 12020 23548
rect 13633 23545 13645 23579
rect 13679 23576 13691 23579
rect 14108 23576 14136 23607
rect 16666 23604 16672 23656
rect 16724 23644 16730 23656
rect 17313 23647 17371 23653
rect 17313 23644 17325 23647
rect 16724 23616 17325 23644
rect 16724 23604 16730 23616
rect 17313 23613 17325 23616
rect 17359 23644 17371 23647
rect 18506 23644 18512 23656
rect 17359 23616 18512 23644
rect 17359 23613 17371 23616
rect 17313 23607 17371 23613
rect 18506 23604 18512 23616
rect 18564 23604 18570 23656
rect 18690 23644 18696 23656
rect 18651 23616 18696 23644
rect 18690 23604 18696 23616
rect 18748 23604 18754 23656
rect 14274 23576 14280 23588
rect 13679 23548 14280 23576
rect 13679 23545 13691 23548
rect 13633 23539 13691 23545
rect 14274 23536 14280 23548
rect 14332 23536 14338 23588
rect 15841 23579 15899 23585
rect 15841 23545 15853 23579
rect 15887 23576 15899 23579
rect 18800 23576 18828 23675
rect 19306 23656 19334 23684
rect 19518 23672 19524 23684
rect 19576 23672 19582 23724
rect 19613 23715 19671 23721
rect 19613 23681 19625 23715
rect 19659 23712 19671 23715
rect 19702 23712 19708 23724
rect 19659 23684 19708 23712
rect 19659 23681 19671 23684
rect 19613 23675 19671 23681
rect 19702 23672 19708 23684
rect 19760 23712 19766 23724
rect 19886 23712 19892 23724
rect 19760 23684 19892 23712
rect 19760 23672 19766 23684
rect 19886 23672 19892 23684
rect 19944 23672 19950 23724
rect 21634 23712 21640 23724
rect 20272 23684 21640 23712
rect 19242 23604 19248 23656
rect 19300 23616 19334 23656
rect 20272 23653 20300 23684
rect 21634 23672 21640 23684
rect 21692 23712 21698 23724
rect 21821 23715 21879 23721
rect 21821 23712 21833 23715
rect 21692 23684 21833 23712
rect 21692 23672 21698 23684
rect 21821 23681 21833 23684
rect 21867 23681 21879 23715
rect 21821 23675 21879 23681
rect 22097 23715 22155 23721
rect 22097 23681 22109 23715
rect 22143 23681 22155 23715
rect 22097 23675 22155 23681
rect 20257 23647 20315 23653
rect 20257 23644 20269 23647
rect 20180 23616 20269 23644
rect 19300 23604 19306 23616
rect 19518 23576 19524 23588
rect 15887 23548 19524 23576
rect 15887 23545 15899 23548
rect 15841 23539 15899 23545
rect 19518 23536 19524 23548
rect 19576 23536 19582 23588
rect 13722 23508 13728 23520
rect 11992 23480 13728 23508
rect 13722 23468 13728 23480
rect 13780 23468 13786 23520
rect 13998 23468 14004 23520
rect 14056 23508 14062 23520
rect 15657 23511 15715 23517
rect 15657 23508 15669 23511
rect 14056 23480 15669 23508
rect 14056 23468 14062 23480
rect 15657 23477 15669 23480
rect 15703 23477 15715 23511
rect 15657 23471 15715 23477
rect 16942 23468 16948 23520
rect 17000 23508 17006 23520
rect 17221 23511 17279 23517
rect 17221 23508 17233 23511
rect 17000 23480 17233 23508
rect 17000 23468 17006 23480
rect 17221 23477 17233 23480
rect 17267 23477 17279 23511
rect 17221 23471 17279 23477
rect 17589 23511 17647 23517
rect 17589 23477 17601 23511
rect 17635 23508 17647 23511
rect 18046 23508 18052 23520
rect 17635 23480 18052 23508
rect 17635 23477 17647 23480
rect 17589 23471 17647 23477
rect 18046 23468 18052 23480
rect 18104 23468 18110 23520
rect 18230 23468 18236 23520
rect 18288 23508 18294 23520
rect 18509 23511 18567 23517
rect 18509 23508 18521 23511
rect 18288 23480 18521 23508
rect 18288 23468 18294 23480
rect 18509 23477 18521 23480
rect 18555 23508 18567 23511
rect 20180 23508 20208 23616
rect 20257 23613 20269 23616
rect 20303 23613 20315 23647
rect 20257 23607 20315 23613
rect 20533 23647 20591 23653
rect 20533 23613 20545 23647
rect 20579 23644 20591 23647
rect 20898 23644 20904 23656
rect 20579 23616 20904 23644
rect 20579 23613 20591 23616
rect 20533 23607 20591 23613
rect 20898 23604 20904 23616
rect 20956 23604 20962 23656
rect 21910 23644 21916 23656
rect 21871 23616 21916 23644
rect 21910 23604 21916 23616
rect 21968 23604 21974 23656
rect 21174 23536 21180 23588
rect 21232 23576 21238 23588
rect 22112 23576 22140 23675
rect 21232 23548 22140 23576
rect 21232 23536 21238 23548
rect 22002 23508 22008 23520
rect 18555 23480 20208 23508
rect 21963 23480 22008 23508
rect 18555 23477 18567 23480
rect 18509 23471 18567 23477
rect 22002 23468 22008 23480
rect 22060 23468 22066 23520
rect 22228 23508 22256 23752
rect 25314 23740 25320 23752
rect 25372 23740 25378 23792
rect 22370 23672 22376 23724
rect 22428 23712 22434 23724
rect 22741 23715 22799 23721
rect 22741 23712 22753 23715
rect 22428 23684 22753 23712
rect 22428 23672 22434 23684
rect 22741 23681 22753 23684
rect 22787 23681 22799 23715
rect 22741 23675 22799 23681
rect 23017 23715 23075 23721
rect 23017 23681 23029 23715
rect 23063 23712 23075 23715
rect 23106 23712 23112 23724
rect 23063 23684 23112 23712
rect 23063 23681 23075 23684
rect 23017 23675 23075 23681
rect 23106 23672 23112 23684
rect 23164 23672 23170 23724
rect 23382 23672 23388 23724
rect 23440 23712 23446 23724
rect 24029 23715 24087 23721
rect 24029 23712 24041 23715
rect 23440 23684 24041 23712
rect 23440 23672 23446 23684
rect 24029 23681 24041 23684
rect 24075 23681 24087 23715
rect 24029 23675 24087 23681
rect 24762 23672 24768 23724
rect 24820 23712 24826 23724
rect 25424 23712 25452 23811
rect 25682 23808 25688 23820
rect 25740 23808 25746 23860
rect 25498 23740 25504 23792
rect 25556 23780 25562 23792
rect 27154 23780 27160 23792
rect 25556 23752 25601 23780
rect 27115 23752 27160 23780
rect 25556 23740 25562 23752
rect 27154 23740 27160 23752
rect 27212 23740 27218 23792
rect 26421 23715 26479 23721
rect 26421 23712 26433 23715
rect 24820 23684 25452 23712
rect 25516 23684 26433 23712
rect 24820 23672 24826 23684
rect 22925 23647 22983 23653
rect 22925 23613 22937 23647
rect 22971 23644 22983 23647
rect 23290 23644 23296 23656
rect 22971 23616 23296 23644
rect 22971 23613 22983 23616
rect 22925 23607 22983 23613
rect 23290 23604 23296 23616
rect 23348 23604 23354 23656
rect 23753 23647 23811 23653
rect 23753 23613 23765 23647
rect 23799 23613 23811 23647
rect 23753 23607 23811 23613
rect 23768 23576 23796 23607
rect 24394 23604 24400 23656
rect 24452 23644 24458 23656
rect 25516 23644 25544 23684
rect 26421 23681 26433 23684
rect 26467 23681 26479 23715
rect 26421 23675 26479 23681
rect 24452 23616 25544 23644
rect 24452 23604 24458 23616
rect 25590 23604 25596 23656
rect 25648 23644 25654 23656
rect 27172 23644 27200 23740
rect 25648 23616 25693 23644
rect 25976 23616 27200 23644
rect 25648 23604 25654 23616
rect 25682 23576 25688 23588
rect 23768 23548 25688 23576
rect 25682 23536 25688 23548
rect 25740 23576 25746 23588
rect 25976 23576 26004 23616
rect 25740 23548 26004 23576
rect 26237 23579 26295 23585
rect 25740 23536 25746 23548
rect 26237 23545 26249 23579
rect 26283 23576 26295 23579
rect 27430 23576 27436 23588
rect 26283 23548 27436 23576
rect 26283 23545 26295 23548
rect 26237 23539 26295 23545
rect 27430 23536 27436 23548
rect 27488 23536 27494 23588
rect 22554 23508 22560 23520
rect 22228 23480 22560 23508
rect 22554 23468 22560 23480
rect 22612 23508 22618 23520
rect 22741 23511 22799 23517
rect 22741 23508 22753 23511
rect 22612 23480 22753 23508
rect 22612 23468 22618 23480
rect 22741 23477 22753 23480
rect 22787 23477 22799 23511
rect 22741 23471 22799 23477
rect 25314 23468 25320 23520
rect 25372 23508 25378 23520
rect 27249 23511 27307 23517
rect 27249 23508 27261 23511
rect 25372 23480 27261 23508
rect 25372 23468 25378 23480
rect 27249 23477 27261 23480
rect 27295 23477 27307 23511
rect 27249 23471 27307 23477
rect 1104 23418 28060 23440
rect 1104 23366 5442 23418
rect 5494 23366 5506 23418
rect 5558 23366 5570 23418
rect 5622 23366 5634 23418
rect 5686 23366 5698 23418
rect 5750 23366 14428 23418
rect 14480 23366 14492 23418
rect 14544 23366 14556 23418
rect 14608 23366 14620 23418
rect 14672 23366 14684 23418
rect 14736 23366 23413 23418
rect 23465 23366 23477 23418
rect 23529 23366 23541 23418
rect 23593 23366 23605 23418
rect 23657 23366 23669 23418
rect 23721 23366 28060 23418
rect 1104 23344 28060 23366
rect 2501 23307 2559 23313
rect 2501 23273 2513 23307
rect 2547 23304 2559 23307
rect 3786 23304 3792 23316
rect 2547 23276 3792 23304
rect 2547 23273 2559 23276
rect 2501 23267 2559 23273
rect 3786 23264 3792 23276
rect 3844 23264 3850 23316
rect 5902 23304 5908 23316
rect 5863 23276 5908 23304
rect 5902 23264 5908 23276
rect 5960 23264 5966 23316
rect 6362 23264 6368 23316
rect 6420 23304 6426 23316
rect 6825 23307 6883 23313
rect 6825 23304 6837 23307
rect 6420 23276 6837 23304
rect 6420 23264 6426 23276
rect 6825 23273 6837 23276
rect 6871 23273 6883 23307
rect 6825 23267 6883 23273
rect 6914 23264 6920 23316
rect 6972 23304 6978 23316
rect 10321 23307 10379 23313
rect 10321 23304 10333 23307
rect 6972 23276 10333 23304
rect 6972 23264 6978 23276
rect 10321 23273 10333 23276
rect 10367 23304 10379 23307
rect 10778 23304 10784 23316
rect 10367 23276 10784 23304
rect 10367 23273 10379 23276
rect 10321 23267 10379 23273
rect 10778 23264 10784 23276
rect 10836 23264 10842 23316
rect 12161 23307 12219 23313
rect 12161 23273 12173 23307
rect 12207 23304 12219 23307
rect 12526 23304 12532 23316
rect 12207 23276 12532 23304
rect 12207 23273 12219 23276
rect 12161 23267 12219 23273
rect 12526 23264 12532 23276
rect 12584 23264 12590 23316
rect 13722 23264 13728 23316
rect 13780 23304 13786 23316
rect 15197 23307 15255 23313
rect 13780 23276 14780 23304
rect 13780 23264 13786 23276
rect 5350 23236 5356 23248
rect 4356 23208 5356 23236
rect 4356 23177 4384 23208
rect 5350 23196 5356 23208
rect 5408 23196 5414 23248
rect 6454 23196 6460 23248
rect 6512 23236 6518 23248
rect 7469 23239 7527 23245
rect 7469 23236 7481 23239
rect 6512 23208 7481 23236
rect 6512 23196 6518 23208
rect 7469 23205 7481 23208
rect 7515 23205 7527 23239
rect 7469 23199 7527 23205
rect 7558 23196 7564 23248
rect 7616 23236 7622 23248
rect 7926 23236 7932 23248
rect 7616 23208 7932 23236
rect 7616 23196 7622 23208
rect 7926 23196 7932 23208
rect 7984 23196 7990 23248
rect 8478 23196 8484 23248
rect 8536 23236 8542 23248
rect 8846 23236 8852 23248
rect 8536 23208 8852 23236
rect 8536 23196 8542 23208
rect 8846 23196 8852 23208
rect 8904 23236 8910 23248
rect 8904 23208 9628 23236
rect 8904 23196 8910 23208
rect 3053 23171 3111 23177
rect 3053 23137 3065 23171
rect 3099 23168 3111 23171
rect 4341 23171 4399 23177
rect 4341 23168 4353 23171
rect 3099 23140 4353 23168
rect 3099 23137 3111 23140
rect 3053 23131 3111 23137
rect 4341 23137 4353 23140
rect 4387 23137 4399 23171
rect 4341 23131 4399 23137
rect 4430 23128 4436 23180
rect 4488 23168 4494 23180
rect 4488 23140 5764 23168
rect 4488 23128 4494 23140
rect 2041 23103 2099 23109
rect 2041 23069 2053 23103
rect 2087 23100 2099 23103
rect 2869 23103 2927 23109
rect 2087 23072 2452 23100
rect 2087 23069 2099 23072
rect 2041 23063 2099 23069
rect 1857 22967 1915 22973
rect 1857 22933 1869 22967
rect 1903 22964 1915 22967
rect 2038 22964 2044 22976
rect 1903 22936 2044 22964
rect 1903 22933 1915 22936
rect 1857 22927 1915 22933
rect 2038 22924 2044 22936
rect 2096 22924 2102 22976
rect 2424 22973 2452 23072
rect 2869 23069 2881 23103
rect 2915 23100 2927 23103
rect 2958 23100 2964 23112
rect 2915 23072 2964 23100
rect 2915 23069 2927 23072
rect 2869 23063 2927 23069
rect 2958 23060 2964 23072
rect 3016 23100 3022 23112
rect 3142 23100 3148 23112
rect 3016 23072 3148 23100
rect 3016 23060 3022 23072
rect 3142 23060 3148 23072
rect 3200 23060 3206 23112
rect 4157 23103 4215 23109
rect 4157 23069 4169 23103
rect 4203 23100 4215 23103
rect 4246 23100 4252 23112
rect 4203 23072 4252 23100
rect 4203 23069 4215 23072
rect 4157 23063 4215 23069
rect 4246 23060 4252 23072
rect 4304 23060 4310 23112
rect 5074 23060 5080 23112
rect 5132 23100 5138 23112
rect 5736 23109 5764 23140
rect 7834 23128 7840 23180
rect 7892 23128 7898 23180
rect 9033 23171 9091 23177
rect 9033 23137 9045 23171
rect 9079 23137 9091 23171
rect 9033 23131 9091 23137
rect 5261 23103 5319 23109
rect 5261 23100 5273 23103
rect 5132 23072 5273 23100
rect 5132 23060 5138 23072
rect 5261 23069 5273 23072
rect 5307 23069 5319 23103
rect 5261 23063 5319 23069
rect 5721 23103 5779 23109
rect 5721 23069 5733 23103
rect 5767 23069 5779 23103
rect 5721 23063 5779 23069
rect 6733 23103 6791 23109
rect 6733 23069 6745 23103
rect 6779 23100 6791 23103
rect 7190 23100 7196 23112
rect 6779 23072 7196 23100
rect 6779 23069 6791 23072
rect 6733 23063 6791 23069
rect 7190 23060 7196 23072
rect 7248 23060 7254 23112
rect 7650 23100 7656 23112
rect 7611 23072 7656 23100
rect 7650 23060 7656 23072
rect 7708 23060 7714 23112
rect 7745 23103 7803 23109
rect 7745 23069 7757 23103
rect 7791 23100 7803 23103
rect 7852 23100 7880 23128
rect 8018 23100 8024 23112
rect 7791 23072 7880 23100
rect 7979 23072 8024 23100
rect 7791 23069 7803 23072
rect 7745 23063 7803 23069
rect 8018 23060 8024 23072
rect 8076 23060 8082 23112
rect 8110 23060 8116 23112
rect 8168 23100 8174 23112
rect 9048 23100 9076 23131
rect 9214 23128 9220 23180
rect 9272 23168 9278 23180
rect 9600 23168 9628 23208
rect 10686 23196 10692 23248
rect 10744 23236 10750 23248
rect 14645 23239 14703 23245
rect 14645 23236 14657 23239
rect 10744 23208 14657 23236
rect 10744 23196 10750 23208
rect 14645 23205 14657 23208
rect 14691 23205 14703 23239
rect 14752 23236 14780 23276
rect 15197 23273 15209 23307
rect 15243 23304 15255 23307
rect 16390 23304 16396 23316
rect 15243 23276 16396 23304
rect 15243 23273 15255 23276
rect 15197 23267 15255 23273
rect 16390 23264 16396 23276
rect 16448 23264 16454 23316
rect 18046 23264 18052 23316
rect 18104 23304 18110 23316
rect 19337 23307 19395 23313
rect 19337 23304 19349 23307
rect 18104 23276 19349 23304
rect 18104 23264 18110 23276
rect 19337 23273 19349 23276
rect 19383 23304 19395 23307
rect 20622 23304 20628 23316
rect 19383 23276 20628 23304
rect 19383 23273 19395 23276
rect 19337 23267 19395 23273
rect 20622 23264 20628 23276
rect 20680 23264 20686 23316
rect 20993 23307 21051 23313
rect 20993 23273 21005 23307
rect 21039 23304 21051 23307
rect 22002 23304 22008 23316
rect 21039 23276 22008 23304
rect 21039 23273 21051 23276
rect 20993 23267 21051 23273
rect 22002 23264 22008 23276
rect 22060 23264 22066 23316
rect 22554 23304 22560 23316
rect 22515 23276 22560 23304
rect 22554 23264 22560 23276
rect 22612 23264 22618 23316
rect 22738 23304 22744 23316
rect 22699 23276 22744 23304
rect 22738 23264 22744 23276
rect 22796 23264 22802 23316
rect 22830 23264 22836 23316
rect 22888 23304 22894 23316
rect 23201 23307 23259 23313
rect 23201 23304 23213 23307
rect 22888 23276 23213 23304
rect 22888 23264 22894 23276
rect 23201 23273 23213 23276
rect 23247 23273 23259 23307
rect 23201 23267 23259 23273
rect 24397 23307 24455 23313
rect 24397 23273 24409 23307
rect 24443 23304 24455 23307
rect 24578 23304 24584 23316
rect 24443 23276 24584 23304
rect 24443 23273 24455 23276
rect 24397 23267 24455 23273
rect 24578 23264 24584 23276
rect 24636 23264 24642 23316
rect 19705 23239 19763 23245
rect 14752 23208 15516 23236
rect 14645 23199 14703 23205
rect 9272 23140 9444 23168
rect 9600 23140 9720 23168
rect 9272 23128 9278 23140
rect 9306 23100 9312 23112
rect 8168 23072 9076 23100
rect 9267 23072 9312 23100
rect 8168 23060 8174 23072
rect 9306 23060 9312 23072
rect 9364 23060 9370 23112
rect 9416 23109 9444 23140
rect 9401 23103 9459 23109
rect 9401 23069 9413 23103
rect 9447 23069 9459 23103
rect 9401 23063 9459 23069
rect 9493 23103 9551 23109
rect 9493 23069 9505 23103
rect 9539 23100 9551 23103
rect 9582 23100 9588 23112
rect 9539 23072 9588 23100
rect 9539 23069 9551 23072
rect 9493 23063 9551 23069
rect 9582 23060 9588 23072
rect 9640 23060 9646 23112
rect 9692 23109 9720 23140
rect 10502 23128 10508 23180
rect 10560 23168 10566 23180
rect 10870 23168 10876 23180
rect 10560 23140 10876 23168
rect 10560 23128 10566 23140
rect 10870 23128 10876 23140
rect 10928 23128 10934 23180
rect 11609 23171 11667 23177
rect 11609 23137 11621 23171
rect 11655 23168 11667 23171
rect 12621 23171 12679 23177
rect 12621 23168 12633 23171
rect 11655 23140 12633 23168
rect 11655 23137 11667 23140
rect 11609 23131 11667 23137
rect 12621 23137 12633 23140
rect 12667 23137 12679 23171
rect 13998 23168 14004 23180
rect 12621 23131 12679 23137
rect 13372 23140 14004 23168
rect 9677 23103 9735 23109
rect 9677 23069 9689 23103
rect 9723 23069 9735 23103
rect 9677 23063 9735 23069
rect 9858 23060 9864 23112
rect 9916 23100 9922 23112
rect 11054 23100 11060 23112
rect 9916 23072 10364 23100
rect 11015 23072 11060 23100
rect 9916 23060 9922 23072
rect 4982 23032 4988 23044
rect 4943 23004 4988 23032
rect 4982 22992 4988 23004
rect 5040 22992 5046 23044
rect 5169 23035 5227 23041
rect 5169 23001 5181 23035
rect 5215 23032 5227 23035
rect 5350 23032 5356 23044
rect 5215 23004 5356 23032
rect 5215 23001 5227 23004
rect 5169 22995 5227 23001
rect 5350 22992 5356 23004
rect 5408 22992 5414 23044
rect 7558 22992 7564 23044
rect 7616 23032 7622 23044
rect 7837 23035 7895 23041
rect 7837 23032 7849 23035
rect 7616 23004 7849 23032
rect 7616 22992 7622 23004
rect 7837 23001 7849 23004
rect 7883 23001 7895 23035
rect 7837 22995 7895 23001
rect 8570 22992 8576 23044
rect 8628 23032 8634 23044
rect 8846 23032 8852 23044
rect 8628 23004 8852 23032
rect 8628 22992 8634 23004
rect 8846 22992 8852 23004
rect 8904 22992 8910 23044
rect 9030 22992 9036 23044
rect 9088 23032 9094 23044
rect 10229 23035 10287 23041
rect 10229 23032 10241 23035
rect 9088 23004 10241 23032
rect 9088 22992 9094 23004
rect 10229 23001 10241 23004
rect 10275 23001 10287 23035
rect 10336 23032 10364 23072
rect 11054 23060 11060 23072
rect 11112 23060 11118 23112
rect 11514 23100 11520 23112
rect 11475 23072 11520 23100
rect 11514 23060 11520 23072
rect 11572 23060 11578 23112
rect 11698 23100 11704 23112
rect 11659 23072 11704 23100
rect 11698 23060 11704 23072
rect 11756 23060 11762 23112
rect 12250 23060 12256 23112
rect 12308 23100 12314 23112
rect 12345 23103 12403 23109
rect 12345 23100 12357 23103
rect 12308 23072 12357 23100
rect 12308 23060 12314 23072
rect 12345 23069 12357 23072
rect 12391 23069 12403 23103
rect 12345 23063 12403 23069
rect 12437 23103 12495 23109
rect 12437 23069 12449 23103
rect 12483 23069 12495 23103
rect 12437 23063 12495 23069
rect 12452 23032 12480 23063
rect 12526 23060 12532 23112
rect 12584 23100 12590 23112
rect 13372 23109 13400 23140
rect 13998 23128 14004 23140
rect 14056 23128 14062 23180
rect 15488 23112 15516 23208
rect 19705 23205 19717 23239
rect 19751 23236 19763 23239
rect 19751 23208 20668 23236
rect 19751 23205 19763 23208
rect 19705 23199 19763 23205
rect 18417 23171 18475 23177
rect 18417 23137 18429 23171
rect 18463 23168 18475 23171
rect 18690 23168 18696 23180
rect 18463 23140 18696 23168
rect 18463 23137 18475 23140
rect 18417 23131 18475 23137
rect 18690 23128 18696 23140
rect 18748 23168 18754 23180
rect 19429 23171 19487 23177
rect 19429 23168 19441 23171
rect 18748 23140 19441 23168
rect 18748 23128 18754 23140
rect 19429 23137 19441 23140
rect 19475 23168 19487 23171
rect 19886 23168 19892 23180
rect 19475 23140 19892 23168
rect 19475 23137 19487 23140
rect 19429 23131 19487 23137
rect 19886 23128 19892 23140
rect 19944 23128 19950 23180
rect 13357 23103 13415 23109
rect 12584 23072 12629 23100
rect 12584 23060 12590 23072
rect 13357 23069 13369 23103
rect 13403 23069 13415 23103
rect 13538 23100 13544 23112
rect 13499 23072 13544 23100
rect 13357 23063 13415 23069
rect 13538 23060 13544 23072
rect 13596 23060 13602 23112
rect 14274 23060 14280 23112
rect 14332 23100 14338 23112
rect 14369 23103 14427 23109
rect 14369 23100 14381 23103
rect 14332 23072 14381 23100
rect 14332 23060 14338 23072
rect 14369 23069 14381 23072
rect 14415 23069 14427 23103
rect 14369 23063 14427 23069
rect 15102 23060 15108 23112
rect 15160 23100 15166 23112
rect 15381 23103 15439 23109
rect 15381 23100 15393 23103
rect 15160 23072 15393 23100
rect 15160 23060 15166 23072
rect 15381 23069 15393 23072
rect 15427 23069 15439 23103
rect 15381 23063 15439 23069
rect 15470 23060 15476 23112
rect 15528 23100 15534 23112
rect 15565 23103 15623 23109
rect 15565 23100 15577 23103
rect 15528 23072 15577 23100
rect 15528 23060 15534 23072
rect 15565 23069 15577 23072
rect 15611 23069 15623 23103
rect 15565 23063 15623 23069
rect 15654 23060 15660 23112
rect 15712 23100 15718 23112
rect 15712 23072 15757 23100
rect 15712 23060 15718 23072
rect 16482 23060 16488 23112
rect 16540 23100 16546 23112
rect 16577 23103 16635 23109
rect 16577 23100 16589 23103
rect 16540 23072 16589 23100
rect 16540 23060 16546 23072
rect 16577 23069 16589 23072
rect 16623 23069 16635 23103
rect 16577 23063 16635 23069
rect 16850 23060 16856 23112
rect 16908 23060 16914 23112
rect 18322 23100 18328 23112
rect 18283 23072 18328 23100
rect 18322 23060 18328 23072
rect 18380 23060 18386 23112
rect 18506 23100 18512 23112
rect 18467 23072 18512 23100
rect 18506 23060 18512 23072
rect 18564 23060 18570 23112
rect 19518 23100 19524 23112
rect 18616 23072 19380 23100
rect 19479 23072 19524 23100
rect 12618 23032 12624 23044
rect 10336 23004 12624 23032
rect 10229 22995 10287 23001
rect 12618 22992 12624 23004
rect 12676 22992 12682 23044
rect 14090 23032 14096 23044
rect 14051 23004 14096 23032
rect 14090 22992 14096 23004
rect 14148 22992 14154 23044
rect 17589 23035 17647 23041
rect 17589 23001 17601 23035
rect 17635 23001 17647 23035
rect 18616 23032 18644 23072
rect 17589 22995 17647 23001
rect 18524 23004 18644 23032
rect 2409 22967 2467 22973
rect 2409 22933 2421 22967
rect 2455 22964 2467 22967
rect 2590 22964 2596 22976
rect 2455 22936 2596 22964
rect 2455 22933 2467 22936
rect 2409 22927 2467 22933
rect 2590 22924 2596 22936
rect 2648 22924 2654 22976
rect 2958 22924 2964 22976
rect 3016 22964 3022 22976
rect 3016 22936 3061 22964
rect 3016 22924 3022 22936
rect 3510 22924 3516 22976
rect 3568 22964 3574 22976
rect 3789 22967 3847 22973
rect 3789 22964 3801 22967
rect 3568 22936 3801 22964
rect 3568 22924 3574 22936
rect 3789 22933 3801 22936
rect 3835 22933 3847 22967
rect 3789 22927 3847 22933
rect 3970 22924 3976 22976
rect 4028 22964 4034 22976
rect 4249 22967 4307 22973
rect 4249 22964 4261 22967
rect 4028 22936 4261 22964
rect 4028 22924 4034 22936
rect 4249 22933 4261 22936
rect 4295 22933 4307 22967
rect 4249 22927 4307 22933
rect 5261 22967 5319 22973
rect 5261 22933 5273 22967
rect 5307 22964 5319 22967
rect 5902 22964 5908 22976
rect 5307 22936 5908 22964
rect 5307 22933 5319 22936
rect 5261 22927 5319 22933
rect 5902 22924 5908 22936
rect 5960 22924 5966 22976
rect 7650 22924 7656 22976
rect 7708 22964 7714 22976
rect 9048 22964 9076 22992
rect 7708 22936 9076 22964
rect 10873 22967 10931 22973
rect 7708 22924 7714 22936
rect 10873 22933 10885 22967
rect 10919 22964 10931 22967
rect 12342 22964 12348 22976
rect 10919 22936 12348 22964
rect 10919 22933 10931 22936
rect 10873 22927 10931 22933
rect 12342 22924 12348 22936
rect 12400 22924 12406 22976
rect 13538 22964 13544 22976
rect 13499 22936 13544 22964
rect 13538 22924 13544 22936
rect 13596 22924 13602 22976
rect 14274 22964 14280 22976
rect 14235 22936 14280 22964
rect 14274 22924 14280 22936
rect 14332 22924 14338 22976
rect 14458 22964 14464 22976
rect 14419 22936 14464 22964
rect 14458 22924 14464 22936
rect 14516 22924 14522 22976
rect 17604 22964 17632 22995
rect 18524 22964 18552 23004
rect 19150 22992 19156 23044
rect 19208 23032 19214 23044
rect 19245 23035 19303 23041
rect 19245 23032 19257 23035
rect 19208 23004 19257 23032
rect 19208 22992 19214 23004
rect 19245 23001 19257 23004
rect 19291 23001 19303 23035
rect 19352 23032 19380 23072
rect 19518 23060 19524 23072
rect 19576 23060 19582 23112
rect 19702 23032 19708 23044
rect 19352 23004 19708 23032
rect 19245 22995 19303 23001
rect 19702 22992 19708 23004
rect 19760 22992 19766 23044
rect 20640 23032 20668 23208
rect 20898 23196 20904 23248
rect 20956 23196 20962 23248
rect 21174 23196 21180 23248
rect 21232 23196 21238 23248
rect 23661 23239 23719 23245
rect 21392 23208 22508 23236
rect 20916 23168 20944 23196
rect 21082 23168 21088 23180
rect 20732 23140 21088 23168
rect 20732 23109 20760 23140
rect 21082 23128 21088 23140
rect 21140 23128 21146 23180
rect 20717 23103 20775 23109
rect 20717 23069 20729 23103
rect 20763 23069 20775 23103
rect 20898 23100 20904 23112
rect 20859 23072 20904 23100
rect 20717 23063 20775 23069
rect 20898 23060 20904 23072
rect 20956 23060 20962 23112
rect 20993 23103 21051 23109
rect 20993 23069 21005 23103
rect 21039 23100 21051 23103
rect 21192 23100 21220 23196
rect 21039 23072 21220 23100
rect 21039 23069 21051 23072
rect 20993 23063 21051 23069
rect 21392 23032 21420 23208
rect 21542 23128 21548 23180
rect 21600 23168 21606 23180
rect 21910 23168 21916 23180
rect 21600 23140 21916 23168
rect 21600 23128 21606 23140
rect 21910 23128 21916 23140
rect 21968 23168 21974 23180
rect 22186 23168 22192 23180
rect 21968 23140 22192 23168
rect 21968 23128 21974 23140
rect 22186 23128 22192 23140
rect 22244 23168 22250 23180
rect 22373 23171 22431 23177
rect 22373 23168 22385 23171
rect 22244 23140 22385 23168
rect 22244 23128 22250 23140
rect 22373 23137 22385 23140
rect 22419 23137 22431 23171
rect 22480 23168 22508 23208
rect 23124 23208 23428 23236
rect 23124 23168 23152 23208
rect 23290 23168 23296 23180
rect 22480 23140 23152 23168
rect 23251 23140 23296 23168
rect 22373 23131 22431 23137
rect 23290 23128 23296 23140
rect 23348 23128 23354 23180
rect 23400 23168 23428 23208
rect 23661 23205 23673 23239
rect 23707 23236 23719 23239
rect 25590 23236 25596 23248
rect 23707 23208 25596 23236
rect 23707 23205 23719 23208
rect 23661 23199 23719 23205
rect 25590 23196 25596 23208
rect 25648 23196 25654 23248
rect 24949 23171 25007 23177
rect 24949 23168 24961 23171
rect 23400 23140 24961 23168
rect 24949 23137 24961 23140
rect 24995 23137 25007 23171
rect 25958 23168 25964 23180
rect 25919 23140 25964 23168
rect 24949 23131 25007 23137
rect 25958 23128 25964 23140
rect 26016 23128 26022 23180
rect 21634 23100 21640 23112
rect 21595 23072 21640 23100
rect 21634 23060 21640 23072
rect 21692 23060 21698 23112
rect 21821 23103 21879 23109
rect 21821 23069 21833 23103
rect 21867 23069 21879 23103
rect 21821 23063 21879 23069
rect 22557 23103 22615 23109
rect 22557 23069 22569 23103
rect 22603 23100 22615 23103
rect 23106 23100 23112 23112
rect 22603 23072 23112 23100
rect 22603 23069 22615 23072
rect 22557 23063 22615 23069
rect 20640 23004 21420 23032
rect 21450 22992 21456 23044
rect 21508 23032 21514 23044
rect 21836 23032 21864 23063
rect 23106 23060 23112 23072
rect 23164 23100 23170 23112
rect 23477 23103 23535 23109
rect 23477 23100 23489 23103
rect 23164 23072 23489 23100
rect 23164 23060 23170 23072
rect 23477 23069 23489 23072
rect 23523 23069 23535 23103
rect 24762 23100 24768 23112
rect 24723 23072 24768 23100
rect 23477 23063 23535 23069
rect 24762 23060 24768 23072
rect 24820 23060 24826 23112
rect 21508 23004 21864 23032
rect 22281 23035 22339 23041
rect 21508 22992 21514 23004
rect 22281 23001 22293 23035
rect 22327 23032 22339 23035
rect 22370 23032 22376 23044
rect 22327 23004 22376 23032
rect 22327 23001 22339 23004
rect 22281 22995 22339 23001
rect 22370 22992 22376 23004
rect 22428 22992 22434 23044
rect 23201 23035 23259 23041
rect 23201 23001 23213 23035
rect 23247 23032 23259 23035
rect 23382 23032 23388 23044
rect 23247 23004 23388 23032
rect 23247 23001 23259 23004
rect 23201 22995 23259 23001
rect 23382 22992 23388 23004
rect 23440 22992 23446 23044
rect 26228 23035 26286 23041
rect 26228 23001 26240 23035
rect 26274 23032 26286 23035
rect 26326 23032 26332 23044
rect 26274 23004 26332 23032
rect 26274 23001 26286 23004
rect 26228 22995 26286 23001
rect 26326 22992 26332 23004
rect 26384 22992 26390 23044
rect 17604 22936 18552 22964
rect 19610 22924 19616 22976
rect 19668 22964 19674 22976
rect 21177 22967 21235 22973
rect 21177 22964 21189 22967
rect 19668 22936 21189 22964
rect 19668 22924 19674 22936
rect 21177 22933 21189 22936
rect 21223 22933 21235 22967
rect 21177 22927 21235 22933
rect 21729 22967 21787 22973
rect 21729 22933 21741 22967
rect 21775 22964 21787 22967
rect 22462 22964 22468 22976
rect 21775 22936 22468 22964
rect 21775 22933 21787 22936
rect 21729 22927 21787 22933
rect 22462 22924 22468 22936
rect 22520 22924 22526 22976
rect 24210 22924 24216 22976
rect 24268 22964 24274 22976
rect 24578 22964 24584 22976
rect 24268 22936 24584 22964
rect 24268 22924 24274 22936
rect 24578 22924 24584 22936
rect 24636 22964 24642 22976
rect 24857 22967 24915 22973
rect 24857 22964 24869 22967
rect 24636 22936 24869 22964
rect 24636 22924 24642 22936
rect 24857 22933 24869 22936
rect 24903 22933 24915 22967
rect 24857 22927 24915 22933
rect 25498 22924 25504 22976
rect 25556 22964 25562 22976
rect 27341 22967 27399 22973
rect 27341 22964 27353 22967
rect 25556 22936 27353 22964
rect 25556 22924 25562 22936
rect 27341 22933 27353 22936
rect 27387 22933 27399 22967
rect 27341 22927 27399 22933
rect 1104 22874 28060 22896
rect 1104 22822 9935 22874
rect 9987 22822 9999 22874
rect 10051 22822 10063 22874
rect 10115 22822 10127 22874
rect 10179 22822 10191 22874
rect 10243 22822 18920 22874
rect 18972 22822 18984 22874
rect 19036 22822 19048 22874
rect 19100 22822 19112 22874
rect 19164 22822 19176 22874
rect 19228 22822 28060 22874
rect 1104 22800 28060 22822
rect 1765 22763 1823 22769
rect 1765 22729 1777 22763
rect 1811 22729 1823 22763
rect 1765 22723 1823 22729
rect 2869 22763 2927 22769
rect 2869 22729 2881 22763
rect 2915 22760 2927 22763
rect 2958 22760 2964 22772
rect 2915 22732 2964 22760
rect 2915 22729 2927 22732
rect 2869 22723 2927 22729
rect 1780 22692 1808 22723
rect 2958 22720 2964 22732
rect 3016 22720 3022 22772
rect 3513 22763 3571 22769
rect 3513 22729 3525 22763
rect 3559 22760 3571 22763
rect 3970 22760 3976 22772
rect 3559 22732 3976 22760
rect 3559 22729 3571 22732
rect 3513 22723 3571 22729
rect 3970 22720 3976 22732
rect 4028 22720 4034 22772
rect 4893 22763 4951 22769
rect 4893 22760 4905 22763
rect 4356 22732 4905 22760
rect 3786 22692 3792 22704
rect 1780 22664 3792 22692
rect 3786 22652 3792 22664
rect 3844 22652 3850 22704
rect 4249 22695 4307 22701
rect 3896 22664 4200 22692
rect 1949 22627 2007 22633
rect 1949 22593 1961 22627
rect 1995 22624 2007 22627
rect 2777 22627 2835 22633
rect 1995 22596 2360 22624
rect 1995 22593 2007 22596
rect 1949 22587 2007 22593
rect 2332 22429 2360 22596
rect 2777 22593 2789 22627
rect 2823 22593 2835 22627
rect 2777 22587 2835 22593
rect 3421 22627 3479 22633
rect 3421 22593 3433 22627
rect 3467 22624 3479 22627
rect 3896 22624 3924 22664
rect 4062 22624 4068 22636
rect 3467 22596 3924 22624
rect 4023 22596 4068 22624
rect 3467 22593 3479 22596
rect 3421 22587 3479 22593
rect 2792 22556 2820 22587
rect 4062 22584 4068 22596
rect 4120 22584 4126 22636
rect 4172 22624 4200 22664
rect 4249 22661 4261 22695
rect 4295 22692 4307 22695
rect 4356 22692 4384 22732
rect 4893 22729 4905 22732
rect 4939 22760 4951 22763
rect 5350 22760 5356 22772
rect 4939 22732 5356 22760
rect 4939 22729 4951 22732
rect 4893 22723 4951 22729
rect 5350 22720 5356 22732
rect 5408 22720 5414 22772
rect 6270 22720 6276 22772
rect 6328 22760 6334 22772
rect 6822 22760 6828 22772
rect 6328 22732 6828 22760
rect 6328 22720 6334 22732
rect 6822 22720 6828 22732
rect 6880 22720 6886 22772
rect 7282 22720 7288 22772
rect 7340 22760 7346 22772
rect 7837 22763 7895 22769
rect 7837 22760 7849 22763
rect 7340 22732 7849 22760
rect 7340 22720 7346 22732
rect 7837 22729 7849 22732
rect 7883 22729 7895 22763
rect 7837 22723 7895 22729
rect 8018 22720 8024 22772
rect 8076 22760 8082 22772
rect 8294 22760 8300 22772
rect 8076 22732 8300 22760
rect 8076 22720 8082 22732
rect 8294 22720 8300 22732
rect 8352 22720 8358 22772
rect 9858 22760 9864 22772
rect 8864 22732 9864 22760
rect 4295 22664 4384 22692
rect 4295 22661 4307 22664
rect 4249 22655 4307 22661
rect 4430 22652 4436 22704
rect 4488 22692 4494 22704
rect 6457 22695 6515 22701
rect 6457 22692 6469 22695
rect 4488 22664 6469 22692
rect 4488 22652 4494 22664
rect 6457 22661 6469 22664
rect 6503 22661 6515 22695
rect 6457 22655 6515 22661
rect 7006 22652 7012 22704
rect 7064 22692 7070 22704
rect 7064 22664 7328 22692
rect 7064 22652 7070 22664
rect 5077 22627 5135 22633
rect 5077 22624 5089 22627
rect 4172 22596 5089 22624
rect 5077 22593 5089 22596
rect 5123 22593 5135 22627
rect 5077 22587 5135 22593
rect 5169 22627 5227 22633
rect 5169 22593 5181 22627
rect 5215 22593 5227 22627
rect 5442 22624 5448 22636
rect 5403 22596 5448 22624
rect 5169 22587 5227 22593
rect 4154 22556 4160 22568
rect 2792 22528 4160 22556
rect 4154 22516 4160 22528
rect 4212 22516 4218 22568
rect 4338 22448 4344 22500
rect 4396 22488 4402 22500
rect 4522 22488 4528 22500
rect 4396 22460 4528 22488
rect 4396 22448 4402 22460
rect 4522 22448 4528 22460
rect 4580 22448 4586 22500
rect 5092 22488 5120 22587
rect 5184 22556 5212 22587
rect 5442 22584 5448 22596
rect 5500 22584 5506 22636
rect 7101 22627 7159 22633
rect 7101 22593 7113 22627
rect 7147 22624 7159 22627
rect 7190 22624 7196 22636
rect 7147 22596 7196 22624
rect 7147 22593 7159 22596
rect 7101 22587 7159 22593
rect 7190 22584 7196 22596
rect 7248 22584 7254 22636
rect 7300 22633 7328 22664
rect 7285 22627 7343 22633
rect 7285 22593 7297 22627
rect 7331 22624 7343 22627
rect 7466 22624 7472 22636
rect 7331 22596 7472 22624
rect 7331 22593 7343 22596
rect 7285 22587 7343 22593
rect 7466 22584 7472 22596
rect 7524 22584 7530 22636
rect 8864 22633 8892 22732
rect 9858 22720 9864 22732
rect 9916 22760 9922 22772
rect 10137 22763 10195 22769
rect 10137 22760 10149 22763
rect 9916 22732 10149 22760
rect 9916 22720 9922 22732
rect 10137 22729 10149 22732
rect 10183 22729 10195 22763
rect 10137 22723 10195 22729
rect 11054 22720 11060 22772
rect 11112 22760 11118 22772
rect 12894 22760 12900 22772
rect 11112 22732 12900 22760
rect 11112 22720 11118 22732
rect 12894 22720 12900 22732
rect 12952 22720 12958 22772
rect 16025 22763 16083 22769
rect 16025 22729 16037 22763
rect 16071 22760 16083 22763
rect 17678 22760 17684 22772
rect 16071 22732 17684 22760
rect 16071 22729 16083 22732
rect 16025 22723 16083 22729
rect 17678 22720 17684 22732
rect 17736 22720 17742 22772
rect 17954 22720 17960 22772
rect 18012 22760 18018 22772
rect 18506 22760 18512 22772
rect 18012 22732 18512 22760
rect 18012 22720 18018 22732
rect 18506 22720 18512 22732
rect 18564 22720 18570 22772
rect 18598 22720 18604 22772
rect 18656 22760 18662 22772
rect 19426 22760 19432 22772
rect 18656 22732 19432 22760
rect 18656 22720 18662 22732
rect 19426 22720 19432 22732
rect 19484 22720 19490 22772
rect 19794 22720 19800 22772
rect 19852 22760 19858 22772
rect 19981 22763 20039 22769
rect 19981 22760 19993 22763
rect 19852 22732 19993 22760
rect 19852 22720 19858 22732
rect 19981 22729 19993 22732
rect 20027 22729 20039 22763
rect 19981 22723 20039 22729
rect 20622 22720 20628 22772
rect 20680 22760 20686 22772
rect 20806 22760 20812 22772
rect 20680 22732 20812 22760
rect 20680 22720 20686 22732
rect 20806 22720 20812 22732
rect 20864 22720 20870 22772
rect 21634 22720 21640 22772
rect 21692 22760 21698 22772
rect 22738 22760 22744 22772
rect 21692 22732 22744 22760
rect 21692 22720 21698 22732
rect 22738 22720 22744 22732
rect 22796 22720 22802 22772
rect 24118 22720 24124 22772
rect 24176 22760 24182 22772
rect 24394 22760 24400 22772
rect 24176 22732 24400 22760
rect 24176 22720 24182 22732
rect 24394 22720 24400 22732
rect 24452 22720 24458 22772
rect 25498 22760 25504 22772
rect 25459 22732 25504 22760
rect 25498 22720 25504 22732
rect 25556 22720 25562 22772
rect 26970 22720 26976 22772
rect 27028 22760 27034 22772
rect 27341 22763 27399 22769
rect 27341 22760 27353 22763
rect 27028 22732 27353 22760
rect 27028 22720 27034 22732
rect 27341 22729 27353 22732
rect 27387 22729 27399 22763
rect 27341 22723 27399 22729
rect 9048 22664 9996 22692
rect 9048 22633 9076 22664
rect 7745 22627 7803 22633
rect 7745 22593 7757 22627
rect 7791 22593 7803 22627
rect 7745 22587 7803 22593
rect 8849 22627 8907 22633
rect 8849 22593 8861 22627
rect 8895 22593 8907 22627
rect 8849 22587 8907 22593
rect 9033 22627 9091 22633
rect 9033 22593 9045 22627
rect 9079 22593 9091 22627
rect 9033 22587 9091 22593
rect 6086 22556 6092 22568
rect 5184 22528 6092 22556
rect 6086 22516 6092 22528
rect 6144 22556 6150 22568
rect 6638 22556 6644 22568
rect 6144 22528 6644 22556
rect 6144 22516 6150 22528
rect 6638 22516 6644 22528
rect 6696 22516 6702 22568
rect 6914 22516 6920 22568
rect 6972 22556 6978 22568
rect 7760 22556 7788 22587
rect 9398 22584 9404 22636
rect 9456 22624 9462 22636
rect 9585 22627 9643 22633
rect 9585 22624 9597 22627
rect 9456 22596 9597 22624
rect 9456 22584 9462 22596
rect 9585 22593 9597 22596
rect 9631 22593 9643 22627
rect 9766 22624 9772 22636
rect 9727 22596 9772 22624
rect 9585 22587 9643 22593
rect 9766 22584 9772 22596
rect 9824 22584 9830 22636
rect 9968 22633 9996 22664
rect 11882 22652 11888 22704
rect 11940 22692 11946 22704
rect 11940 22664 12388 22692
rect 11940 22652 11946 22664
rect 9861 22627 9919 22633
rect 9861 22593 9873 22627
rect 9907 22593 9919 22627
rect 9861 22587 9919 22593
rect 9953 22627 10011 22633
rect 9953 22593 9965 22627
rect 9999 22624 10011 22627
rect 10318 22624 10324 22636
rect 9999 22596 10324 22624
rect 9999 22593 10011 22596
rect 9953 22587 10011 22593
rect 6972 22528 7788 22556
rect 6972 22516 6978 22528
rect 8202 22516 8208 22568
rect 8260 22556 8266 22568
rect 8570 22556 8576 22568
rect 8260 22528 8576 22556
rect 8260 22516 8266 22528
rect 8570 22516 8576 22528
rect 8628 22516 8634 22568
rect 9125 22559 9183 22565
rect 9125 22525 9137 22559
rect 9171 22556 9183 22559
rect 9876 22556 9904 22587
rect 10318 22584 10324 22596
rect 10376 22584 10382 22636
rect 10597 22627 10655 22633
rect 10597 22593 10609 22627
rect 10643 22593 10655 22627
rect 10597 22587 10655 22593
rect 10781 22627 10839 22633
rect 10781 22593 10793 22627
rect 10827 22624 10839 22627
rect 10827 22596 11008 22624
rect 10827 22593 10839 22596
rect 10781 22587 10839 22593
rect 10226 22556 10232 22568
rect 9171 22528 10232 22556
rect 9171 22525 9183 22528
rect 9125 22519 9183 22525
rect 10226 22516 10232 22528
rect 10284 22556 10290 22568
rect 10410 22556 10416 22568
rect 10284 22528 10416 22556
rect 10284 22516 10290 22528
rect 10410 22516 10416 22528
rect 10468 22516 10474 22568
rect 10612 22556 10640 22587
rect 10870 22556 10876 22568
rect 10612 22528 10876 22556
rect 10870 22516 10876 22528
rect 10928 22516 10934 22568
rect 5442 22488 5448 22500
rect 5092 22460 5448 22488
rect 5442 22448 5448 22460
rect 5500 22448 5506 22500
rect 7926 22448 7932 22500
rect 7984 22488 7990 22500
rect 7984 22460 8800 22488
rect 7984 22448 7990 22460
rect 2317 22423 2375 22429
rect 2317 22389 2329 22423
rect 2363 22420 2375 22423
rect 2406 22420 2412 22432
rect 2363 22392 2412 22420
rect 2363 22389 2375 22392
rect 2317 22383 2375 22389
rect 2406 22380 2412 22392
rect 2464 22380 2470 22432
rect 4433 22423 4491 22429
rect 4433 22389 4445 22423
rect 4479 22420 4491 22423
rect 4798 22420 4804 22432
rect 4479 22392 4804 22420
rect 4479 22389 4491 22392
rect 4433 22383 4491 22389
rect 4798 22380 4804 22392
rect 4856 22380 4862 22432
rect 4890 22380 4896 22432
rect 4948 22420 4954 22432
rect 5258 22420 5264 22432
rect 4948 22392 5264 22420
rect 4948 22380 4954 22392
rect 5258 22380 5264 22392
rect 5316 22420 5322 22432
rect 5353 22423 5411 22429
rect 5353 22420 5365 22423
rect 5316 22392 5365 22420
rect 5316 22380 5322 22392
rect 5353 22389 5365 22392
rect 5399 22389 5411 22423
rect 6546 22420 6552 22432
rect 6507 22392 6552 22420
rect 5353 22383 5411 22389
rect 6546 22380 6552 22392
rect 6604 22380 6610 22432
rect 7006 22380 7012 22432
rect 7064 22420 7070 22432
rect 7101 22423 7159 22429
rect 7101 22420 7113 22423
rect 7064 22392 7113 22420
rect 7064 22380 7070 22392
rect 7101 22389 7113 22392
rect 7147 22389 7159 22423
rect 7101 22383 7159 22389
rect 7466 22380 7472 22432
rect 7524 22420 7530 22432
rect 8110 22420 8116 22432
rect 7524 22392 8116 22420
rect 7524 22380 7530 22392
rect 8110 22380 8116 22392
rect 8168 22380 8174 22432
rect 8662 22420 8668 22432
rect 8623 22392 8668 22420
rect 8662 22380 8668 22392
rect 8720 22380 8726 22432
rect 8772 22420 8800 22460
rect 9490 22448 9496 22500
rect 9548 22488 9554 22500
rect 10689 22491 10747 22497
rect 10689 22488 10701 22491
rect 9548 22460 10701 22488
rect 9548 22448 9554 22460
rect 10689 22457 10701 22460
rect 10735 22457 10747 22491
rect 10689 22451 10747 22457
rect 10980 22420 11008 22596
rect 11330 22584 11336 22636
rect 11388 22624 11394 22636
rect 12066 22624 12072 22636
rect 11388 22596 12072 22624
rect 11388 22584 11394 22596
rect 12066 22584 12072 22596
rect 12124 22624 12130 22636
rect 12360 22633 12388 22664
rect 13538 22652 13544 22704
rect 13596 22692 13602 22704
rect 15105 22695 15163 22701
rect 15105 22692 15117 22695
rect 13596 22664 15117 22692
rect 13596 22652 13602 22664
rect 15105 22661 15117 22664
rect 15151 22692 15163 22695
rect 15194 22692 15200 22704
rect 15151 22664 15200 22692
rect 15151 22661 15163 22664
rect 15105 22655 15163 22661
rect 15194 22652 15200 22664
rect 15252 22652 15258 22704
rect 15289 22695 15347 22701
rect 15289 22661 15301 22695
rect 15335 22692 15347 22695
rect 15470 22692 15476 22704
rect 15335 22664 15476 22692
rect 15335 22661 15347 22664
rect 15289 22655 15347 22661
rect 15470 22652 15476 22664
rect 15528 22692 15534 22704
rect 19702 22692 19708 22704
rect 15528 22664 19708 22692
rect 15528 22652 15534 22664
rect 12253 22627 12311 22633
rect 12253 22624 12265 22627
rect 12124 22596 12265 22624
rect 12124 22584 12130 22596
rect 12253 22593 12265 22596
rect 12299 22593 12311 22627
rect 12253 22587 12311 22593
rect 12345 22627 12403 22633
rect 12345 22593 12357 22627
rect 12391 22624 12403 22627
rect 12526 22624 12532 22636
rect 12391 22596 12532 22624
rect 12391 22593 12403 22596
rect 12345 22587 12403 22593
rect 12526 22584 12532 22596
rect 12584 22584 12590 22636
rect 14090 22624 14096 22636
rect 14051 22596 14096 22624
rect 14090 22584 14096 22596
rect 14148 22584 14154 22636
rect 14182 22584 14188 22636
rect 14240 22624 14246 22636
rect 14458 22624 14464 22636
rect 14240 22596 14464 22624
rect 14240 22584 14246 22596
rect 14458 22584 14464 22596
rect 14516 22584 14522 22636
rect 15654 22584 15660 22636
rect 15712 22624 15718 22636
rect 16040 22633 16068 22664
rect 19702 22652 19708 22664
rect 19760 22692 19766 22704
rect 20346 22692 20352 22704
rect 19760 22664 20352 22692
rect 19760 22652 19766 22664
rect 20346 22652 20352 22664
rect 20404 22652 20410 22704
rect 22186 22652 22192 22704
rect 22244 22692 22250 22704
rect 22646 22692 22652 22704
rect 22244 22664 22652 22692
rect 22244 22652 22250 22664
rect 22646 22652 22652 22664
rect 22704 22652 22710 22704
rect 25314 22652 25320 22704
rect 25372 22692 25378 22704
rect 25593 22695 25651 22701
rect 25593 22692 25605 22695
rect 25372 22664 25605 22692
rect 25372 22652 25378 22664
rect 25593 22661 25605 22664
rect 25639 22661 25651 22695
rect 25593 22655 25651 22661
rect 15749 22627 15807 22633
rect 15749 22624 15761 22627
rect 15712 22596 15761 22624
rect 15712 22584 15718 22596
rect 15749 22593 15761 22596
rect 15795 22593 15807 22627
rect 15749 22587 15807 22593
rect 16025 22627 16083 22633
rect 16025 22593 16037 22627
rect 16071 22593 16083 22627
rect 16025 22587 16083 22593
rect 16853 22627 16911 22633
rect 16853 22593 16865 22627
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 12158 22556 12164 22568
rect 12119 22528 12164 22556
rect 12158 22516 12164 22528
rect 12216 22516 12222 22568
rect 12434 22556 12440 22568
rect 12395 22528 12440 22556
rect 12434 22516 12440 22528
rect 12492 22516 12498 22568
rect 12986 22556 12992 22568
rect 12947 22528 12992 22556
rect 12986 22516 12992 22528
rect 13044 22516 13050 22568
rect 16482 22516 16488 22568
rect 16540 22556 16546 22568
rect 16868 22556 16896 22587
rect 17954 22584 17960 22636
rect 18012 22624 18018 22636
rect 18230 22624 18236 22636
rect 18012 22596 18236 22624
rect 18012 22584 18018 22596
rect 18230 22584 18236 22596
rect 18288 22624 18294 22636
rect 18325 22627 18383 22633
rect 18325 22624 18337 22627
rect 18288 22596 18337 22624
rect 18288 22584 18294 22596
rect 18325 22593 18337 22596
rect 18371 22593 18383 22627
rect 18325 22587 18383 22593
rect 18785 22627 18843 22633
rect 18785 22593 18797 22627
rect 18831 22624 18843 22627
rect 19426 22624 19432 22636
rect 18831 22596 19432 22624
rect 18831 22593 18843 22596
rect 18785 22587 18843 22593
rect 19426 22584 19432 22596
rect 19484 22624 19490 22636
rect 19613 22627 19671 22633
rect 19613 22624 19625 22627
rect 19484 22596 19625 22624
rect 19484 22584 19490 22596
rect 19613 22593 19625 22596
rect 19659 22624 19671 22627
rect 20717 22627 20775 22633
rect 19659 22596 20392 22624
rect 19659 22593 19671 22596
rect 19613 22587 19671 22593
rect 20364 22568 20392 22596
rect 20717 22593 20729 22627
rect 20763 22624 20775 22627
rect 21542 22624 21548 22636
rect 20763 22596 21548 22624
rect 20763 22593 20775 22596
rect 20717 22587 20775 22593
rect 21542 22584 21548 22596
rect 21600 22584 21606 22636
rect 22370 22584 22376 22636
rect 22428 22624 22434 22636
rect 22554 22624 22560 22636
rect 22428 22596 22560 22624
rect 22428 22584 22434 22596
rect 22554 22584 22560 22596
rect 22612 22584 22618 22636
rect 23661 22627 23719 22633
rect 23661 22593 23673 22627
rect 23707 22624 23719 22627
rect 23842 22624 23848 22636
rect 23707 22596 23848 22624
rect 23707 22593 23719 22596
rect 23661 22587 23719 22593
rect 23842 22584 23848 22596
rect 23900 22584 23906 22636
rect 27154 22624 27160 22636
rect 27115 22596 27160 22624
rect 27154 22584 27160 22596
rect 27212 22584 27218 22636
rect 16540 22528 16896 22556
rect 16945 22559 17003 22565
rect 16540 22516 16546 22528
rect 16945 22525 16957 22559
rect 16991 22525 17003 22559
rect 18877 22559 18935 22565
rect 18877 22556 18889 22559
rect 16945 22519 17003 22525
rect 18156 22528 18889 22556
rect 11977 22491 12035 22497
rect 11977 22457 11989 22491
rect 12023 22457 12035 22491
rect 13265 22491 13323 22497
rect 13265 22488 13277 22491
rect 11977 22451 12035 22457
rect 12406 22460 13277 22488
rect 8772 22392 11008 22420
rect 11992 22420 12020 22451
rect 12406 22420 12434 22460
rect 13265 22457 13277 22460
rect 13311 22457 13323 22491
rect 13265 22451 13323 22457
rect 13449 22491 13507 22497
rect 13449 22457 13461 22491
rect 13495 22488 13507 22491
rect 16022 22488 16028 22500
rect 13495 22460 16028 22488
rect 13495 22457 13507 22460
rect 13449 22451 13507 22457
rect 16022 22448 16028 22460
rect 16080 22448 16086 22500
rect 11992 22392 12434 22420
rect 13998 22380 14004 22432
rect 14056 22420 14062 22432
rect 14369 22423 14427 22429
rect 14369 22420 14381 22423
rect 14056 22392 14381 22420
rect 14056 22380 14062 22392
rect 14369 22389 14381 22392
rect 14415 22389 14427 22423
rect 14369 22383 14427 22389
rect 16482 22380 16488 22432
rect 16540 22420 16546 22432
rect 16960 22420 16988 22519
rect 18156 22497 18184 22528
rect 18877 22525 18889 22528
rect 18923 22556 18935 22559
rect 19705 22559 19763 22565
rect 19705 22556 19717 22559
rect 18923 22528 19717 22556
rect 18923 22525 18935 22528
rect 18877 22519 18935 22525
rect 19705 22525 19717 22528
rect 19751 22556 19763 22559
rect 19794 22556 19800 22568
rect 19751 22528 19800 22556
rect 19751 22525 19763 22528
rect 19705 22519 19763 22525
rect 19794 22516 19800 22528
rect 19852 22516 19858 22568
rect 20346 22516 20352 22568
rect 20404 22516 20410 22568
rect 20441 22559 20499 22565
rect 20441 22525 20453 22559
rect 20487 22556 20499 22559
rect 20530 22556 20536 22568
rect 20487 22528 20536 22556
rect 20487 22525 20499 22528
rect 20441 22519 20499 22525
rect 20530 22516 20536 22528
rect 20588 22516 20594 22568
rect 20806 22516 20812 22568
rect 20864 22556 20870 22568
rect 22189 22559 22247 22565
rect 22189 22556 22201 22559
rect 20864 22528 22201 22556
rect 20864 22516 20870 22528
rect 22189 22525 22201 22528
rect 22235 22525 22247 22559
rect 22189 22519 22247 22525
rect 22465 22559 22523 22565
rect 22465 22525 22477 22559
rect 22511 22556 22523 22559
rect 23382 22556 23388 22568
rect 22511 22528 23388 22556
rect 22511 22525 22523 22528
rect 22465 22519 22523 22525
rect 23382 22516 23388 22528
rect 23440 22516 23446 22568
rect 23937 22559 23995 22565
rect 23937 22525 23949 22559
rect 23983 22556 23995 22559
rect 25038 22556 25044 22568
rect 23983 22528 25044 22556
rect 23983 22525 23995 22528
rect 23937 22519 23995 22525
rect 25038 22516 25044 22528
rect 25096 22516 25102 22568
rect 25777 22559 25835 22565
rect 25777 22525 25789 22559
rect 25823 22556 25835 22559
rect 25866 22556 25872 22568
rect 25823 22528 25872 22556
rect 25823 22525 25835 22528
rect 25777 22519 25835 22525
rect 25866 22516 25872 22528
rect 25924 22516 25930 22568
rect 26142 22516 26148 22568
rect 26200 22556 26206 22568
rect 26786 22556 26792 22568
rect 26200 22528 26792 22556
rect 26200 22516 26206 22528
rect 26786 22516 26792 22528
rect 26844 22556 26850 22568
rect 26973 22559 27031 22565
rect 26973 22556 26985 22559
rect 26844 22528 26985 22556
rect 26844 22516 26850 22528
rect 26973 22525 26985 22528
rect 27019 22525 27031 22559
rect 26973 22519 27031 22525
rect 18141 22491 18199 22497
rect 18141 22457 18153 22491
rect 18187 22457 18199 22491
rect 19153 22491 19211 22497
rect 18141 22451 18199 22457
rect 18800 22460 19104 22488
rect 16540 22392 16988 22420
rect 17129 22423 17187 22429
rect 16540 22380 16546 22392
rect 17129 22389 17141 22423
rect 17175 22420 17187 22423
rect 18800 22420 18828 22460
rect 18966 22420 18972 22432
rect 17175 22392 18828 22420
rect 18927 22392 18972 22420
rect 17175 22389 17187 22392
rect 17129 22383 17187 22389
rect 18966 22380 18972 22392
rect 19024 22380 19030 22432
rect 19076 22420 19104 22460
rect 19153 22457 19165 22491
rect 19199 22488 19211 22491
rect 19518 22488 19524 22500
rect 19199 22460 19524 22488
rect 19199 22457 19211 22460
rect 19153 22451 19211 22457
rect 19518 22448 19524 22460
rect 19576 22448 19582 22500
rect 20898 22448 20904 22500
rect 20956 22488 20962 22500
rect 20956 22460 21772 22488
rect 20956 22448 20962 22460
rect 19613 22423 19671 22429
rect 19613 22420 19625 22423
rect 19076 22392 19625 22420
rect 19613 22389 19625 22392
rect 19659 22420 19671 22423
rect 21634 22420 21640 22432
rect 19659 22392 21640 22420
rect 19659 22389 19671 22392
rect 19613 22383 19671 22389
rect 21634 22380 21640 22392
rect 21692 22380 21698 22432
rect 21744 22420 21772 22460
rect 22554 22448 22560 22500
rect 22612 22488 22618 22500
rect 23106 22488 23112 22500
rect 22612 22460 23112 22488
rect 22612 22448 22618 22460
rect 23106 22448 23112 22460
rect 23164 22448 23170 22500
rect 23290 22420 23296 22432
rect 21744 22392 23296 22420
rect 23290 22380 23296 22392
rect 23348 22380 23354 22432
rect 25133 22423 25191 22429
rect 25133 22389 25145 22423
rect 25179 22420 25191 22423
rect 25866 22420 25872 22432
rect 25179 22392 25872 22420
rect 25179 22389 25191 22392
rect 25133 22383 25191 22389
rect 25866 22380 25872 22392
rect 25924 22380 25930 22432
rect 1104 22330 28060 22352
rect 1104 22278 5442 22330
rect 5494 22278 5506 22330
rect 5558 22278 5570 22330
rect 5622 22278 5634 22330
rect 5686 22278 5698 22330
rect 5750 22278 14428 22330
rect 14480 22278 14492 22330
rect 14544 22278 14556 22330
rect 14608 22278 14620 22330
rect 14672 22278 14684 22330
rect 14736 22278 23413 22330
rect 23465 22278 23477 22330
rect 23529 22278 23541 22330
rect 23593 22278 23605 22330
rect 23657 22278 23669 22330
rect 23721 22278 28060 22330
rect 1104 22256 28060 22278
rect 4062 22176 4068 22228
rect 4120 22216 4126 22228
rect 4120 22188 4476 22216
rect 4120 22176 4126 22188
rect 3142 22108 3148 22160
rect 3200 22148 3206 22160
rect 3200 22120 4108 22148
rect 3200 22108 3206 22120
rect 4080 22080 4108 22120
rect 4448 22080 4476 22188
rect 4982 22176 4988 22228
rect 5040 22216 5046 22228
rect 5077 22219 5135 22225
rect 5077 22216 5089 22219
rect 5040 22188 5089 22216
rect 5040 22176 5046 22188
rect 5077 22185 5089 22188
rect 5123 22185 5135 22219
rect 8202 22216 8208 22228
rect 5077 22179 5135 22185
rect 5210 22188 5580 22216
rect 4525 22151 4583 22157
rect 4525 22117 4537 22151
rect 4571 22148 4583 22151
rect 5210 22148 5238 22188
rect 5552 22160 5580 22188
rect 6288 22188 8208 22216
rect 4571 22120 5238 22148
rect 4571 22117 4583 22120
rect 4525 22111 4583 22117
rect 5534 22108 5540 22160
rect 5592 22108 5598 22160
rect 6086 22080 6092 22092
rect 1964 22052 3372 22080
rect 4080 22052 4384 22080
rect 4448 22052 5120 22080
rect 1964 22021 1992 22052
rect 3344 22021 3372 22052
rect 1949 22015 2007 22021
rect 1949 21981 1961 22015
rect 1995 21981 2007 22015
rect 1949 21975 2007 21981
rect 2593 22015 2651 22021
rect 2593 21981 2605 22015
rect 2639 22012 2651 22015
rect 3329 22015 3387 22021
rect 2639 21984 3004 22012
rect 2639 21981 2651 21984
rect 2593 21975 2651 21981
rect 1765 21879 1823 21885
rect 1765 21845 1777 21879
rect 1811 21876 1823 21879
rect 2314 21876 2320 21888
rect 1811 21848 2320 21876
rect 1811 21845 1823 21848
rect 1765 21839 1823 21845
rect 2314 21836 2320 21848
rect 2372 21836 2378 21888
rect 2409 21879 2467 21885
rect 2409 21845 2421 21879
rect 2455 21876 2467 21879
rect 2682 21876 2688 21888
rect 2455 21848 2688 21876
rect 2455 21845 2467 21848
rect 2409 21839 2467 21845
rect 2682 21836 2688 21848
rect 2740 21836 2746 21888
rect 2976 21885 3004 21984
rect 3329 21981 3341 22015
rect 3375 22012 3387 22015
rect 3418 22012 3424 22024
rect 3375 21984 3424 22012
rect 3375 21981 3387 21984
rect 3329 21975 3387 21981
rect 3418 21972 3424 21984
rect 3476 21972 3482 22024
rect 3605 22015 3663 22021
rect 3605 21981 3617 22015
rect 3651 22012 3663 22015
rect 3970 22012 3976 22024
rect 3651 21984 3976 22012
rect 3651 21981 3663 21984
rect 3605 21975 3663 21981
rect 3970 21972 3976 21984
rect 4028 21972 4034 22024
rect 4246 22012 4252 22024
rect 4207 21984 4252 22012
rect 4246 21972 4252 21984
rect 4304 21972 4310 22024
rect 4356 22021 4384 22052
rect 4341 22015 4399 22021
rect 4341 21981 4353 22015
rect 4387 21981 4399 22015
rect 4614 22012 4620 22024
rect 4575 21984 4620 22012
rect 4341 21975 4399 21981
rect 4614 21972 4620 21984
rect 4672 21972 4678 22024
rect 5092 22021 5120 22052
rect 5184 22052 6092 22080
rect 5184 22021 5212 22052
rect 6086 22040 6092 22052
rect 6144 22040 6150 22092
rect 5077 22015 5135 22021
rect 5077 21981 5089 22015
rect 5123 21981 5135 22015
rect 5077 21975 5135 21981
rect 5169 22015 5227 22021
rect 5169 21981 5181 22015
rect 5215 21981 5227 22015
rect 5350 22012 5356 22024
rect 5311 21984 5356 22012
rect 5169 21975 5227 21981
rect 5350 21972 5356 21984
rect 5408 21972 5414 22024
rect 5534 21972 5540 22024
rect 5592 22012 5598 22024
rect 6288 22012 6316 22188
rect 8202 22176 8208 22188
rect 8260 22176 8266 22228
rect 8297 22219 8355 22225
rect 8297 22185 8309 22219
rect 8343 22216 8355 22219
rect 8662 22216 8668 22228
rect 8343 22188 8668 22216
rect 8343 22185 8355 22188
rect 8297 22179 8355 22185
rect 8662 22176 8668 22188
rect 8720 22176 8726 22228
rect 9125 22219 9183 22225
rect 9125 22185 9137 22219
rect 9171 22216 9183 22219
rect 11609 22219 11667 22225
rect 9171 22188 10640 22216
rect 9171 22185 9183 22188
rect 9125 22179 9183 22185
rect 7466 22148 7472 22160
rect 7208 22120 7472 22148
rect 7208 22089 7236 22120
rect 7466 22108 7472 22120
rect 7524 22108 7530 22160
rect 7929 22151 7987 22157
rect 7929 22117 7941 22151
rect 7975 22148 7987 22151
rect 9033 22151 9091 22157
rect 9033 22148 9045 22151
rect 7975 22120 9045 22148
rect 7975 22117 7987 22120
rect 7929 22111 7987 22117
rect 9033 22117 9045 22120
rect 9079 22117 9091 22151
rect 10134 22148 10140 22160
rect 9033 22111 9091 22117
rect 9968 22120 10140 22148
rect 7193 22083 7251 22089
rect 5592 21984 6316 22012
rect 6748 22052 7144 22080
rect 5592 21972 5598 21984
rect 4632 21944 4660 21972
rect 4982 21944 4988 21956
rect 4632 21916 4988 21944
rect 4982 21904 4988 21916
rect 5040 21944 5046 21956
rect 5445 21947 5503 21953
rect 5445 21944 5457 21947
rect 5040 21916 5457 21944
rect 5040 21904 5046 21916
rect 5445 21913 5457 21916
rect 5491 21913 5503 21947
rect 5445 21907 5503 21913
rect 5902 21904 5908 21956
rect 5960 21944 5966 21956
rect 6748 21944 6776 22052
rect 6825 22015 6883 22021
rect 6825 21981 6837 22015
rect 6871 21981 6883 22015
rect 6825 21975 6883 21981
rect 5960 21916 6776 21944
rect 5960 21904 5966 21916
rect 6840 21888 6868 21975
rect 6914 21972 6920 22024
rect 6972 22012 6978 22024
rect 7116 22012 7144 22052
rect 7193 22049 7205 22083
rect 7239 22049 7251 22083
rect 7193 22043 7251 22049
rect 7374 22040 7380 22092
rect 7432 22080 7438 22092
rect 9217 22083 9275 22089
rect 9217 22080 9229 22083
rect 7432 22052 9229 22080
rect 7432 22040 7438 22052
rect 9217 22049 9229 22052
rect 9263 22049 9275 22083
rect 9217 22043 9275 22049
rect 9766 22040 9772 22092
rect 9824 22080 9830 22092
rect 9968 22089 9996 22120
rect 10134 22108 10140 22120
rect 10192 22108 10198 22160
rect 9953 22083 10011 22089
rect 9824 22052 9904 22080
rect 9824 22040 9830 22052
rect 6972 21984 7017 22012
rect 7116 21984 7604 22012
rect 6972 21972 6978 21984
rect 7282 21944 7288 21956
rect 7243 21916 7288 21944
rect 7282 21904 7288 21916
rect 7340 21904 7346 21956
rect 7576 21944 7604 21984
rect 7650 21972 7656 22024
rect 7708 22012 7714 22024
rect 8113 22015 8171 22021
rect 8113 22012 8125 22015
rect 7708 21984 8125 22012
rect 7708 21972 7714 21984
rect 8113 21981 8125 21984
rect 8159 21981 8171 22015
rect 8294 22014 8300 22024
rect 8266 22012 8300 22014
rect 8113 21975 8171 21981
rect 8220 21984 8300 22012
rect 8220 21944 8248 21984
rect 8294 21972 8300 21984
rect 8352 21972 8358 22024
rect 8389 22015 8447 22021
rect 8389 21981 8401 22015
rect 8435 21981 8447 22015
rect 8938 22012 8944 22024
rect 8899 21984 8944 22012
rect 8389 21975 8447 21981
rect 7576 21916 8248 21944
rect 8404 21944 8432 21975
rect 8938 21972 8944 21984
rect 8996 21972 9002 22024
rect 9674 22012 9680 22024
rect 9635 21984 9680 22012
rect 9674 21972 9680 21984
rect 9732 21972 9738 22024
rect 9876 22021 9904 22052
rect 9953 22049 9965 22083
rect 9999 22049 10011 22083
rect 9953 22043 10011 22049
rect 10045 22083 10103 22089
rect 10045 22049 10057 22083
rect 10091 22080 10103 22083
rect 10318 22080 10324 22092
rect 10091 22052 10324 22080
rect 10091 22049 10103 22052
rect 10045 22043 10103 22049
rect 10318 22040 10324 22052
rect 10376 22040 10382 22092
rect 10410 22040 10416 22092
rect 10468 22080 10474 22092
rect 10468 22052 10513 22080
rect 10468 22040 10474 22052
rect 10612 22024 10640 22188
rect 11609 22185 11621 22219
rect 11655 22216 11667 22219
rect 12986 22216 12992 22228
rect 11655 22188 12992 22216
rect 11655 22185 11667 22188
rect 11609 22179 11667 22185
rect 12986 22176 12992 22188
rect 13044 22176 13050 22228
rect 13998 22176 14004 22228
rect 14056 22176 14062 22228
rect 14182 22176 14188 22228
rect 14240 22216 14246 22228
rect 14240 22188 14495 22216
rect 14240 22176 14246 22188
rect 12158 22108 12164 22160
rect 12216 22148 12222 22160
rect 12216 22120 12296 22148
rect 12216 22108 12222 22120
rect 11606 22040 11612 22092
rect 11664 22080 11670 22092
rect 11882 22080 11888 22092
rect 11664 22052 11888 22080
rect 11664 22040 11670 22052
rect 11882 22040 11888 22052
rect 11940 22040 11946 22092
rect 12268 22089 12296 22120
rect 12253 22083 12311 22089
rect 12253 22049 12265 22083
rect 12299 22080 12311 22083
rect 14016 22080 14044 22176
rect 14090 22108 14096 22160
rect 14148 22148 14154 22160
rect 14366 22148 14372 22160
rect 14148 22120 14372 22148
rect 14148 22108 14154 22120
rect 14366 22108 14372 22120
rect 14424 22108 14430 22160
rect 14467 22080 14495 22188
rect 18966 22176 18972 22228
rect 19024 22216 19030 22228
rect 19610 22216 19616 22228
rect 19024 22188 19616 22216
rect 19024 22176 19030 22188
rect 19610 22176 19616 22188
rect 19668 22176 19674 22228
rect 20530 22216 20536 22228
rect 19720 22188 20536 22216
rect 18141 22151 18199 22157
rect 18141 22117 18153 22151
rect 18187 22148 18199 22151
rect 18322 22148 18328 22160
rect 18187 22120 18328 22148
rect 18187 22117 18199 22120
rect 18141 22111 18199 22117
rect 18322 22108 18328 22120
rect 18380 22148 18386 22160
rect 19720 22148 19748 22188
rect 20530 22176 20536 22188
rect 20588 22176 20594 22228
rect 25682 22176 25688 22228
rect 25740 22216 25746 22228
rect 26142 22216 26148 22228
rect 25740 22188 26148 22216
rect 25740 22176 25746 22188
rect 26142 22176 26148 22188
rect 26200 22176 26206 22228
rect 26237 22219 26295 22225
rect 26237 22185 26249 22219
rect 26283 22216 26295 22219
rect 27154 22216 27160 22228
rect 26283 22188 27160 22216
rect 26283 22185 26295 22188
rect 26237 22179 26295 22185
rect 27154 22176 27160 22188
rect 27212 22176 27218 22228
rect 18380 22120 19748 22148
rect 18380 22108 18386 22120
rect 23474 22108 23480 22160
rect 23532 22148 23538 22160
rect 23842 22148 23848 22160
rect 23532 22120 23848 22148
rect 23532 22108 23538 22120
rect 23842 22108 23848 22120
rect 23900 22108 23906 22160
rect 26050 22108 26056 22160
rect 26108 22148 26114 22160
rect 26108 22120 26188 22148
rect 26108 22108 26114 22120
rect 15102 22080 15108 22092
rect 12299 22052 12333 22080
rect 14016 22052 14136 22080
rect 12299 22049 12311 22052
rect 12253 22043 12311 22049
rect 14108 22024 14136 22052
rect 14200 22052 15108 22080
rect 9861 22015 9919 22021
rect 9861 21981 9873 22015
rect 9907 21981 9919 22015
rect 10226 22012 10232 22024
rect 10187 21984 10232 22012
rect 9861 21975 9919 21981
rect 10226 21972 10232 21984
rect 10284 21972 10290 22024
rect 10594 21972 10600 22024
rect 10652 21972 10658 22024
rect 11793 22015 11851 22021
rect 11793 21981 11805 22015
rect 11839 21981 11851 22015
rect 11793 21975 11851 21981
rect 8662 21944 8668 21956
rect 8404 21916 8668 21944
rect 8662 21904 8668 21916
rect 8720 21904 8726 21956
rect 10962 21944 10968 21956
rect 10923 21916 10968 21944
rect 10962 21904 10968 21916
rect 11020 21904 11026 21956
rect 11808 21944 11836 21975
rect 12066 21972 12072 22024
rect 12124 22012 12130 22024
rect 12161 22015 12219 22021
rect 12161 22012 12173 22015
rect 12124 21984 12173 22012
rect 12124 21972 12130 21984
rect 12161 21981 12173 21984
rect 12207 21981 12219 22015
rect 12161 21975 12219 21981
rect 12713 22015 12771 22021
rect 12713 21981 12725 22015
rect 12759 22012 12771 22015
rect 12802 22012 12808 22024
rect 12759 21984 12808 22012
rect 12759 21981 12771 21984
rect 12713 21975 12771 21981
rect 12802 21972 12808 21984
rect 12860 21972 12866 22024
rect 12897 22015 12955 22021
rect 12897 21981 12909 22015
rect 12943 21981 12955 22015
rect 12897 21975 12955 21981
rect 13541 22015 13599 22021
rect 13541 21981 13553 22015
rect 13587 22012 13599 22015
rect 13906 22012 13912 22024
rect 13587 21984 13912 22012
rect 13587 21981 13599 21984
rect 13541 21975 13599 21981
rect 12526 21944 12532 21956
rect 11808 21916 12532 21944
rect 12526 21904 12532 21916
rect 12584 21944 12590 21956
rect 12912 21944 12940 21975
rect 13906 21972 13912 21984
rect 13964 21972 13970 22024
rect 14090 21972 14096 22024
rect 14148 21972 14154 22024
rect 14200 22021 14228 22052
rect 15102 22040 15108 22052
rect 15160 22040 15166 22092
rect 15286 22040 15292 22092
rect 15344 22080 15350 22092
rect 15838 22080 15844 22092
rect 15344 22052 15844 22080
rect 15344 22040 15350 22052
rect 15838 22040 15844 22052
rect 15896 22040 15902 22092
rect 16482 22040 16488 22092
rect 16540 22080 16546 22092
rect 16577 22083 16635 22089
rect 16577 22080 16589 22083
rect 16540 22052 16589 22080
rect 16540 22040 16546 22052
rect 16577 22049 16589 22052
rect 16623 22080 16635 22083
rect 17681 22083 17739 22089
rect 17681 22080 17693 22083
rect 16623 22052 17693 22080
rect 16623 22049 16635 22052
rect 16577 22043 16635 22049
rect 17681 22049 17693 22052
rect 17727 22080 17739 22083
rect 17862 22080 17868 22092
rect 17727 22052 17868 22080
rect 17727 22049 17739 22052
rect 17681 22043 17739 22049
rect 17862 22040 17868 22052
rect 17920 22040 17926 22092
rect 20165 22083 20223 22089
rect 20165 22049 20177 22083
rect 20211 22080 20223 22083
rect 20898 22080 20904 22092
rect 20211 22052 20904 22080
rect 20211 22049 20223 22052
rect 20165 22043 20223 22049
rect 20898 22040 20904 22052
rect 20956 22040 20962 22092
rect 21913 22083 21971 22089
rect 21913 22049 21925 22083
rect 21959 22080 21971 22083
rect 22002 22080 22008 22092
rect 21959 22052 22008 22080
rect 21959 22049 21971 22052
rect 21913 22043 21971 22049
rect 22002 22040 22008 22052
rect 22060 22040 22066 22092
rect 23382 22040 23388 22092
rect 23440 22080 23446 22092
rect 23661 22083 23719 22089
rect 23661 22080 23673 22083
rect 23440 22052 23673 22080
rect 23440 22040 23446 22052
rect 23661 22049 23673 22052
rect 23707 22049 23719 22083
rect 25041 22083 25099 22089
rect 25041 22080 25053 22083
rect 23661 22043 23719 22049
rect 23768 22052 25053 22080
rect 14185 22015 14243 22021
rect 14185 21981 14197 22015
rect 14231 21981 14243 22015
rect 14185 21975 14243 21981
rect 14366 21972 14372 22024
rect 14424 22012 14430 22024
rect 14734 22012 14740 22024
rect 14424 21984 14740 22012
rect 14424 21972 14430 21984
rect 14734 21972 14740 21984
rect 14792 21972 14798 22024
rect 16298 21972 16304 22024
rect 16356 22012 16362 22024
rect 17773 22015 17831 22021
rect 17773 22012 17785 22015
rect 16356 21984 17785 22012
rect 16356 21972 16362 21984
rect 17773 21981 17785 21984
rect 17819 22012 17831 22015
rect 17954 22012 17960 22024
rect 17819 21984 17960 22012
rect 17819 21981 17831 21984
rect 17773 21975 17831 21981
rect 17954 21972 17960 21984
rect 18012 21972 18018 22024
rect 18230 21972 18236 22024
rect 18288 22012 18294 22024
rect 19245 22015 19303 22021
rect 19245 22012 19257 22015
rect 18288 21984 19257 22012
rect 18288 21972 18294 21984
rect 19245 21981 19257 21984
rect 19291 21981 19303 22015
rect 19429 22015 19487 22021
rect 19429 22006 19441 22015
rect 19245 21975 19303 21981
rect 19352 21981 19441 22006
rect 19475 21981 19487 22015
rect 19886 22012 19892 22024
rect 19847 21984 19892 22012
rect 19352 21978 19487 21981
rect 14277 21947 14335 21953
rect 12584 21916 14219 21944
rect 12584 21904 12590 21916
rect 2961 21879 3019 21885
rect 2961 21845 2973 21879
rect 3007 21876 3019 21879
rect 3234 21876 3240 21888
rect 3007 21848 3240 21876
rect 3007 21845 3019 21848
rect 2961 21839 3019 21845
rect 3234 21836 3240 21848
rect 3292 21836 3298 21888
rect 3421 21879 3479 21885
rect 3421 21845 3433 21879
rect 3467 21876 3479 21879
rect 3510 21876 3516 21888
rect 3467 21848 3516 21876
rect 3467 21845 3479 21848
rect 3421 21839 3479 21845
rect 3510 21836 3516 21848
rect 3568 21836 3574 21888
rect 4065 21879 4123 21885
rect 4065 21845 4077 21879
rect 4111 21876 4123 21879
rect 5074 21876 5080 21888
rect 4111 21848 5080 21876
rect 4111 21845 4123 21848
rect 4065 21839 4123 21845
rect 5074 21836 5080 21848
rect 5132 21836 5138 21888
rect 6638 21876 6644 21888
rect 6599 21848 6644 21876
rect 6638 21836 6644 21848
rect 6696 21836 6702 21888
rect 6822 21836 6828 21888
rect 6880 21876 6886 21888
rect 8478 21876 8484 21888
rect 6880 21848 8484 21876
rect 6880 21836 6886 21848
rect 8478 21836 8484 21848
rect 8536 21836 8542 21888
rect 11057 21879 11115 21885
rect 11057 21845 11069 21879
rect 11103 21876 11115 21879
rect 11790 21876 11796 21888
rect 11103 21848 11796 21876
rect 11103 21845 11115 21848
rect 11057 21839 11115 21845
rect 11790 21836 11796 21848
rect 11848 21836 11854 21888
rect 12069 21879 12127 21885
rect 12069 21845 12081 21879
rect 12115 21876 12127 21879
rect 12434 21876 12440 21888
rect 12115 21848 12440 21876
rect 12115 21845 12127 21848
rect 12069 21839 12127 21845
rect 12434 21836 12440 21848
rect 12492 21876 12498 21888
rect 12618 21876 12624 21888
rect 12492 21848 12624 21876
rect 12492 21836 12498 21848
rect 12618 21836 12624 21848
rect 12676 21836 12682 21888
rect 12805 21879 12863 21885
rect 12805 21845 12817 21879
rect 12851 21876 12863 21879
rect 13078 21876 13084 21888
rect 12851 21848 13084 21876
rect 12851 21845 12863 21848
rect 12805 21839 12863 21845
rect 13078 21836 13084 21848
rect 13136 21836 13142 21888
rect 13357 21879 13415 21885
rect 13357 21845 13369 21879
rect 13403 21876 13415 21879
rect 14090 21876 14096 21888
rect 13403 21848 14096 21876
rect 13403 21845 13415 21848
rect 13357 21839 13415 21845
rect 14090 21836 14096 21848
rect 14148 21836 14154 21888
rect 14191 21876 14219 21916
rect 14277 21913 14289 21947
rect 14323 21944 14335 21947
rect 14826 21944 14832 21956
rect 14323 21916 14832 21944
rect 14323 21913 14335 21916
rect 14277 21907 14335 21913
rect 14826 21904 14832 21916
rect 14884 21944 14890 21956
rect 14921 21947 14979 21953
rect 14921 21944 14933 21947
rect 14884 21916 14933 21944
rect 14884 21904 14890 21916
rect 14921 21913 14933 21916
rect 14967 21913 14979 21947
rect 14921 21907 14979 21913
rect 15657 21947 15715 21953
rect 15657 21913 15669 21947
rect 15703 21944 15715 21947
rect 16393 21947 16451 21953
rect 15703 21916 15884 21944
rect 15703 21913 15715 21916
rect 15657 21907 15715 21913
rect 15013 21879 15071 21885
rect 15013 21876 15025 21879
rect 14191 21848 15025 21876
rect 15013 21845 15025 21848
rect 15059 21845 15071 21879
rect 15856 21876 15884 21916
rect 16393 21913 16405 21947
rect 16439 21944 16451 21947
rect 16850 21944 16856 21956
rect 16439 21916 16856 21944
rect 16439 21913 16451 21916
rect 16393 21907 16451 21913
rect 16850 21904 16856 21916
rect 16908 21904 16914 21956
rect 19352 21944 19380 21978
rect 19429 21975 19487 21978
rect 19886 21972 19892 21984
rect 19944 21972 19950 22024
rect 21634 22012 21640 22024
rect 21595 21984 21640 22012
rect 21634 21972 21640 21984
rect 21692 21972 21698 22024
rect 23566 21972 23572 22024
rect 23624 22012 23630 22024
rect 23768 22012 23796 22052
rect 25041 22049 25053 22052
rect 25087 22049 25099 22083
rect 26160 22080 26188 22120
rect 26620 22120 26924 22148
rect 26620 22080 26648 22120
rect 26160 22052 26648 22080
rect 26697 22083 26755 22089
rect 25041 22043 25099 22049
rect 26697 22049 26709 22083
rect 26743 22080 26755 22083
rect 26786 22080 26792 22092
rect 26743 22052 26792 22080
rect 26743 22049 26755 22052
rect 26697 22043 26755 22049
rect 26786 22040 26792 22052
rect 26844 22040 26850 22092
rect 26896 22080 26924 22120
rect 27065 22083 27123 22089
rect 27065 22080 27077 22083
rect 26896 22052 27077 22080
rect 27065 22049 27077 22052
rect 27111 22049 27123 22083
rect 27065 22043 27123 22049
rect 25685 22015 25743 22021
rect 25685 22012 25697 22015
rect 23624 21984 23796 22012
rect 25056 21984 25697 22012
rect 23624 21972 23630 21984
rect 25056 21956 25084 21984
rect 25685 21981 25697 21984
rect 25731 21981 25743 22015
rect 25866 22012 25872 22024
rect 25827 21984 25872 22012
rect 25685 21975 25743 21981
rect 25866 21972 25872 21984
rect 25924 21972 25930 22024
rect 26050 22012 26056 22024
rect 26011 21984 26056 22012
rect 26050 21972 26056 21984
rect 26108 21972 26114 22024
rect 26881 22015 26939 22021
rect 26881 21981 26893 22015
rect 26927 21981 26939 22015
rect 26881 21975 26939 21981
rect 16960 21916 19380 21944
rect 16114 21876 16120 21888
rect 15856 21848 16120 21876
rect 15013 21839 15071 21845
rect 16114 21836 16120 21848
rect 16172 21876 16178 21888
rect 16960 21876 16988 21916
rect 19610 21904 19616 21956
rect 19668 21944 19674 21956
rect 20898 21944 20904 21956
rect 19668 21916 20904 21944
rect 19668 21904 19674 21916
rect 20898 21904 20904 21916
rect 20956 21904 20962 21956
rect 23477 21947 23535 21953
rect 23477 21913 23489 21947
rect 23523 21944 23535 21947
rect 24670 21944 24676 21956
rect 23523 21916 24676 21944
rect 23523 21913 23535 21916
rect 23477 21907 23535 21913
rect 24044 21888 24072 21916
rect 24670 21904 24676 21916
rect 24728 21944 24734 21956
rect 24728 21916 24900 21944
rect 24728 21904 24734 21916
rect 16172 21848 16988 21876
rect 16172 21836 16178 21848
rect 18046 21836 18052 21888
rect 18104 21876 18110 21888
rect 19429 21879 19487 21885
rect 19429 21876 19441 21879
rect 18104 21848 19441 21876
rect 18104 21836 18110 21848
rect 19429 21845 19441 21848
rect 19475 21876 19487 21879
rect 21818 21876 21824 21888
rect 19475 21848 21824 21876
rect 19475 21845 19487 21848
rect 19429 21839 19487 21845
rect 21818 21836 21824 21848
rect 21876 21836 21882 21888
rect 23106 21876 23112 21888
rect 23067 21848 23112 21876
rect 23106 21836 23112 21848
rect 23164 21836 23170 21888
rect 23569 21879 23627 21885
rect 23569 21845 23581 21879
rect 23615 21876 23627 21879
rect 23658 21876 23664 21888
rect 23615 21848 23664 21876
rect 23615 21845 23627 21848
rect 23569 21839 23627 21845
rect 23658 21836 23664 21848
rect 23716 21836 23722 21888
rect 24026 21836 24032 21888
rect 24084 21836 24090 21888
rect 24489 21879 24547 21885
rect 24489 21845 24501 21879
rect 24535 21876 24547 21879
rect 24762 21876 24768 21888
rect 24535 21848 24768 21876
rect 24535 21845 24547 21848
rect 24489 21839 24547 21845
rect 24762 21836 24768 21848
rect 24820 21836 24826 21888
rect 24872 21885 24900 21916
rect 25038 21904 25044 21956
rect 25096 21904 25102 21956
rect 25498 21904 25504 21956
rect 25556 21944 25562 21956
rect 25961 21947 26019 21953
rect 25961 21944 25973 21947
rect 25556 21916 25973 21944
rect 25556 21904 25562 21916
rect 25961 21913 25973 21916
rect 26007 21913 26019 21947
rect 25961 21907 26019 21913
rect 26234 21904 26240 21956
rect 26292 21944 26298 21956
rect 26786 21944 26792 21956
rect 26292 21916 26792 21944
rect 26292 21904 26298 21916
rect 26786 21904 26792 21916
rect 26844 21904 26850 21956
rect 24857 21879 24915 21885
rect 24857 21845 24869 21879
rect 24903 21845 24915 21879
rect 24857 21839 24915 21845
rect 24949 21879 25007 21885
rect 24949 21845 24961 21879
rect 24995 21876 25007 21879
rect 25590 21876 25596 21888
rect 24995 21848 25596 21876
rect 24995 21845 25007 21848
rect 24949 21839 25007 21845
rect 25590 21836 25596 21848
rect 25648 21836 25654 21888
rect 25682 21836 25688 21888
rect 25740 21876 25746 21888
rect 26896 21876 26924 21975
rect 25740 21848 26924 21876
rect 25740 21836 25746 21848
rect 1104 21786 28060 21808
rect 1104 21734 9935 21786
rect 9987 21734 9999 21786
rect 10051 21734 10063 21786
rect 10115 21734 10127 21786
rect 10179 21734 10191 21786
rect 10243 21734 18920 21786
rect 18972 21734 18984 21786
rect 19036 21734 19048 21786
rect 19100 21734 19112 21786
rect 19164 21734 19176 21786
rect 19228 21734 28060 21786
rect 1104 21712 28060 21734
rect 1489 21675 1547 21681
rect 1489 21641 1501 21675
rect 1535 21672 1547 21675
rect 2866 21672 2872 21684
rect 1535 21644 2872 21672
rect 1535 21641 1547 21644
rect 1489 21635 1547 21641
rect 2866 21632 2872 21644
rect 2924 21632 2930 21684
rect 3234 21632 3240 21684
rect 3292 21672 3298 21684
rect 4062 21672 4068 21684
rect 3292 21644 3924 21672
rect 4023 21644 4068 21672
rect 3292 21632 3298 21644
rect 3142 21564 3148 21616
rect 3200 21604 3206 21616
rect 3789 21607 3847 21613
rect 3789 21604 3801 21607
rect 3200 21576 3801 21604
rect 3200 21564 3206 21576
rect 3789 21573 3801 21576
rect 3835 21573 3847 21607
rect 3896 21604 3924 21644
rect 4062 21632 4068 21644
rect 4120 21632 4126 21684
rect 4154 21632 4160 21684
rect 4212 21672 4218 21684
rect 4890 21672 4896 21684
rect 4212 21644 4896 21672
rect 4212 21632 4218 21644
rect 4890 21632 4896 21644
rect 4948 21632 4954 21684
rect 5445 21675 5503 21681
rect 5445 21641 5457 21675
rect 5491 21672 5503 21675
rect 7374 21672 7380 21684
rect 5491 21644 7380 21672
rect 5491 21641 5503 21644
rect 5445 21635 5503 21641
rect 7374 21632 7380 21644
rect 7432 21632 7438 21684
rect 7650 21672 7656 21684
rect 7611 21644 7656 21672
rect 7650 21632 7656 21644
rect 7708 21632 7714 21684
rect 10410 21672 10416 21684
rect 8128 21644 10416 21672
rect 3896 21576 4660 21604
rect 3789 21567 3847 21573
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21536 1731 21539
rect 3053 21539 3111 21545
rect 1719 21508 2084 21536
rect 1719 21505 1731 21508
rect 1673 21499 1731 21505
rect 2056 21341 2084 21508
rect 3053 21505 3065 21539
rect 3099 21536 3111 21539
rect 3513 21539 3571 21545
rect 3099 21508 3133 21536
rect 3099 21505 3111 21508
rect 3053 21499 3111 21505
rect 3513 21505 3525 21539
rect 3559 21536 3571 21539
rect 3602 21536 3608 21548
rect 3559 21508 3608 21536
rect 3559 21505 3571 21508
rect 3513 21499 3571 21505
rect 2593 21471 2651 21477
rect 2593 21437 2605 21471
rect 2639 21468 2651 21471
rect 3068 21468 3096 21499
rect 3602 21496 3608 21508
rect 3660 21496 3666 21548
rect 3697 21539 3755 21545
rect 3697 21505 3709 21539
rect 3743 21505 3755 21539
rect 3697 21499 3755 21505
rect 3881 21539 3939 21545
rect 3881 21505 3893 21539
rect 3927 21536 3939 21539
rect 4246 21536 4252 21548
rect 3927 21508 4252 21536
rect 3927 21505 3939 21508
rect 3881 21499 3939 21505
rect 3712 21468 3740 21499
rect 4246 21496 4252 21508
rect 4304 21536 4310 21548
rect 4522 21536 4528 21548
rect 4304 21508 4528 21536
rect 4304 21496 4310 21508
rect 4522 21496 4528 21508
rect 4580 21496 4586 21548
rect 4154 21468 4160 21480
rect 2639 21440 3648 21468
rect 3712 21440 4160 21468
rect 2639 21437 2651 21440
rect 2593 21431 2651 21437
rect 2869 21403 2927 21409
rect 2869 21369 2881 21403
rect 2915 21400 2927 21403
rect 3234 21400 3240 21412
rect 2915 21372 3240 21400
rect 2915 21369 2927 21372
rect 2869 21363 2927 21369
rect 3234 21360 3240 21372
rect 3292 21360 3298 21412
rect 2041 21335 2099 21341
rect 2041 21301 2053 21335
rect 2087 21332 2099 21335
rect 2590 21332 2596 21344
rect 2087 21304 2596 21332
rect 2087 21301 2099 21304
rect 2041 21295 2099 21301
rect 2590 21292 2596 21304
rect 2648 21292 2654 21344
rect 3620 21332 3648 21440
rect 4154 21428 4160 21440
rect 4212 21428 4218 21480
rect 4632 21468 4660 21576
rect 4982 21564 4988 21616
rect 5040 21604 5046 21616
rect 5169 21607 5227 21613
rect 5169 21604 5181 21607
rect 5040 21576 5181 21604
rect 5040 21564 5046 21576
rect 5169 21573 5181 21576
rect 5215 21573 5227 21607
rect 5169 21567 5227 21573
rect 6638 21564 6644 21616
rect 6696 21604 6702 21616
rect 6696 21576 7144 21604
rect 6696 21564 6702 21576
rect 4798 21496 4804 21548
rect 4856 21536 4862 21548
rect 4893 21539 4951 21545
rect 4893 21536 4905 21539
rect 4856 21508 4905 21536
rect 4856 21496 4862 21508
rect 4893 21505 4905 21508
rect 4939 21505 4951 21539
rect 5074 21536 5080 21548
rect 5035 21508 5080 21536
rect 4893 21499 4951 21505
rect 5074 21496 5080 21508
rect 5132 21496 5138 21548
rect 5261 21539 5319 21545
rect 5261 21505 5273 21539
rect 5307 21536 5319 21539
rect 5534 21536 5540 21548
rect 5307 21508 5540 21536
rect 5307 21505 5319 21508
rect 5261 21499 5319 21505
rect 5534 21496 5540 21508
rect 5592 21496 5598 21548
rect 6733 21539 6791 21545
rect 6733 21505 6745 21539
rect 6779 21505 6791 21539
rect 6733 21499 6791 21505
rect 6638 21468 6644 21480
rect 4632 21440 6644 21468
rect 6638 21428 6644 21440
rect 6696 21428 6702 21480
rect 6748 21468 6776 21499
rect 6822 21496 6828 21548
rect 6880 21536 6886 21548
rect 7006 21536 7012 21548
rect 6880 21508 6925 21536
rect 6967 21508 7012 21536
rect 6880 21496 6886 21508
rect 7006 21496 7012 21508
rect 7064 21496 7070 21548
rect 7116 21545 7144 21576
rect 7466 21564 7472 21616
rect 7524 21604 7530 21616
rect 8128 21604 8156 21644
rect 10410 21632 10416 21644
rect 10468 21632 10474 21684
rect 10594 21632 10600 21684
rect 10652 21672 10658 21684
rect 10689 21675 10747 21681
rect 10689 21672 10701 21675
rect 10652 21644 10701 21672
rect 10652 21632 10658 21644
rect 10689 21641 10701 21644
rect 10735 21641 10747 21675
rect 10689 21635 10747 21641
rect 10781 21675 10839 21681
rect 10781 21641 10793 21675
rect 10827 21641 10839 21675
rect 10781 21635 10839 21641
rect 10965 21675 11023 21681
rect 10965 21641 10977 21675
rect 11011 21672 11023 21675
rect 11330 21672 11336 21684
rect 11011 21644 11336 21672
rect 11011 21641 11023 21644
rect 10965 21635 11023 21641
rect 8570 21604 8576 21616
rect 7524 21576 8156 21604
rect 8220 21576 8576 21604
rect 7524 21564 7530 21576
rect 7101 21539 7159 21545
rect 7101 21505 7113 21539
rect 7147 21505 7159 21539
rect 7101 21499 7159 21505
rect 7190 21496 7196 21548
rect 7248 21536 7254 21548
rect 7742 21536 7748 21548
rect 7248 21508 7748 21536
rect 7248 21496 7254 21508
rect 7742 21496 7748 21508
rect 7800 21496 7806 21548
rect 7834 21496 7840 21548
rect 7892 21536 7898 21548
rect 7929 21539 7987 21545
rect 7929 21536 7941 21539
rect 7892 21508 7941 21536
rect 7892 21496 7898 21508
rect 7929 21505 7941 21508
rect 7975 21505 7987 21539
rect 8110 21536 8116 21548
rect 8071 21508 8116 21536
rect 7929 21499 7987 21505
rect 8110 21496 8116 21508
rect 8168 21496 8174 21548
rect 8220 21545 8248 21576
rect 8570 21564 8576 21576
rect 8628 21564 8634 21616
rect 8938 21564 8944 21616
rect 8996 21604 9002 21616
rect 8996 21576 9536 21604
rect 8996 21564 9002 21576
rect 8205 21539 8263 21545
rect 8205 21505 8217 21539
rect 8251 21505 8263 21539
rect 8205 21499 8263 21505
rect 8389 21539 8447 21545
rect 8389 21505 8401 21539
rect 8435 21536 8447 21539
rect 8478 21536 8484 21548
rect 8435 21508 8484 21536
rect 8435 21505 8447 21508
rect 8389 21499 8447 21505
rect 6914 21468 6920 21480
rect 6748 21440 6920 21468
rect 6914 21428 6920 21440
rect 6972 21428 6978 21480
rect 7466 21428 7472 21480
rect 7524 21468 7530 21480
rect 8216 21468 8244 21499
rect 8478 21496 8484 21508
rect 8536 21496 8542 21548
rect 9398 21536 9404 21548
rect 9359 21508 9404 21536
rect 9398 21496 9404 21508
rect 9456 21496 9462 21548
rect 9508 21536 9536 21576
rect 9582 21564 9588 21616
rect 9640 21604 9646 21616
rect 10796 21604 10824 21635
rect 11330 21632 11336 21644
rect 11388 21632 11394 21684
rect 11517 21675 11575 21681
rect 11517 21641 11529 21675
rect 11563 21672 11575 21675
rect 12158 21672 12164 21684
rect 11563 21644 12164 21672
rect 11563 21641 11575 21644
rect 11517 21635 11575 21641
rect 12158 21632 12164 21644
rect 12216 21632 12222 21684
rect 13446 21632 13452 21684
rect 13504 21672 13510 21684
rect 18325 21675 18383 21681
rect 18325 21672 18337 21675
rect 13504 21644 15036 21672
rect 13504 21632 13510 21644
rect 9640 21576 10640 21604
rect 10796 21576 12020 21604
rect 9640 21564 9646 21576
rect 10612 21548 10640 21576
rect 9769 21539 9827 21545
rect 9769 21536 9781 21539
rect 9508 21508 9781 21536
rect 9769 21505 9781 21508
rect 9815 21505 9827 21539
rect 9769 21499 9827 21505
rect 9858 21496 9864 21548
rect 9916 21536 9922 21548
rect 9953 21539 10011 21545
rect 9953 21536 9965 21539
rect 9916 21508 9965 21536
rect 9916 21496 9922 21508
rect 9953 21505 9965 21508
rect 9999 21505 10011 21539
rect 10594 21536 10600 21548
rect 10555 21508 10600 21536
rect 9953 21499 10011 21505
rect 10594 21496 10600 21508
rect 10652 21536 10658 21548
rect 10652 21508 11652 21536
rect 10652 21496 10658 21508
rect 9582 21477 9588 21480
rect 7524 21440 8244 21468
rect 9559 21471 9588 21477
rect 7524 21428 7530 21440
rect 9559 21437 9571 21471
rect 9559 21431 9588 21437
rect 9582 21428 9588 21431
rect 9640 21428 9646 21480
rect 9674 21428 9680 21480
rect 9732 21468 9738 21480
rect 10965 21471 11023 21477
rect 10965 21468 10977 21471
rect 9732 21440 10977 21468
rect 9732 21428 9738 21440
rect 10965 21437 10977 21440
rect 11011 21468 11023 21471
rect 11514 21468 11520 21480
rect 11011 21440 11520 21468
rect 11011 21437 11023 21440
rect 10965 21431 11023 21437
rect 11514 21428 11520 21440
rect 11572 21428 11578 21480
rect 11624 21468 11652 21508
rect 11992 21477 12020 21576
rect 12342 21564 12348 21616
rect 12400 21604 12406 21616
rect 13326 21607 13384 21613
rect 13326 21604 13338 21607
rect 12400 21576 13338 21604
rect 12400 21564 12406 21576
rect 13326 21573 13338 21576
rect 13372 21573 13384 21607
rect 13326 21567 13384 21573
rect 13081 21539 13139 21545
rect 13081 21505 13093 21539
rect 13127 21536 13139 21539
rect 13814 21536 13820 21548
rect 13127 21508 13820 21536
rect 13127 21505 13139 21508
rect 13081 21499 13139 21505
rect 13814 21496 13820 21508
rect 13872 21496 13878 21548
rect 14826 21496 14832 21548
rect 14884 21536 14890 21548
rect 14921 21539 14979 21545
rect 14921 21536 14933 21539
rect 14884 21508 14933 21536
rect 14884 21496 14890 21508
rect 14921 21505 14933 21508
rect 14967 21505 14979 21539
rect 15008 21536 15036 21644
rect 15948 21644 18337 21672
rect 15948 21545 15976 21644
rect 18325 21641 18337 21644
rect 18371 21672 18383 21675
rect 18371 21644 19104 21672
rect 18371 21641 18383 21644
rect 18325 21635 18383 21641
rect 17129 21607 17187 21613
rect 17129 21573 17141 21607
rect 17175 21604 17187 21607
rect 18782 21604 18788 21616
rect 17175 21576 18788 21604
rect 17175 21573 17187 21576
rect 17129 21567 17187 21573
rect 18782 21564 18788 21576
rect 18840 21564 18846 21616
rect 15105 21539 15163 21545
rect 15105 21536 15117 21539
rect 15008 21508 15117 21536
rect 14921 21499 14979 21505
rect 15105 21505 15117 21508
rect 15151 21505 15163 21539
rect 15105 21499 15163 21505
rect 15933 21539 15991 21545
rect 15933 21505 15945 21539
rect 15979 21505 15991 21539
rect 16114 21536 16120 21548
rect 16075 21508 16120 21536
rect 15933 21499 15991 21505
rect 16114 21496 16120 21508
rect 16172 21496 16178 21548
rect 17954 21536 17960 21548
rect 17915 21508 17960 21536
rect 17954 21496 17960 21508
rect 18012 21496 18018 21548
rect 18046 21496 18052 21548
rect 18104 21536 18110 21548
rect 18877 21539 18935 21545
rect 18877 21536 18889 21539
rect 18104 21508 18889 21536
rect 18104 21496 18110 21508
rect 18877 21505 18889 21508
rect 18923 21505 18935 21539
rect 19076 21536 19104 21644
rect 19886 21632 19892 21684
rect 19944 21632 19950 21684
rect 19981 21675 20039 21681
rect 19981 21641 19993 21675
rect 20027 21672 20039 21675
rect 20622 21672 20628 21684
rect 20027 21644 20628 21672
rect 20027 21641 20039 21644
rect 19981 21635 20039 21641
rect 20622 21632 20628 21644
rect 20680 21632 20686 21684
rect 21269 21675 21327 21681
rect 21269 21641 21281 21675
rect 21315 21672 21327 21675
rect 23382 21672 23388 21684
rect 21315 21644 23388 21672
rect 21315 21641 21327 21644
rect 21269 21635 21327 21641
rect 23382 21632 23388 21644
rect 23440 21632 23446 21684
rect 23658 21632 23664 21684
rect 23716 21632 23722 21684
rect 24762 21632 24768 21684
rect 24820 21672 24826 21684
rect 25682 21672 25688 21684
rect 24820 21644 25360 21672
rect 25643 21644 25688 21672
rect 24820 21632 24826 21644
rect 19904 21604 19932 21632
rect 20806 21604 20812 21616
rect 19628 21576 19932 21604
rect 20767 21576 20812 21604
rect 19521 21539 19579 21545
rect 19521 21536 19533 21539
rect 19076 21508 19533 21536
rect 18877 21499 18935 21505
rect 19521 21505 19533 21508
rect 19567 21536 19579 21539
rect 19628 21536 19656 21576
rect 20806 21564 20812 21576
rect 20864 21604 20870 21616
rect 22002 21604 22008 21616
rect 20864 21576 22008 21604
rect 20864 21564 20870 21576
rect 22002 21564 22008 21576
rect 22060 21564 22066 21616
rect 22646 21604 22652 21616
rect 22204 21576 22652 21604
rect 19567 21508 19656 21536
rect 19790 21539 19848 21545
rect 19567 21505 19579 21508
rect 19521 21499 19579 21505
rect 19790 21505 19802 21539
rect 19836 21505 19848 21539
rect 19790 21499 19848 21505
rect 21085 21539 21143 21545
rect 21085 21505 21097 21539
rect 21131 21536 21143 21539
rect 21818 21536 21824 21548
rect 21131 21508 21824 21536
rect 21131 21505 21143 21508
rect 21085 21499 21143 21505
rect 11701 21471 11759 21477
rect 11701 21468 11713 21471
rect 11624 21440 11713 21468
rect 11701 21437 11713 21440
rect 11747 21437 11759 21471
rect 11701 21431 11759 21437
rect 11793 21471 11851 21477
rect 11793 21437 11805 21471
rect 11839 21437 11851 21471
rect 11793 21431 11851 21437
rect 11885 21471 11943 21477
rect 11885 21437 11897 21471
rect 11931 21437 11943 21471
rect 11885 21431 11943 21437
rect 11977 21471 12035 21477
rect 11977 21437 11989 21471
rect 12023 21468 12035 21471
rect 12250 21468 12256 21480
rect 12023 21440 12256 21468
rect 12023 21437 12035 21440
rect 11977 21431 12035 21437
rect 6549 21403 6607 21409
rect 6549 21369 6561 21403
rect 6595 21400 6607 21403
rect 8662 21400 8668 21412
rect 6595 21372 8668 21400
rect 6595 21369 6607 21372
rect 6549 21363 6607 21369
rect 8662 21360 8668 21372
rect 8720 21400 8726 21412
rect 8720 21372 9812 21400
rect 8720 21360 8726 21372
rect 4890 21332 4896 21344
rect 3620 21304 4896 21332
rect 4890 21292 4896 21304
rect 4948 21292 4954 21344
rect 4982 21292 4988 21344
rect 5040 21332 5046 21344
rect 7190 21332 7196 21344
rect 5040 21304 7196 21332
rect 5040 21292 5046 21304
rect 7190 21292 7196 21304
rect 7248 21292 7254 21344
rect 7374 21292 7380 21344
rect 7432 21332 7438 21344
rect 8021 21335 8079 21341
rect 8021 21332 8033 21335
rect 7432 21304 8033 21332
rect 7432 21292 7438 21304
rect 8021 21301 8033 21304
rect 8067 21332 8079 21335
rect 9674 21332 9680 21344
rect 8067 21304 9680 21332
rect 8067 21301 8079 21304
rect 8021 21295 8079 21301
rect 9674 21292 9680 21304
rect 9732 21292 9738 21344
rect 9784 21341 9812 21372
rect 10686 21360 10692 21412
rect 10744 21400 10750 21412
rect 11808 21400 11836 21431
rect 10744 21372 11836 21400
rect 10744 21360 10750 21372
rect 9769 21335 9827 21341
rect 9769 21301 9781 21335
rect 9815 21301 9827 21335
rect 9769 21295 9827 21301
rect 9858 21292 9864 21344
rect 9916 21332 9922 21344
rect 10870 21332 10876 21344
rect 9916 21304 10876 21332
rect 9916 21292 9922 21304
rect 10870 21292 10876 21304
rect 10928 21332 10934 21344
rect 11330 21332 11336 21344
rect 10928 21304 11336 21332
rect 10928 21292 10934 21304
rect 11330 21292 11336 21304
rect 11388 21292 11394 21344
rect 11514 21292 11520 21344
rect 11572 21332 11578 21344
rect 11900 21332 11928 21431
rect 12250 21428 12256 21440
rect 12308 21428 12314 21480
rect 15013 21471 15071 21477
rect 15013 21437 15025 21471
rect 15059 21468 15071 21471
rect 16132 21468 16160 21496
rect 17862 21468 17868 21480
rect 15059 21440 16160 21468
rect 17823 21440 17868 21468
rect 15059 21437 15071 21440
rect 15013 21431 15071 21437
rect 17862 21428 17868 21440
rect 17920 21428 17926 21480
rect 19610 21428 19616 21480
rect 19668 21468 19674 21480
rect 19812 21468 19840 21499
rect 21818 21496 21824 21508
rect 21876 21496 21882 21548
rect 22094 21496 22100 21548
rect 22152 21536 22158 21548
rect 22204 21545 22232 21576
rect 22646 21564 22652 21576
rect 22704 21564 22710 21616
rect 23106 21564 23112 21616
rect 23164 21604 23170 21616
rect 23477 21607 23535 21613
rect 23477 21604 23489 21607
rect 23164 21576 23489 21604
rect 23164 21564 23170 21576
rect 23477 21573 23489 21576
rect 23523 21573 23535 21607
rect 23477 21567 23535 21573
rect 23569 21607 23627 21613
rect 23569 21573 23581 21607
rect 23615 21604 23627 21607
rect 23676 21604 23704 21632
rect 23615 21576 24532 21604
rect 23615 21573 23627 21576
rect 23569 21567 23627 21573
rect 22189 21539 22247 21545
rect 22189 21536 22201 21539
rect 22152 21508 22201 21536
rect 22152 21496 22158 21508
rect 22189 21505 22201 21508
rect 22235 21505 22247 21539
rect 22189 21499 22247 21505
rect 22281 21539 22339 21545
rect 22281 21505 22293 21539
rect 22327 21536 22339 21539
rect 22554 21536 22560 21548
rect 22327 21508 22560 21536
rect 22327 21505 22339 21508
rect 22281 21499 22339 21505
rect 22554 21496 22560 21508
rect 22612 21496 22618 21548
rect 23293 21539 23351 21545
rect 23293 21505 23305 21539
rect 23339 21536 23351 21539
rect 23382 21536 23388 21548
rect 23339 21508 23388 21536
rect 23339 21505 23351 21508
rect 23293 21499 23351 21505
rect 23382 21496 23388 21508
rect 23440 21496 23446 21548
rect 23661 21539 23719 21545
rect 23661 21505 23673 21539
rect 23707 21536 23719 21539
rect 24397 21539 24455 21545
rect 24397 21536 24409 21539
rect 23707 21508 24409 21536
rect 23707 21505 23719 21508
rect 23661 21499 23719 21505
rect 24397 21505 24409 21508
rect 24443 21505 24455 21539
rect 24504 21536 24532 21576
rect 24578 21564 24584 21616
rect 24636 21604 24642 21616
rect 24854 21604 24860 21616
rect 24636 21576 24860 21604
rect 24636 21564 24642 21576
rect 24854 21564 24860 21576
rect 24912 21564 24918 21616
rect 25332 21613 25360 21644
rect 25682 21632 25688 21644
rect 25740 21632 25746 21684
rect 25958 21632 25964 21684
rect 26016 21672 26022 21684
rect 26329 21675 26387 21681
rect 26329 21672 26341 21675
rect 26016 21644 26341 21672
rect 26016 21632 26022 21644
rect 26329 21641 26341 21644
rect 26375 21641 26387 21675
rect 26329 21635 26387 21641
rect 25317 21607 25375 21613
rect 25317 21573 25329 21607
rect 25363 21573 25375 21607
rect 25317 21567 25375 21573
rect 25409 21607 25467 21613
rect 25409 21573 25421 21607
rect 25455 21604 25467 21607
rect 25590 21604 25596 21616
rect 25455 21576 25596 21604
rect 25455 21573 25467 21576
rect 25409 21567 25467 21573
rect 25590 21564 25596 21576
rect 25648 21604 25654 21616
rect 26142 21604 26148 21616
rect 25648 21576 26148 21604
rect 25648 21564 25654 21576
rect 26142 21564 26148 21576
rect 26200 21564 26206 21616
rect 24762 21536 24768 21548
rect 24504 21508 24768 21536
rect 24397 21499 24455 21505
rect 19886 21468 19892 21480
rect 19668 21440 19713 21468
rect 19812 21440 19892 21468
rect 19668 21428 19674 21440
rect 19886 21428 19892 21440
rect 19944 21428 19950 21480
rect 20530 21428 20536 21480
rect 20588 21468 20594 21480
rect 20901 21471 20959 21477
rect 20901 21468 20913 21471
rect 20588 21440 20913 21468
rect 20588 21428 20594 21440
rect 20901 21437 20913 21440
rect 20947 21437 20959 21471
rect 23566 21468 23572 21480
rect 20901 21431 20959 21437
rect 22480 21440 23572 21468
rect 22480 21409 22508 21440
rect 23566 21428 23572 21440
rect 23624 21428 23630 21480
rect 16025 21403 16083 21409
rect 16025 21369 16037 21403
rect 16071 21400 16083 21403
rect 22465 21403 22523 21409
rect 16071 21372 19334 21400
rect 16071 21369 16083 21372
rect 16025 21363 16083 21369
rect 11572 21304 11928 21332
rect 11572 21292 11578 21304
rect 14274 21292 14280 21344
rect 14332 21332 14338 21344
rect 14461 21335 14519 21341
rect 14461 21332 14473 21335
rect 14332 21304 14473 21332
rect 14332 21292 14338 21304
rect 14461 21301 14473 21304
rect 14507 21332 14519 21335
rect 15010 21332 15016 21344
rect 14507 21304 15016 21332
rect 14507 21301 14519 21304
rect 14461 21295 14519 21301
rect 15010 21292 15016 21304
rect 15068 21292 15074 21344
rect 17218 21332 17224 21344
rect 17179 21304 17224 21332
rect 17218 21292 17224 21304
rect 17276 21292 17282 21344
rect 18966 21332 18972 21344
rect 18927 21304 18972 21332
rect 18966 21292 18972 21304
rect 19024 21292 19030 21344
rect 19306 21332 19334 21372
rect 22465 21369 22477 21403
rect 22511 21369 22523 21403
rect 22465 21363 22523 21369
rect 23198 21360 23204 21412
rect 23256 21400 23262 21412
rect 23676 21400 23704 21499
rect 24762 21496 24768 21508
rect 24820 21496 24826 21548
rect 25038 21496 25044 21548
rect 25096 21536 25102 21548
rect 25133 21539 25191 21545
rect 25133 21536 25145 21539
rect 25096 21508 25145 21536
rect 25096 21496 25102 21508
rect 25133 21505 25145 21508
rect 25179 21505 25191 21539
rect 25133 21499 25191 21505
rect 25501 21539 25559 21545
rect 25501 21505 25513 21539
rect 25547 21536 25559 21539
rect 26050 21536 26056 21548
rect 25547 21508 26056 21536
rect 25547 21505 25559 21508
rect 25501 21499 25559 21505
rect 25516 21468 25544 21499
rect 26050 21496 26056 21508
rect 26108 21496 26114 21548
rect 26234 21536 26240 21548
rect 26195 21508 26240 21536
rect 26234 21496 26240 21508
rect 26292 21496 26298 21548
rect 26970 21536 26976 21548
rect 26931 21508 26976 21536
rect 26970 21496 26976 21508
rect 27028 21496 27034 21548
rect 27157 21539 27215 21545
rect 27157 21505 27169 21539
rect 27203 21505 27215 21539
rect 27157 21499 27215 21505
rect 24688 21440 25544 21468
rect 24688 21412 24716 21440
rect 26602 21428 26608 21480
rect 26660 21468 26666 21480
rect 27172 21468 27200 21499
rect 26660 21440 27200 21468
rect 26660 21428 26666 21440
rect 23256 21372 23704 21400
rect 24581 21403 24639 21409
rect 23256 21360 23262 21372
rect 24581 21369 24593 21403
rect 24627 21400 24639 21403
rect 24670 21400 24676 21412
rect 24627 21372 24676 21400
rect 24627 21369 24639 21372
rect 24581 21363 24639 21369
rect 24670 21360 24676 21372
rect 24728 21360 24734 21412
rect 19426 21332 19432 21344
rect 19306 21304 19432 21332
rect 19426 21292 19432 21304
rect 19484 21292 19490 21344
rect 19797 21335 19855 21341
rect 19797 21301 19809 21335
rect 19843 21332 19855 21335
rect 20622 21332 20628 21344
rect 19843 21304 20628 21332
rect 19843 21301 19855 21304
rect 19797 21295 19855 21301
rect 20622 21292 20628 21304
rect 20680 21292 20686 21344
rect 20898 21332 20904 21344
rect 20859 21304 20904 21332
rect 20898 21292 20904 21304
rect 20956 21292 20962 21344
rect 21634 21292 21640 21344
rect 21692 21332 21698 21344
rect 22005 21335 22063 21341
rect 22005 21332 22017 21335
rect 21692 21304 22017 21332
rect 21692 21292 21698 21304
rect 22005 21301 22017 21304
rect 22051 21301 22063 21335
rect 23842 21332 23848 21344
rect 23803 21304 23848 21332
rect 22005 21295 22063 21301
rect 23842 21292 23848 21304
rect 23900 21292 23906 21344
rect 25682 21292 25688 21344
rect 25740 21332 25746 21344
rect 26973 21335 27031 21341
rect 26973 21332 26985 21335
rect 25740 21304 26985 21332
rect 25740 21292 25746 21304
rect 26973 21301 26985 21304
rect 27019 21301 27031 21335
rect 26973 21295 27031 21301
rect 1104 21242 28060 21264
rect 1104 21190 5442 21242
rect 5494 21190 5506 21242
rect 5558 21190 5570 21242
rect 5622 21190 5634 21242
rect 5686 21190 5698 21242
rect 5750 21190 14428 21242
rect 14480 21190 14492 21242
rect 14544 21190 14556 21242
rect 14608 21190 14620 21242
rect 14672 21190 14684 21242
rect 14736 21190 23413 21242
rect 23465 21190 23477 21242
rect 23529 21190 23541 21242
rect 23593 21190 23605 21242
rect 23657 21190 23669 21242
rect 23721 21190 28060 21242
rect 1104 21168 28060 21190
rect 2409 21131 2467 21137
rect 2409 21097 2421 21131
rect 2455 21128 2467 21131
rect 4982 21128 4988 21140
rect 2455 21100 4988 21128
rect 2455 21097 2467 21100
rect 2409 21091 2467 21097
rect 4982 21088 4988 21100
rect 5040 21088 5046 21140
rect 5721 21131 5779 21137
rect 5721 21097 5733 21131
rect 5767 21128 5779 21131
rect 6638 21128 6644 21140
rect 5767 21100 6644 21128
rect 5767 21097 5779 21100
rect 5721 21091 5779 21097
rect 6638 21088 6644 21100
rect 6696 21088 6702 21140
rect 7650 21128 7656 21140
rect 7611 21100 7656 21128
rect 7650 21088 7656 21100
rect 7708 21088 7714 21140
rect 7837 21131 7895 21137
rect 7837 21097 7849 21131
rect 7883 21128 7895 21131
rect 8386 21128 8392 21140
rect 7883 21100 8392 21128
rect 7883 21097 7895 21100
rect 7837 21091 7895 21097
rect 8386 21088 8392 21100
rect 8444 21088 8450 21140
rect 9953 21131 10011 21137
rect 9953 21097 9965 21131
rect 9999 21128 10011 21131
rect 10686 21128 10692 21140
rect 9999 21100 10692 21128
rect 9999 21097 10011 21100
rect 9953 21091 10011 21097
rect 10686 21088 10692 21100
rect 10744 21088 10750 21140
rect 13998 21088 14004 21140
rect 14056 21128 14062 21140
rect 14277 21131 14335 21137
rect 14277 21128 14289 21131
rect 14056 21100 14289 21128
rect 14056 21088 14062 21100
rect 14277 21097 14289 21100
rect 14323 21097 14335 21131
rect 16850 21128 16856 21140
rect 14277 21091 14335 21097
rect 15028 21100 16712 21128
rect 16811 21100 16856 21128
rect 1210 21020 1216 21072
rect 1268 21060 1274 21072
rect 3421 21063 3479 21069
rect 1268 21032 2452 21060
rect 1268 21020 1274 21032
rect 1949 20927 2007 20933
rect 1949 20893 1961 20927
rect 1995 20924 2007 20927
rect 2222 20924 2228 20936
rect 1995 20896 2228 20924
rect 1995 20893 2007 20896
rect 1949 20887 2007 20893
rect 2222 20884 2228 20896
rect 2280 20884 2286 20936
rect 2424 20934 2452 21032
rect 3421 21029 3433 21063
rect 3467 21060 3479 21063
rect 3970 21060 3976 21072
rect 3467 21032 3976 21060
rect 3467 21029 3479 21032
rect 3421 21023 3479 21029
rect 3970 21020 3976 21032
rect 4028 21020 4034 21072
rect 6288 21032 6868 21060
rect 4154 20992 4160 21004
rect 3620 20964 4160 20992
rect 2332 20933 2452 20934
rect 2317 20927 2452 20933
rect 2317 20893 2329 20927
rect 2363 20906 2452 20927
rect 2593 20927 2651 20933
rect 2363 20893 2375 20906
rect 2317 20887 2375 20893
rect 2593 20893 2605 20927
rect 2639 20924 2651 20927
rect 2961 20927 3019 20933
rect 2961 20924 2973 20927
rect 2639 20896 2973 20924
rect 2639 20893 2651 20896
rect 2593 20887 2651 20893
rect 2961 20893 2973 20896
rect 3007 20924 3019 20927
rect 3142 20924 3148 20936
rect 3007 20896 3148 20924
rect 3007 20893 3019 20896
rect 2961 20887 3019 20893
rect 3142 20884 3148 20896
rect 3200 20884 3206 20936
rect 3620 20933 3648 20964
rect 4154 20952 4160 20964
rect 4212 20952 4218 21004
rect 6178 20992 6184 21004
rect 4540 20964 6184 20992
rect 3605 20927 3663 20933
rect 3605 20893 3617 20927
rect 3651 20893 3663 20927
rect 3605 20887 3663 20893
rect 3786 20884 3792 20936
rect 3844 20884 3850 20936
rect 3973 20927 4031 20933
rect 3973 20893 3985 20927
rect 4019 20924 4031 20927
rect 4540 20924 4568 20964
rect 6178 20952 6184 20964
rect 6236 20952 6242 21004
rect 4019 20896 4568 20924
rect 4617 20927 4675 20933
rect 4019 20893 4031 20896
rect 3973 20887 4031 20893
rect 4617 20893 4629 20927
rect 4663 20924 4675 20927
rect 4798 20924 4804 20936
rect 4663 20896 4804 20924
rect 4663 20893 4675 20896
rect 4617 20887 4675 20893
rect 4798 20884 4804 20896
rect 4856 20884 4862 20936
rect 5169 20927 5227 20933
rect 5169 20893 5181 20927
rect 5215 20893 5227 20927
rect 5169 20887 5227 20893
rect 5537 20927 5595 20933
rect 5537 20893 5549 20927
rect 5583 20924 5595 20927
rect 6288 20924 6316 21032
rect 6840 20992 6868 21032
rect 10134 21020 10140 21072
rect 10192 21060 10198 21072
rect 10192 21032 10237 21060
rect 10192 21020 10198 21032
rect 10318 21020 10324 21072
rect 10376 21060 10382 21072
rect 10965 21063 11023 21069
rect 10965 21060 10977 21063
rect 10376 21032 10977 21060
rect 10376 21020 10382 21032
rect 10965 21029 10977 21032
rect 11011 21029 11023 21063
rect 10965 21023 11023 21029
rect 7282 20992 7288 21004
rect 5583 20896 6316 20924
rect 6386 20964 6684 20992
rect 5583 20893 5595 20896
rect 5537 20887 5595 20893
rect 2866 20856 2872 20868
rect 1780 20828 2872 20856
rect 1780 20797 1808 20828
rect 2866 20816 2872 20828
rect 2924 20816 2930 20868
rect 3804 20856 3832 20884
rect 4706 20856 4712 20868
rect 3068 20828 3648 20856
rect 3804 20828 4712 20856
rect 1765 20791 1823 20797
rect 1765 20757 1777 20791
rect 1811 20757 1823 20791
rect 1765 20751 1823 20757
rect 2133 20791 2191 20797
rect 2133 20757 2145 20791
rect 2179 20788 2191 20791
rect 2314 20788 2320 20800
rect 2179 20760 2320 20788
rect 2179 20757 2191 20760
rect 2133 20751 2191 20757
rect 2314 20748 2320 20760
rect 2372 20748 2378 20800
rect 2406 20748 2412 20800
rect 2464 20788 2470 20800
rect 3068 20788 3096 20828
rect 3620 20800 3648 20828
rect 4706 20816 4712 20828
rect 4764 20816 4770 20868
rect 5184 20856 5212 20887
rect 5184 20828 5488 20856
rect 5460 20800 5488 20828
rect 3234 20788 3240 20800
rect 2464 20760 3096 20788
rect 3195 20760 3240 20788
rect 2464 20748 2470 20760
rect 3234 20748 3240 20760
rect 3292 20748 3298 20800
rect 3602 20748 3608 20800
rect 3660 20748 3666 20800
rect 3786 20788 3792 20800
rect 3747 20760 3792 20788
rect 3786 20748 3792 20760
rect 3844 20748 3850 20800
rect 5350 20788 5356 20800
rect 5311 20760 5356 20788
rect 5350 20748 5356 20760
rect 5408 20748 5414 20800
rect 5442 20748 5448 20800
rect 5500 20788 5506 20800
rect 6386 20788 6414 20964
rect 6656 20933 6684 20964
rect 6840 20964 7288 20992
rect 6840 20933 6868 20964
rect 7282 20952 7288 20964
rect 7340 20952 7346 21004
rect 7484 20964 11652 20992
rect 7484 20936 7512 20964
rect 6641 20927 6699 20933
rect 6641 20893 6653 20927
rect 6687 20893 6699 20927
rect 6641 20887 6699 20893
rect 6733 20927 6791 20933
rect 6733 20893 6745 20927
rect 6779 20893 6791 20927
rect 6733 20887 6791 20893
rect 6825 20927 6883 20933
rect 6825 20893 6837 20927
rect 6871 20893 6883 20927
rect 7466 20924 7472 20936
rect 7427 20896 7472 20924
rect 6825 20887 6883 20893
rect 6748 20856 6776 20887
rect 7466 20884 7472 20896
rect 7524 20884 7530 20936
rect 7653 20927 7711 20933
rect 7653 20893 7665 20927
rect 7699 20924 7711 20927
rect 7926 20924 7932 20936
rect 7699 20896 7932 20924
rect 7699 20893 7711 20896
rect 7653 20887 7711 20893
rect 7926 20884 7932 20896
rect 7984 20884 7990 20936
rect 8938 20924 8944 20936
rect 8899 20896 8944 20924
rect 8938 20884 8944 20896
rect 8996 20884 9002 20936
rect 9125 20927 9183 20933
rect 9125 20893 9137 20927
rect 9171 20893 9183 20927
rect 9582 20924 9588 20936
rect 9543 20896 9588 20924
rect 9125 20887 9183 20893
rect 8018 20856 8024 20868
rect 6748 20828 8024 20856
rect 8018 20816 8024 20828
rect 8076 20816 8082 20868
rect 9140 20856 9168 20887
rect 9582 20884 9588 20896
rect 9640 20884 9646 20936
rect 9674 20884 9680 20936
rect 9732 20924 9738 20936
rect 9950 20924 9956 20936
rect 9732 20896 9956 20924
rect 9732 20884 9738 20896
rect 9950 20884 9956 20896
rect 10008 20884 10014 20936
rect 10594 20924 10600 20936
rect 10555 20896 10600 20924
rect 10594 20884 10600 20896
rect 10652 20884 10658 20936
rect 10781 20927 10839 20933
rect 10781 20893 10793 20927
rect 10827 20924 10839 20927
rect 10870 20924 10876 20936
rect 10827 20896 10876 20924
rect 10827 20893 10839 20896
rect 10781 20887 10839 20893
rect 10870 20884 10876 20896
rect 10928 20884 10934 20936
rect 11330 20884 11336 20936
rect 11388 20924 11394 20936
rect 11624 20933 11652 20964
rect 11425 20927 11483 20933
rect 11425 20924 11437 20927
rect 11388 20896 11437 20924
rect 11388 20884 11394 20896
rect 11425 20893 11437 20896
rect 11471 20893 11483 20927
rect 11425 20887 11483 20893
rect 11609 20927 11667 20933
rect 11609 20893 11621 20927
rect 11655 20893 11667 20927
rect 11609 20887 11667 20893
rect 11790 20884 11796 20936
rect 11848 20924 11854 20936
rect 12069 20927 12127 20933
rect 12069 20924 12081 20927
rect 11848 20896 12081 20924
rect 11848 20884 11854 20896
rect 12069 20893 12081 20896
rect 12115 20924 12127 20927
rect 12115 20896 12434 20924
rect 12115 20893 12127 20896
rect 12069 20887 12127 20893
rect 9140 20828 10548 20856
rect 6730 20788 6736 20800
rect 5500 20760 6736 20788
rect 5500 20748 5506 20760
rect 6730 20748 6736 20760
rect 6788 20748 6794 20800
rect 7009 20791 7067 20797
rect 7009 20757 7021 20791
rect 7055 20788 7067 20791
rect 7190 20788 7196 20800
rect 7055 20760 7196 20788
rect 7055 20757 7067 20760
rect 7009 20751 7067 20757
rect 7190 20748 7196 20760
rect 7248 20748 7254 20800
rect 7558 20748 7564 20800
rect 7616 20788 7622 20800
rect 9030 20788 9036 20800
rect 7616 20760 9036 20788
rect 7616 20748 7622 20760
rect 9030 20748 9036 20760
rect 9088 20748 9094 20800
rect 9125 20791 9183 20797
rect 9125 20757 9137 20791
rect 9171 20788 9183 20791
rect 9674 20788 9680 20800
rect 9171 20760 9680 20788
rect 9171 20757 9183 20760
rect 9125 20751 9183 20757
rect 9674 20748 9680 20760
rect 9732 20748 9738 20800
rect 10520 20788 10548 20828
rect 10796 20828 11652 20856
rect 10796 20788 10824 20828
rect 11514 20788 11520 20800
rect 10520 20760 10824 20788
rect 11475 20760 11520 20788
rect 11514 20748 11520 20760
rect 11572 20748 11578 20800
rect 11624 20788 11652 20828
rect 11882 20816 11888 20868
rect 11940 20856 11946 20868
rect 12314 20859 12372 20865
rect 12314 20856 12326 20859
rect 11940 20828 12326 20856
rect 11940 20816 11946 20828
rect 12314 20825 12326 20828
rect 12360 20825 12372 20859
rect 12406 20856 12434 20896
rect 13078 20884 13084 20936
rect 13136 20924 13142 20936
rect 15028 20933 15056 21100
rect 16684 21060 16712 21100
rect 16850 21088 16856 21100
rect 16908 21088 16914 21140
rect 18966 21088 18972 21140
rect 19024 21128 19030 21140
rect 20806 21128 20812 21140
rect 19024 21100 20812 21128
rect 19024 21088 19030 21100
rect 20806 21088 20812 21100
rect 20864 21128 20870 21140
rect 21082 21128 21088 21140
rect 20864 21100 21088 21128
rect 20864 21088 20870 21100
rect 21082 21088 21088 21100
rect 21140 21088 21146 21140
rect 22370 21128 22376 21140
rect 22331 21100 22376 21128
rect 22370 21088 22376 21100
rect 22428 21088 22434 21140
rect 23750 21128 23756 21140
rect 23711 21100 23756 21128
rect 23750 21088 23756 21100
rect 23808 21088 23814 21140
rect 24394 21088 24400 21140
rect 24452 21088 24458 21140
rect 18322 21060 18328 21072
rect 16684 21032 18328 21060
rect 18322 21020 18328 21032
rect 18380 21020 18386 21072
rect 19886 21020 19892 21072
rect 19944 21060 19950 21072
rect 23106 21060 23112 21072
rect 19944 21032 23112 21060
rect 19944 21020 19950 21032
rect 23106 21020 23112 21032
rect 23164 21060 23170 21072
rect 24412 21060 24440 21088
rect 23164 21032 23428 21060
rect 23164 21020 23170 21032
rect 19904 20992 19932 21020
rect 21910 20992 21916 21004
rect 17788 20964 19932 20992
rect 20916 20964 21916 20992
rect 14093 20927 14151 20933
rect 14093 20924 14105 20927
rect 13136 20896 14105 20924
rect 13136 20884 13142 20896
rect 14093 20893 14105 20896
rect 14139 20893 14151 20927
rect 14093 20887 14151 20893
rect 15013 20927 15071 20933
rect 15013 20893 15025 20927
rect 15059 20893 15071 20927
rect 15013 20887 15071 20893
rect 15473 20927 15531 20933
rect 15473 20893 15485 20927
rect 15519 20924 15531 20927
rect 16298 20924 16304 20936
rect 15519 20896 16304 20924
rect 15519 20893 15531 20896
rect 15473 20887 15531 20893
rect 16298 20884 16304 20896
rect 16356 20924 16362 20936
rect 16758 20924 16764 20936
rect 16356 20896 16764 20924
rect 16356 20884 16362 20896
rect 16758 20884 16764 20896
rect 16816 20924 16822 20936
rect 17218 20924 17224 20936
rect 16816 20896 17224 20924
rect 16816 20884 16822 20896
rect 17218 20884 17224 20896
rect 17276 20884 17282 20936
rect 17788 20933 17816 20964
rect 17773 20927 17831 20933
rect 17773 20893 17785 20927
rect 17819 20893 17831 20927
rect 17773 20887 17831 20893
rect 18046 20884 18052 20936
rect 18104 20924 18110 20936
rect 18509 20927 18567 20933
rect 18509 20924 18521 20927
rect 18104 20896 18521 20924
rect 18104 20884 18110 20896
rect 18509 20893 18521 20896
rect 18555 20893 18567 20927
rect 19610 20924 19616 20936
rect 18509 20887 18567 20893
rect 19352 20896 19616 20924
rect 13814 20856 13820 20868
rect 12406 20828 13820 20856
rect 12314 20819 12372 20825
rect 13814 20816 13820 20828
rect 13872 20816 13878 20868
rect 15194 20816 15200 20868
rect 15252 20856 15258 20868
rect 15718 20859 15776 20865
rect 15718 20856 15730 20859
rect 15252 20828 15730 20856
rect 15252 20816 15258 20828
rect 15718 20825 15730 20828
rect 15764 20825 15776 20859
rect 15718 20819 15776 20825
rect 18693 20859 18751 20865
rect 18693 20825 18705 20859
rect 18739 20856 18751 20859
rect 19352 20856 19380 20896
rect 19610 20884 19616 20896
rect 19668 20924 19674 20936
rect 19797 20927 19855 20933
rect 19797 20924 19809 20927
rect 19668 20896 19809 20924
rect 19668 20884 19674 20896
rect 19797 20893 19809 20896
rect 19843 20893 19855 20927
rect 19797 20887 19855 20893
rect 19889 20927 19947 20933
rect 19889 20893 19901 20927
rect 19935 20893 19947 20927
rect 19889 20887 19947 20893
rect 20073 20927 20131 20933
rect 20073 20893 20085 20927
rect 20119 20893 20131 20927
rect 20073 20887 20131 20893
rect 20165 20927 20223 20933
rect 20165 20893 20177 20927
rect 20211 20924 20223 20927
rect 20346 20924 20352 20936
rect 20211 20896 20352 20924
rect 20211 20893 20223 20896
rect 20165 20887 20223 20893
rect 18739 20828 19380 20856
rect 18739 20825 18751 20828
rect 18693 20819 18751 20825
rect 19426 20816 19432 20868
rect 19484 20856 19490 20868
rect 19904 20856 19932 20887
rect 19484 20828 19932 20856
rect 20088 20856 20116 20887
rect 20346 20884 20352 20896
rect 20404 20884 20410 20936
rect 20530 20884 20536 20936
rect 20588 20924 20594 20936
rect 20916 20933 20944 20964
rect 21910 20952 21916 20964
rect 21968 20952 21974 21004
rect 22373 20995 22431 21001
rect 22373 20961 22385 20995
rect 22419 20992 22431 20995
rect 23290 20992 23296 21004
rect 22419 20964 23296 20992
rect 22419 20961 22431 20964
rect 22373 20955 22431 20961
rect 20809 20927 20867 20933
rect 20809 20924 20821 20927
rect 20588 20896 20821 20924
rect 20588 20884 20594 20896
rect 20809 20893 20821 20896
rect 20855 20893 20867 20927
rect 20809 20887 20867 20893
rect 20901 20927 20959 20933
rect 20901 20893 20913 20927
rect 20947 20893 20959 20927
rect 21082 20924 21088 20936
rect 21043 20896 21088 20924
rect 20901 20887 20959 20893
rect 21082 20884 21088 20896
rect 21140 20884 21146 20936
rect 21174 20884 21180 20936
rect 21232 20924 21238 20936
rect 21818 20924 21824 20936
rect 21232 20896 21277 20924
rect 21779 20896 21824 20924
rect 21232 20884 21238 20896
rect 21818 20884 21824 20896
rect 21876 20884 21882 20936
rect 22002 20884 22008 20936
rect 22060 20924 22066 20936
rect 22281 20927 22339 20933
rect 22281 20924 22293 20927
rect 22060 20896 22293 20924
rect 22060 20884 22066 20896
rect 22281 20893 22293 20896
rect 22327 20893 22339 20927
rect 22281 20887 22339 20893
rect 20990 20856 20996 20868
rect 20088 20828 20996 20856
rect 19484 20816 19490 20828
rect 20990 20816 20996 20828
rect 21048 20816 21054 20868
rect 22388 20856 22416 20955
rect 23290 20952 23296 20964
rect 23348 20952 23354 21004
rect 23400 21001 23428 21032
rect 23768 21032 24440 21060
rect 23768 21004 23796 21032
rect 23385 20995 23443 21001
rect 23385 20961 23397 20995
rect 23431 20961 23443 20995
rect 23385 20955 23443 20961
rect 23750 20952 23756 21004
rect 23808 20952 23814 21004
rect 24118 20952 24124 21004
rect 24176 20992 24182 21004
rect 24394 20992 24400 21004
rect 24176 20964 24400 20992
rect 24176 20952 24182 20964
rect 24394 20952 24400 20964
rect 24452 20952 24458 21004
rect 24946 20952 24952 21004
rect 25004 20992 25010 21004
rect 25317 20995 25375 21001
rect 25317 20992 25329 20995
rect 25004 20964 25329 20992
rect 25004 20952 25010 20964
rect 25317 20961 25329 20964
rect 25363 20961 25375 20995
rect 25958 20992 25964 21004
rect 25919 20964 25964 20992
rect 25317 20955 25375 20961
rect 25958 20952 25964 20964
rect 26016 20952 26022 21004
rect 22554 20924 22560 20936
rect 22515 20896 22560 20924
rect 22554 20884 22560 20896
rect 22612 20884 22618 20936
rect 23569 20927 23627 20933
rect 23569 20893 23581 20927
rect 23615 20924 23627 20927
rect 23842 20924 23848 20936
rect 23615 20896 23848 20924
rect 23615 20893 23627 20896
rect 23569 20887 23627 20893
rect 23842 20884 23848 20896
rect 23900 20884 23906 20936
rect 25774 20884 25780 20936
rect 25832 20924 25838 20936
rect 26217 20927 26275 20933
rect 26217 20924 26229 20927
rect 25832 20896 26229 20924
rect 25832 20884 25838 20896
rect 26217 20893 26229 20896
rect 26263 20893 26275 20927
rect 26217 20887 26275 20893
rect 22020 20828 22416 20856
rect 25225 20859 25283 20865
rect 22020 20800 22048 20828
rect 25225 20825 25237 20859
rect 25271 20856 25283 20859
rect 25314 20856 25320 20868
rect 25271 20828 25320 20856
rect 25271 20825 25283 20828
rect 25225 20819 25283 20825
rect 25314 20816 25320 20828
rect 25372 20816 25378 20868
rect 12158 20788 12164 20800
rect 11624 20760 12164 20788
rect 12158 20748 12164 20760
rect 12216 20748 12222 20800
rect 13449 20791 13507 20797
rect 13449 20757 13461 20791
rect 13495 20788 13507 20791
rect 13538 20788 13544 20800
rect 13495 20760 13544 20788
rect 13495 20757 13507 20760
rect 13449 20751 13507 20757
rect 13538 20748 13544 20760
rect 13596 20748 13602 20800
rect 14829 20791 14887 20797
rect 14829 20757 14841 20791
rect 14875 20788 14887 20791
rect 17586 20788 17592 20800
rect 14875 20760 17592 20788
rect 14875 20757 14887 20760
rect 14829 20751 14887 20757
rect 17586 20748 17592 20760
rect 17644 20748 17650 20800
rect 17862 20788 17868 20800
rect 17823 20760 17868 20788
rect 17862 20748 17868 20760
rect 17920 20748 17926 20800
rect 19613 20791 19671 20797
rect 19613 20757 19625 20791
rect 19659 20788 19671 20791
rect 20346 20788 20352 20800
rect 19659 20760 20352 20788
rect 19659 20757 19671 20760
rect 19613 20751 19671 20757
rect 20346 20748 20352 20760
rect 20404 20748 20410 20800
rect 20625 20791 20683 20797
rect 20625 20757 20637 20791
rect 20671 20788 20683 20791
rect 21358 20788 21364 20800
rect 20671 20760 21364 20788
rect 20671 20757 20683 20760
rect 20625 20751 20683 20757
rect 21358 20748 21364 20760
rect 21416 20748 21422 20800
rect 21634 20788 21640 20800
rect 21595 20760 21640 20788
rect 21634 20748 21640 20760
rect 21692 20748 21698 20800
rect 22002 20748 22008 20800
rect 22060 20748 22066 20800
rect 22741 20791 22799 20797
rect 22741 20757 22753 20791
rect 22787 20788 22799 20791
rect 24210 20788 24216 20800
rect 22787 20760 24216 20788
rect 22787 20757 22799 20760
rect 22741 20751 22799 20757
rect 24210 20748 24216 20760
rect 24268 20748 24274 20800
rect 24765 20791 24823 20797
rect 24765 20757 24777 20791
rect 24811 20788 24823 20791
rect 25038 20788 25044 20800
rect 24811 20760 25044 20788
rect 24811 20757 24823 20760
rect 24765 20751 24823 20757
rect 25038 20748 25044 20760
rect 25096 20748 25102 20800
rect 25133 20791 25191 20797
rect 25133 20757 25145 20791
rect 25179 20788 25191 20791
rect 25590 20788 25596 20800
rect 25179 20760 25596 20788
rect 25179 20757 25191 20760
rect 25133 20751 25191 20757
rect 25590 20748 25596 20760
rect 25648 20748 25654 20800
rect 26142 20748 26148 20800
rect 26200 20788 26206 20800
rect 27341 20791 27399 20797
rect 27341 20788 27353 20791
rect 26200 20760 27353 20788
rect 26200 20748 26206 20760
rect 27341 20757 27353 20760
rect 27387 20757 27399 20791
rect 27341 20751 27399 20757
rect 1104 20698 28060 20720
rect 1104 20646 9935 20698
rect 9987 20646 9999 20698
rect 10051 20646 10063 20698
rect 10115 20646 10127 20698
rect 10179 20646 10191 20698
rect 10243 20646 18920 20698
rect 18972 20646 18984 20698
rect 19036 20646 19048 20698
rect 19100 20646 19112 20698
rect 19164 20646 19176 20698
rect 19228 20646 28060 20698
rect 1104 20624 28060 20646
rect 6914 20584 6920 20596
rect 1780 20556 6500 20584
rect 6875 20556 6920 20584
rect 1780 20457 1808 20556
rect 5442 20516 5448 20528
rect 5092 20488 5448 20516
rect 1765 20451 1823 20457
rect 1765 20417 1777 20451
rect 1811 20417 1823 20451
rect 1765 20411 1823 20417
rect 2133 20451 2191 20457
rect 2133 20417 2145 20451
rect 2179 20448 2191 20451
rect 2593 20451 2651 20457
rect 2593 20448 2605 20451
rect 2179 20420 2605 20448
rect 2179 20417 2191 20420
rect 2133 20411 2191 20417
rect 2593 20417 2605 20420
rect 2639 20448 2651 20451
rect 2682 20448 2688 20460
rect 2639 20420 2688 20448
rect 2639 20417 2651 20420
rect 2593 20411 2651 20417
rect 2682 20408 2688 20420
rect 2740 20408 2746 20460
rect 3605 20451 3663 20457
rect 3605 20417 3617 20451
rect 3651 20417 3663 20451
rect 3605 20411 3663 20417
rect 4157 20451 4215 20457
rect 4157 20417 4169 20451
rect 4203 20417 4215 20451
rect 4890 20448 4896 20460
rect 4851 20420 4896 20448
rect 4157 20411 4215 20417
rect 1486 20340 1492 20392
rect 1544 20380 1550 20392
rect 1670 20380 1676 20392
rect 1544 20352 1676 20380
rect 1544 20340 1550 20352
rect 1670 20340 1676 20352
rect 1728 20340 1734 20392
rect 2222 20340 2228 20392
rect 2280 20380 2286 20392
rect 3620 20380 3648 20411
rect 2280 20352 3648 20380
rect 4172 20380 4200 20411
rect 4890 20408 4896 20420
rect 4948 20408 4954 20460
rect 5092 20457 5120 20488
rect 5442 20476 5448 20488
rect 5500 20476 5506 20528
rect 5077 20451 5135 20457
rect 5077 20417 5089 20451
rect 5123 20417 5135 20451
rect 5077 20411 5135 20417
rect 5353 20451 5411 20457
rect 5353 20417 5365 20451
rect 5399 20448 5411 20451
rect 6086 20448 6092 20460
rect 5399 20420 6092 20448
rect 5399 20417 5411 20420
rect 5353 20411 5411 20417
rect 6086 20408 6092 20420
rect 6144 20448 6150 20460
rect 6365 20451 6423 20457
rect 6365 20448 6377 20451
rect 6144 20420 6377 20448
rect 6144 20408 6150 20420
rect 6365 20417 6377 20420
rect 6411 20417 6423 20451
rect 6365 20411 6423 20417
rect 6178 20380 6184 20392
rect 4172 20352 6184 20380
rect 2280 20340 2286 20352
rect 6178 20340 6184 20352
rect 6236 20340 6242 20392
rect 6472 20380 6500 20556
rect 6914 20544 6920 20556
rect 6972 20544 6978 20596
rect 8846 20544 8852 20596
rect 8904 20584 8910 20596
rect 8904 20556 12664 20584
rect 8904 20544 8910 20556
rect 8018 20476 8024 20528
rect 8076 20516 8082 20528
rect 9030 20516 9036 20528
rect 8076 20488 9036 20516
rect 8076 20476 8082 20488
rect 9030 20476 9036 20488
rect 9088 20516 9094 20528
rect 9582 20516 9588 20528
rect 9088 20488 9588 20516
rect 9088 20476 9094 20488
rect 9582 20476 9588 20488
rect 9640 20516 9646 20528
rect 10594 20516 10600 20528
rect 9640 20488 10600 20516
rect 9640 20476 9646 20488
rect 10594 20476 10600 20488
rect 10652 20476 10658 20528
rect 11238 20476 11244 20528
rect 11296 20516 11302 20528
rect 11296 20488 12296 20516
rect 11296 20476 11302 20488
rect 6730 20448 6736 20460
rect 6643 20420 6736 20448
rect 6730 20408 6736 20420
rect 6788 20448 6794 20460
rect 7558 20448 7564 20460
rect 6788 20420 7564 20448
rect 6788 20408 6794 20420
rect 7558 20408 7564 20420
rect 7616 20408 7622 20460
rect 7650 20408 7656 20460
rect 7708 20448 7714 20460
rect 7708 20420 7753 20448
rect 7708 20408 7714 20420
rect 7834 20408 7840 20460
rect 7892 20448 7898 20460
rect 7929 20451 7987 20457
rect 7929 20448 7941 20451
rect 7892 20420 7941 20448
rect 7892 20408 7898 20420
rect 7929 20417 7941 20420
rect 7975 20417 7987 20451
rect 7929 20411 7987 20417
rect 9214 20408 9220 20460
rect 9272 20448 9278 20460
rect 9401 20451 9459 20457
rect 9401 20448 9413 20451
rect 9272 20420 9413 20448
rect 9272 20408 9278 20420
rect 9401 20417 9413 20420
rect 9447 20417 9459 20451
rect 9766 20448 9772 20460
rect 9727 20420 9772 20448
rect 9401 20411 9459 20417
rect 9766 20408 9772 20420
rect 9824 20408 9830 20460
rect 10781 20451 10839 20457
rect 10781 20417 10793 20451
rect 10827 20448 10839 20451
rect 11790 20448 11796 20460
rect 10827 20420 11796 20448
rect 10827 20417 10839 20420
rect 10781 20411 10839 20417
rect 10594 20380 10600 20392
rect 6472 20352 10600 20380
rect 10594 20340 10600 20352
rect 10652 20340 10658 20392
rect 4522 20272 4528 20324
rect 4580 20312 4586 20324
rect 4985 20315 5043 20321
rect 4985 20312 4997 20315
rect 4580 20284 4997 20312
rect 4580 20272 4586 20284
rect 4985 20281 4997 20284
rect 5031 20281 5043 20315
rect 7466 20312 7472 20324
rect 4985 20275 5043 20281
rect 6472 20284 7472 20312
rect 1486 20204 1492 20256
rect 1544 20244 1550 20256
rect 1581 20247 1639 20253
rect 1581 20244 1593 20247
rect 1544 20216 1593 20244
rect 1544 20204 1550 20216
rect 1581 20213 1593 20216
rect 1627 20213 1639 20247
rect 1581 20207 1639 20213
rect 2409 20247 2467 20253
rect 2409 20213 2421 20247
rect 2455 20244 2467 20247
rect 2866 20244 2872 20256
rect 2455 20216 2872 20244
rect 2455 20213 2467 20216
rect 2409 20207 2467 20213
rect 2866 20204 2872 20216
rect 2924 20204 2930 20256
rect 3421 20247 3479 20253
rect 3421 20213 3433 20247
rect 3467 20244 3479 20247
rect 4062 20244 4068 20256
rect 3467 20216 4068 20244
rect 3467 20213 3479 20216
rect 3421 20207 3479 20213
rect 4062 20204 4068 20216
rect 4120 20204 4126 20256
rect 4249 20247 4307 20253
rect 4249 20213 4261 20247
rect 4295 20244 4307 20247
rect 6472 20244 6500 20284
rect 7466 20272 7472 20284
rect 7524 20272 7530 20324
rect 8846 20312 8852 20324
rect 8266 20284 8852 20312
rect 6638 20244 6644 20256
rect 4295 20216 6500 20244
rect 6599 20216 6644 20244
rect 4295 20213 4307 20216
rect 4249 20207 4307 20213
rect 6638 20204 6644 20216
rect 6696 20204 6702 20256
rect 7006 20204 7012 20256
rect 7064 20244 7070 20256
rect 8266 20244 8294 20284
rect 8846 20272 8852 20284
rect 8904 20272 8910 20324
rect 9953 20315 10011 20321
rect 9953 20281 9965 20315
rect 9999 20312 10011 20315
rect 10796 20312 10824 20411
rect 11790 20408 11796 20420
rect 11848 20408 11854 20460
rect 12268 20457 12296 20488
rect 12161 20451 12219 20457
rect 12161 20417 12173 20451
rect 12207 20417 12219 20451
rect 12161 20411 12219 20417
rect 12253 20451 12311 20457
rect 12253 20417 12265 20451
rect 12299 20417 12311 20451
rect 12253 20411 12311 20417
rect 11882 20380 11888 20392
rect 11843 20352 11888 20380
rect 11882 20340 11888 20352
rect 11940 20340 11946 20392
rect 9999 20284 10824 20312
rect 10965 20315 11023 20321
rect 9999 20281 10011 20284
rect 9953 20275 10011 20281
rect 10965 20281 10977 20315
rect 11011 20312 11023 20315
rect 11146 20312 11152 20324
rect 11011 20284 11152 20312
rect 11011 20281 11023 20284
rect 10965 20275 11023 20281
rect 11146 20272 11152 20284
rect 11204 20272 11210 20324
rect 12176 20312 12204 20411
rect 12268 20380 12296 20411
rect 12342 20408 12348 20460
rect 12400 20457 12406 20460
rect 12400 20448 12408 20457
rect 12529 20451 12587 20457
rect 12400 20420 12445 20448
rect 12400 20411 12408 20420
rect 12529 20417 12541 20451
rect 12575 20448 12587 20451
rect 12636 20448 12664 20556
rect 12894 20544 12900 20596
rect 12952 20584 12958 20596
rect 13449 20587 13507 20593
rect 13449 20584 13461 20587
rect 12952 20556 13461 20584
rect 12952 20544 12958 20556
rect 13449 20553 13461 20556
rect 13495 20553 13507 20587
rect 13449 20547 13507 20553
rect 16942 20544 16948 20596
rect 17000 20584 17006 20596
rect 17402 20584 17408 20596
rect 17000 20556 17408 20584
rect 17000 20544 17006 20556
rect 17402 20544 17408 20556
rect 17460 20544 17466 20596
rect 19702 20544 19708 20596
rect 19760 20584 19766 20596
rect 19760 20556 20944 20584
rect 19760 20544 19766 20556
rect 13078 20476 13084 20528
rect 13136 20516 13142 20528
rect 13297 20519 13355 20525
rect 13136 20488 13181 20516
rect 13136 20476 13142 20488
rect 13297 20485 13309 20519
rect 13343 20516 13355 20519
rect 13998 20516 14004 20528
rect 13343 20488 14004 20516
rect 13343 20485 13355 20488
rect 13297 20479 13355 20485
rect 13998 20476 14004 20488
rect 14056 20476 14062 20528
rect 15654 20516 15660 20528
rect 14108 20488 15660 20516
rect 12575 20420 13768 20448
rect 12575 20417 12587 20420
rect 12529 20411 12587 20417
rect 12400 20408 12406 20411
rect 12802 20380 12808 20392
rect 12268 20352 12808 20380
rect 12802 20340 12808 20352
rect 12860 20340 12866 20392
rect 13740 20380 13768 20420
rect 13814 20408 13820 20460
rect 13872 20448 13878 20460
rect 13909 20451 13967 20457
rect 13909 20448 13921 20451
rect 13872 20420 13921 20448
rect 13872 20408 13878 20420
rect 13909 20417 13921 20420
rect 13955 20417 13967 20451
rect 14108 20448 14136 20488
rect 15654 20476 15660 20488
rect 15712 20516 15718 20528
rect 17862 20516 17868 20528
rect 15712 20488 17868 20516
rect 15712 20476 15718 20488
rect 14182 20457 14188 20460
rect 13909 20411 13967 20417
rect 14016 20420 14136 20448
rect 14016 20380 14044 20420
rect 14176 20411 14188 20457
rect 14240 20448 14246 20460
rect 14240 20420 14276 20448
rect 14182 20408 14188 20411
rect 14240 20408 14246 20420
rect 15286 20408 15292 20460
rect 15344 20448 15350 20460
rect 15933 20451 15991 20457
rect 15933 20448 15945 20451
rect 15344 20420 15945 20448
rect 15344 20408 15350 20420
rect 15933 20417 15945 20420
rect 15979 20417 15991 20451
rect 15933 20411 15991 20417
rect 16758 20408 16764 20460
rect 16816 20448 16822 20460
rect 16899 20451 16957 20457
rect 16899 20448 16911 20451
rect 16816 20420 16911 20448
rect 16816 20408 16822 20420
rect 16899 20417 16911 20420
rect 16945 20417 16957 20451
rect 17034 20448 17040 20460
rect 16995 20420 17040 20448
rect 16899 20411 16957 20417
rect 17034 20408 17040 20420
rect 17092 20408 17098 20460
rect 17328 20457 17356 20488
rect 17862 20476 17868 20488
rect 17920 20476 17926 20528
rect 17954 20476 17960 20528
rect 18012 20516 18018 20528
rect 18598 20516 18604 20528
rect 18012 20488 18604 20516
rect 18012 20476 18018 20488
rect 18598 20476 18604 20488
rect 18656 20476 18662 20528
rect 20916 20525 20944 20556
rect 20990 20544 20996 20596
rect 21048 20584 21054 20596
rect 21269 20587 21327 20593
rect 21269 20584 21281 20587
rect 21048 20556 21281 20584
rect 21048 20544 21054 20556
rect 21269 20553 21281 20556
rect 21315 20553 21327 20587
rect 21269 20547 21327 20553
rect 21358 20544 21364 20596
rect 21416 20584 21422 20596
rect 23033 20587 23091 20593
rect 23033 20584 23045 20587
rect 21416 20556 23045 20584
rect 21416 20544 21422 20556
rect 23033 20553 23045 20556
rect 23079 20553 23091 20587
rect 23033 20547 23091 20553
rect 23201 20587 23259 20593
rect 23201 20553 23213 20587
rect 23247 20553 23259 20587
rect 24026 20584 24032 20596
rect 23987 20556 24032 20584
rect 23201 20547 23259 20553
rect 20901 20519 20959 20525
rect 20901 20485 20913 20519
rect 20947 20485 20959 20519
rect 21117 20519 21175 20525
rect 21117 20516 21129 20519
rect 20901 20479 20959 20485
rect 21008 20488 21129 20516
rect 18046 20457 18052 20460
rect 17129 20451 17187 20457
rect 17129 20417 17141 20451
rect 17175 20417 17187 20451
rect 17129 20411 17187 20417
rect 17313 20451 17371 20457
rect 17313 20417 17325 20451
rect 17359 20417 17371 20451
rect 17313 20411 17371 20417
rect 18040 20411 18052 20457
rect 18104 20448 18110 20460
rect 18104 20420 18140 20448
rect 13740 20352 14044 20380
rect 15838 20340 15844 20392
rect 15896 20380 15902 20392
rect 15896 20352 16344 20380
rect 15896 20340 15902 20352
rect 12618 20312 12624 20324
rect 12176 20284 12624 20312
rect 12618 20272 12624 20284
rect 12676 20312 12682 20324
rect 13538 20312 13544 20324
rect 12676 20284 13544 20312
rect 12676 20272 12682 20284
rect 13538 20272 13544 20284
rect 13596 20272 13602 20324
rect 15289 20315 15347 20321
rect 15289 20281 15301 20315
rect 15335 20312 15347 20315
rect 16022 20312 16028 20324
rect 15335 20284 16028 20312
rect 15335 20281 15347 20284
rect 15289 20275 15347 20281
rect 7064 20216 8294 20244
rect 7064 20204 7070 20216
rect 9306 20204 9312 20256
rect 9364 20244 9370 20256
rect 9493 20247 9551 20253
rect 9493 20244 9505 20247
rect 9364 20216 9505 20244
rect 9364 20204 9370 20216
rect 9493 20213 9505 20216
rect 9539 20213 9551 20247
rect 11164 20244 11192 20272
rect 12066 20244 12072 20256
rect 11164 20216 12072 20244
rect 9493 20207 9551 20213
rect 12066 20204 12072 20216
rect 12124 20244 12130 20256
rect 13265 20247 13323 20253
rect 13265 20244 13277 20247
rect 12124 20216 13277 20244
rect 12124 20204 12130 20216
rect 13265 20213 13277 20216
rect 13311 20213 13323 20247
rect 13265 20207 13323 20213
rect 13814 20204 13820 20256
rect 13872 20244 13878 20256
rect 15102 20244 15108 20256
rect 13872 20216 15108 20244
rect 13872 20204 13878 20216
rect 15102 20204 15108 20216
rect 15160 20244 15166 20256
rect 15304 20244 15332 20275
rect 16022 20272 16028 20284
rect 16080 20272 16086 20324
rect 16316 20312 16344 20352
rect 16390 20340 16396 20392
rect 16448 20380 16454 20392
rect 17144 20380 17172 20411
rect 18046 20408 18052 20411
rect 18104 20408 18110 20420
rect 19518 20408 19524 20460
rect 19576 20448 19582 20460
rect 19613 20451 19671 20457
rect 19613 20448 19625 20451
rect 19576 20420 19625 20448
rect 19576 20408 19582 20420
rect 19613 20417 19625 20420
rect 19659 20417 19671 20451
rect 19886 20448 19892 20460
rect 19847 20420 19892 20448
rect 19613 20411 19671 20417
rect 19886 20408 19892 20420
rect 19944 20408 19950 20460
rect 20622 20408 20628 20460
rect 20680 20448 20686 20460
rect 21008 20448 21036 20488
rect 21117 20485 21129 20488
rect 21163 20485 21175 20519
rect 22833 20519 22891 20525
rect 21117 20479 21175 20485
rect 21836 20488 22140 20516
rect 21836 20460 21864 20488
rect 20680 20420 21036 20448
rect 20680 20408 20686 20420
rect 21818 20408 21824 20460
rect 21876 20408 21882 20460
rect 21910 20408 21916 20460
rect 21968 20448 21974 20460
rect 22112 20457 22140 20488
rect 22833 20485 22845 20519
rect 22879 20485 22891 20519
rect 23216 20516 23244 20547
rect 24026 20544 24032 20556
rect 24084 20544 24090 20596
rect 27338 20584 27344 20596
rect 27299 20556 27344 20584
rect 27338 20544 27344 20556
rect 27396 20544 27402 20596
rect 24854 20516 24860 20528
rect 23216 20488 24860 20516
rect 22833 20479 22891 20485
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 21968 20420 22017 20448
rect 21968 20408 21974 20420
rect 22005 20417 22017 20420
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 22097 20451 22155 20457
rect 22097 20417 22109 20451
rect 22143 20417 22155 20451
rect 22097 20411 22155 20417
rect 22186 20408 22192 20460
rect 22244 20448 22250 20460
rect 22281 20451 22339 20457
rect 22281 20448 22293 20451
rect 22244 20420 22293 20448
rect 22244 20408 22250 20420
rect 22281 20417 22293 20420
rect 22327 20417 22339 20451
rect 22281 20411 22339 20417
rect 22370 20408 22376 20460
rect 22428 20448 22434 20460
rect 22428 20420 22473 20448
rect 22428 20408 22434 20420
rect 16448 20352 17172 20380
rect 16448 20340 16454 20352
rect 17218 20340 17224 20392
rect 17276 20380 17282 20392
rect 17773 20383 17831 20389
rect 17773 20380 17785 20383
rect 17276 20352 17785 20380
rect 17276 20340 17282 20352
rect 17773 20349 17785 20352
rect 17819 20349 17831 20383
rect 22848 20380 22876 20479
rect 24854 20476 24860 20488
rect 24912 20476 24918 20528
rect 25038 20476 25044 20528
rect 25096 20516 25102 20528
rect 25501 20519 25559 20525
rect 25501 20516 25513 20519
rect 25096 20488 25513 20516
rect 25096 20476 25102 20488
rect 25501 20485 25513 20488
rect 25547 20485 25559 20519
rect 25501 20479 25559 20485
rect 23842 20408 23848 20460
rect 23900 20448 23906 20460
rect 24946 20448 24952 20460
rect 23900 20420 24952 20448
rect 23900 20408 23906 20420
rect 24946 20408 24952 20420
rect 25004 20448 25010 20460
rect 25317 20451 25375 20457
rect 25317 20448 25329 20451
rect 25004 20420 25329 20448
rect 25004 20408 25010 20420
rect 25317 20417 25329 20420
rect 25363 20417 25375 20451
rect 25590 20448 25596 20460
rect 25551 20420 25596 20448
rect 25317 20411 25375 20417
rect 25590 20408 25596 20420
rect 25648 20408 25654 20460
rect 25685 20451 25743 20457
rect 25685 20417 25697 20451
rect 25731 20448 25743 20451
rect 25774 20448 25780 20460
rect 25731 20420 25780 20448
rect 25731 20417 25743 20420
rect 25685 20411 25743 20417
rect 25774 20408 25780 20420
rect 25832 20408 25838 20460
rect 27157 20451 27215 20457
rect 27157 20448 27169 20451
rect 25884 20420 27169 20448
rect 17773 20343 17831 20349
rect 21376 20352 22876 20380
rect 24121 20383 24179 20389
rect 16316 20284 17816 20312
rect 15160 20216 15332 20244
rect 15160 20204 15166 20216
rect 15470 20204 15476 20256
rect 15528 20244 15534 20256
rect 15749 20247 15807 20253
rect 15749 20244 15761 20247
rect 15528 20216 15761 20244
rect 15528 20204 15534 20216
rect 15749 20213 15761 20216
rect 15795 20213 15807 20247
rect 15749 20207 15807 20213
rect 16574 20204 16580 20256
rect 16632 20244 16638 20256
rect 16669 20247 16727 20253
rect 16669 20244 16681 20247
rect 16632 20216 16681 20244
rect 16632 20204 16638 20216
rect 16669 20213 16681 20216
rect 16715 20213 16727 20247
rect 17788 20244 17816 20284
rect 18892 20284 21128 20312
rect 18892 20244 18920 20284
rect 19150 20244 19156 20256
rect 17788 20216 18920 20244
rect 19063 20216 19156 20244
rect 16669 20207 16727 20213
rect 19150 20204 19156 20216
rect 19208 20244 19214 20256
rect 19426 20244 19432 20256
rect 19208 20216 19432 20244
rect 19208 20204 19214 20216
rect 19426 20204 19432 20216
rect 19484 20204 19490 20256
rect 21100 20253 21128 20284
rect 21376 20256 21404 20352
rect 24121 20349 24133 20383
rect 24167 20349 24179 20383
rect 24121 20343 24179 20349
rect 24136 20312 24164 20343
rect 24210 20340 24216 20392
rect 24268 20380 24274 20392
rect 24268 20352 24313 20380
rect 24268 20340 24274 20352
rect 24946 20312 24952 20324
rect 24136 20284 24952 20312
rect 24946 20272 24952 20284
rect 25004 20272 25010 20324
rect 25884 20321 25912 20420
rect 27157 20417 27169 20420
rect 27203 20417 27215 20451
rect 27157 20411 27215 20417
rect 26326 20340 26332 20392
rect 26384 20380 26390 20392
rect 26973 20383 27031 20389
rect 26973 20380 26985 20383
rect 26384 20352 26985 20380
rect 26384 20340 26390 20352
rect 26973 20349 26985 20352
rect 27019 20349 27031 20383
rect 26973 20343 27031 20349
rect 25869 20315 25927 20321
rect 25869 20281 25881 20315
rect 25915 20281 25927 20315
rect 25869 20275 25927 20281
rect 21085 20247 21143 20253
rect 21085 20213 21097 20247
rect 21131 20244 21143 20247
rect 21358 20244 21364 20256
rect 21131 20216 21364 20244
rect 21131 20213 21143 20216
rect 21085 20207 21143 20213
rect 21358 20204 21364 20216
rect 21416 20204 21422 20256
rect 21821 20247 21879 20253
rect 21821 20213 21833 20247
rect 21867 20244 21879 20247
rect 23017 20247 23075 20253
rect 23017 20244 23029 20247
rect 21867 20216 23029 20244
rect 21867 20213 21879 20216
rect 21821 20207 21879 20213
rect 23017 20213 23029 20216
rect 23063 20213 23075 20247
rect 23017 20207 23075 20213
rect 23661 20247 23719 20253
rect 23661 20213 23673 20247
rect 23707 20244 23719 20247
rect 24118 20244 24124 20256
rect 23707 20216 24124 20244
rect 23707 20213 23719 20216
rect 23661 20207 23719 20213
rect 24118 20204 24124 20216
rect 24176 20204 24182 20256
rect 1104 20154 28060 20176
rect 1104 20102 5442 20154
rect 5494 20102 5506 20154
rect 5558 20102 5570 20154
rect 5622 20102 5634 20154
rect 5686 20102 5698 20154
rect 5750 20102 14428 20154
rect 14480 20102 14492 20154
rect 14544 20102 14556 20154
rect 14608 20102 14620 20154
rect 14672 20102 14684 20154
rect 14736 20102 23413 20154
rect 23465 20102 23477 20154
rect 23529 20102 23541 20154
rect 23593 20102 23605 20154
rect 23657 20102 23669 20154
rect 23721 20102 28060 20154
rect 1104 20080 28060 20102
rect 1854 20000 1860 20052
rect 1912 20040 1918 20052
rect 3602 20040 3608 20052
rect 1912 20012 3608 20040
rect 1912 20000 1918 20012
rect 3602 20000 3608 20012
rect 3660 20000 3666 20052
rect 4062 20000 4068 20052
rect 4120 20040 4126 20052
rect 5258 20040 5264 20052
rect 4120 20012 5120 20040
rect 5219 20012 5264 20040
rect 4120 20000 4126 20012
rect 1673 19975 1731 19981
rect 1673 19941 1685 19975
rect 1719 19972 1731 19975
rect 2406 19972 2412 19984
rect 1719 19944 2412 19972
rect 1719 19941 1731 19944
rect 1673 19935 1731 19941
rect 2406 19932 2412 19944
rect 2464 19932 2470 19984
rect 4430 19972 4436 19984
rect 4391 19944 4436 19972
rect 4430 19932 4436 19944
rect 4488 19932 4494 19984
rect 5092 19972 5120 20012
rect 5258 20000 5264 20012
rect 5316 20000 5322 20052
rect 6181 20043 6239 20049
rect 6181 20009 6193 20043
rect 6227 20040 6239 20043
rect 7650 20040 7656 20052
rect 6227 20012 7656 20040
rect 6227 20009 6239 20012
rect 6181 20003 6239 20009
rect 7650 20000 7656 20012
rect 7708 20000 7714 20052
rect 8110 20000 8116 20052
rect 8168 20040 8174 20052
rect 11514 20040 11520 20052
rect 8168 20012 11520 20040
rect 8168 20000 8174 20012
rect 11514 20000 11520 20012
rect 11572 20000 11578 20052
rect 13446 20040 13452 20052
rect 12452 20012 13452 20040
rect 5092 19944 7696 19972
rect 7668 19916 7696 19944
rect 8478 19932 8484 19984
rect 8536 19972 8542 19984
rect 8536 19944 9628 19972
rect 8536 19932 8542 19944
rect 2225 19907 2283 19913
rect 2225 19904 2237 19907
rect 1872 19876 2237 19904
rect 1872 19845 1900 19876
rect 2225 19873 2237 19876
rect 2271 19904 2283 19907
rect 4062 19904 4068 19916
rect 2271 19876 4068 19904
rect 2271 19873 2283 19876
rect 2225 19867 2283 19873
rect 4062 19864 4068 19876
rect 4120 19864 4126 19916
rect 5000 19876 6132 19904
rect 5000 19845 5028 19876
rect 6104 19848 6132 19876
rect 6178 19864 6184 19916
rect 6236 19904 6242 19916
rect 6733 19907 6791 19913
rect 6733 19904 6745 19907
rect 6236 19876 6745 19904
rect 6236 19864 6242 19876
rect 6733 19873 6745 19876
rect 6779 19904 6791 19907
rect 6822 19904 6828 19916
rect 6779 19876 6828 19904
rect 6779 19873 6791 19876
rect 6733 19867 6791 19873
rect 6822 19864 6828 19876
rect 6880 19864 6886 19916
rect 7650 19864 7656 19916
rect 7708 19864 7714 19916
rect 8570 19864 8576 19916
rect 8628 19904 8634 19916
rect 8938 19904 8944 19916
rect 8628 19876 8944 19904
rect 8628 19864 8634 19876
rect 8938 19864 8944 19876
rect 8996 19904 9002 19916
rect 8996 19876 9352 19904
rect 8996 19864 9002 19876
rect 1857 19839 1915 19845
rect 1857 19805 1869 19839
rect 1903 19805 1915 19839
rect 1857 19799 1915 19805
rect 2501 19839 2559 19845
rect 2501 19805 2513 19839
rect 2547 19805 2559 19839
rect 2501 19799 2559 19805
rect 3237 19839 3295 19845
rect 3237 19805 3249 19839
rect 3283 19836 3295 19839
rect 4985 19839 5043 19845
rect 3283 19808 4844 19836
rect 3283 19805 3295 19808
rect 3237 19799 3295 19805
rect 2516 19768 2544 19799
rect 4246 19768 4252 19780
rect 2516 19740 3648 19768
rect 4207 19740 4252 19768
rect 3620 19712 3648 19740
rect 4246 19728 4252 19740
rect 4304 19728 4310 19780
rect 1118 19660 1124 19712
rect 1176 19700 1182 19712
rect 2317 19703 2375 19709
rect 2317 19700 2329 19703
rect 1176 19672 2329 19700
rect 1176 19660 1182 19672
rect 2317 19669 2329 19672
rect 2363 19669 2375 19703
rect 3050 19700 3056 19712
rect 3011 19672 3056 19700
rect 2317 19663 2375 19669
rect 3050 19660 3056 19672
rect 3108 19660 3114 19712
rect 3602 19660 3608 19712
rect 3660 19660 3666 19712
rect 4816 19700 4844 19808
rect 4985 19805 4997 19839
rect 5031 19805 5043 19839
rect 4985 19799 5043 19805
rect 5169 19839 5227 19845
rect 5169 19805 5181 19839
rect 5215 19836 5227 19839
rect 5258 19836 5264 19848
rect 5215 19808 5264 19836
rect 5215 19805 5227 19808
rect 5169 19799 5227 19805
rect 5258 19796 5264 19808
rect 5316 19796 5322 19848
rect 5353 19839 5411 19845
rect 5353 19805 5365 19839
rect 5399 19805 5411 19839
rect 6086 19836 6092 19848
rect 6047 19808 6092 19836
rect 5353 19799 5411 19805
rect 4890 19728 4896 19780
rect 4948 19768 4954 19780
rect 5368 19768 5396 19799
rect 6086 19796 6092 19808
rect 6144 19796 6150 19848
rect 6638 19796 6644 19848
rect 6696 19836 6702 19848
rect 9324 19845 9352 19876
rect 9600 19848 9628 19944
rect 12452 19913 12480 20012
rect 13446 20000 13452 20012
rect 13504 20000 13510 20052
rect 13998 20000 14004 20052
rect 14056 20040 14062 20052
rect 14093 20043 14151 20049
rect 14093 20040 14105 20043
rect 14056 20012 14105 20040
rect 14056 20000 14062 20012
rect 14093 20009 14105 20012
rect 14139 20009 14151 20043
rect 15194 20040 15200 20052
rect 15155 20012 15200 20040
rect 14093 20003 14151 20009
rect 15194 20000 15200 20012
rect 15252 20000 15258 20052
rect 17034 20040 17040 20052
rect 15580 20012 17040 20040
rect 14274 19972 14280 19984
rect 12535 19944 14280 19972
rect 12437 19907 12495 19913
rect 12437 19873 12449 19907
rect 12483 19873 12495 19907
rect 12437 19867 12495 19873
rect 7009 19839 7067 19845
rect 7009 19836 7021 19839
rect 6696 19808 7021 19836
rect 6696 19796 6702 19808
rect 7009 19805 7021 19808
rect 7055 19836 7067 19839
rect 8113 19839 8171 19845
rect 8113 19836 8125 19839
rect 7055 19808 8125 19836
rect 7055 19805 7067 19808
rect 7009 19799 7067 19805
rect 8113 19805 8125 19808
rect 8159 19805 8171 19839
rect 8113 19799 8171 19805
rect 9217 19839 9275 19845
rect 9217 19805 9229 19839
rect 9263 19805 9275 19839
rect 9217 19799 9275 19805
rect 9309 19839 9367 19845
rect 9309 19805 9321 19839
rect 9355 19805 9367 19839
rect 9309 19799 9367 19805
rect 9401 19839 9459 19845
rect 9401 19805 9413 19839
rect 9447 19836 9459 19839
rect 9490 19836 9496 19848
rect 9447 19808 9496 19836
rect 9447 19805 9459 19808
rect 9401 19799 9459 19805
rect 6656 19768 6684 19796
rect 4948 19740 6684 19768
rect 4948 19728 4954 19740
rect 6914 19728 6920 19780
rect 6972 19768 6978 19780
rect 7374 19768 7380 19780
rect 6972 19740 7380 19768
rect 6972 19728 6978 19740
rect 7374 19728 7380 19740
rect 7432 19728 7438 19780
rect 8297 19771 8355 19777
rect 8297 19737 8309 19771
rect 8343 19768 8355 19771
rect 9030 19768 9036 19780
rect 8343 19740 9036 19768
rect 8343 19737 8355 19740
rect 8297 19731 8355 19737
rect 9030 19728 9036 19740
rect 9088 19728 9094 19780
rect 7466 19700 7472 19712
rect 4816 19672 7472 19700
rect 7466 19660 7472 19672
rect 7524 19660 7530 19712
rect 8386 19660 8392 19712
rect 8444 19700 8450 19712
rect 8941 19703 8999 19709
rect 8941 19700 8953 19703
rect 8444 19672 8953 19700
rect 8444 19660 8450 19672
rect 8941 19669 8953 19672
rect 8987 19669 8999 19703
rect 9232 19700 9260 19799
rect 9490 19796 9496 19808
rect 9548 19796 9554 19848
rect 9582 19796 9588 19848
rect 9640 19836 9646 19848
rect 10318 19836 10324 19848
rect 9640 19808 9733 19836
rect 10279 19808 10324 19836
rect 9640 19796 9646 19808
rect 10318 19796 10324 19808
rect 10376 19796 10382 19848
rect 12066 19836 12072 19848
rect 10520 19808 12072 19836
rect 9858 19728 9864 19780
rect 9916 19768 9922 19780
rect 10520 19768 10548 19808
rect 12066 19796 12072 19808
rect 12124 19836 12130 19848
rect 12253 19839 12311 19845
rect 12253 19836 12265 19839
rect 12124 19808 12265 19836
rect 12124 19796 12130 19808
rect 12253 19805 12265 19808
rect 12299 19805 12311 19839
rect 12253 19799 12311 19805
rect 12345 19839 12403 19845
rect 12345 19805 12357 19839
rect 12391 19836 12403 19839
rect 12535 19836 12563 19944
rect 14274 19932 14280 19944
rect 14332 19932 14338 19984
rect 12802 19864 12808 19916
rect 12860 19904 12866 19916
rect 14366 19904 14372 19916
rect 12860 19876 13400 19904
rect 14327 19876 14372 19904
rect 12860 19864 12866 19876
rect 12391 19808 12563 19836
rect 12621 19839 12679 19845
rect 12391 19805 12403 19808
rect 12345 19799 12403 19805
rect 12621 19805 12633 19839
rect 12667 19836 12679 19839
rect 13262 19836 13268 19848
rect 12667 19808 13268 19836
rect 12667 19805 12679 19808
rect 12621 19799 12679 19805
rect 13262 19796 13268 19808
rect 13320 19796 13326 19848
rect 13372 19845 13400 19876
rect 14366 19864 14372 19876
rect 14424 19864 14430 19916
rect 15580 19904 15608 20012
rect 17034 20000 17040 20012
rect 17092 20000 17098 20052
rect 18046 20000 18052 20052
rect 18104 20040 18110 20052
rect 18141 20043 18199 20049
rect 18141 20040 18153 20043
rect 18104 20012 18153 20040
rect 18104 20000 18110 20012
rect 18141 20009 18153 20012
rect 18187 20009 18199 20043
rect 18141 20003 18199 20009
rect 18690 20000 18696 20052
rect 18748 20040 18754 20052
rect 19334 20040 19340 20052
rect 18748 20012 19340 20040
rect 18748 20000 18754 20012
rect 19334 20000 19340 20012
rect 19392 20000 19398 20052
rect 19889 20043 19947 20049
rect 19889 20009 19901 20043
rect 19935 20040 19947 20043
rect 21082 20040 21088 20052
rect 19935 20012 21088 20040
rect 19935 20009 19947 20012
rect 19889 20003 19947 20009
rect 21082 20000 21088 20012
rect 21140 20000 21146 20052
rect 21358 20040 21364 20052
rect 21319 20012 21364 20040
rect 21358 20000 21364 20012
rect 21416 20000 21422 20052
rect 22189 20043 22247 20049
rect 22189 20009 22201 20043
rect 22235 20040 22247 20043
rect 22370 20040 22376 20052
rect 22235 20012 22376 20040
rect 22235 20009 22247 20012
rect 22189 20003 22247 20009
rect 22370 20000 22376 20012
rect 22428 20000 22434 20052
rect 23845 20043 23903 20049
rect 23845 20009 23857 20043
rect 23891 20040 23903 20043
rect 24302 20040 24308 20052
rect 23891 20012 24308 20040
rect 23891 20009 23903 20012
rect 23845 20003 23903 20009
rect 24302 20000 24308 20012
rect 24360 20000 24366 20052
rect 26326 20040 26332 20052
rect 25976 20012 26332 20040
rect 15654 19932 15660 19984
rect 15712 19932 15718 19984
rect 18064 19944 20300 19972
rect 15120 19876 15608 19904
rect 15672 19904 15700 19932
rect 18064 19916 18092 19944
rect 15672 19876 15884 19904
rect 13357 19839 13415 19845
rect 13357 19805 13369 19839
rect 13403 19836 13415 19839
rect 14274 19836 14280 19848
rect 13403 19808 13860 19836
rect 14235 19808 14280 19836
rect 13403 19805 13415 19808
rect 13357 19799 13415 19805
rect 9916 19740 10548 19768
rect 10588 19771 10646 19777
rect 9916 19728 9922 19740
rect 10588 19737 10600 19771
rect 10634 19768 10646 19771
rect 10870 19768 10876 19780
rect 10634 19740 10876 19768
rect 10634 19737 10646 19740
rect 10588 19731 10646 19737
rect 10870 19728 10876 19740
rect 10928 19728 10934 19780
rect 13173 19771 13231 19777
rect 11624 19740 13032 19768
rect 11624 19700 11652 19740
rect 9232 19672 11652 19700
rect 11701 19703 11759 19709
rect 8941 19663 8999 19669
rect 11701 19669 11713 19703
rect 11747 19700 11759 19703
rect 12250 19700 12256 19712
rect 11747 19672 12256 19700
rect 11747 19669 11759 19672
rect 11701 19663 11759 19669
rect 12250 19660 12256 19672
rect 12308 19660 12314 19712
rect 12529 19703 12587 19709
rect 12529 19669 12541 19703
rect 12575 19700 12587 19703
rect 12894 19700 12900 19712
rect 12575 19672 12900 19700
rect 12575 19669 12587 19672
rect 12529 19663 12587 19669
rect 12894 19660 12900 19672
rect 12952 19660 12958 19712
rect 13004 19700 13032 19740
rect 13173 19737 13185 19771
rect 13219 19768 13231 19771
rect 13722 19768 13728 19780
rect 13219 19740 13728 19768
rect 13219 19737 13231 19740
rect 13173 19731 13231 19737
rect 13722 19728 13728 19740
rect 13780 19728 13786 19780
rect 13832 19768 13860 19808
rect 14274 19796 14280 19808
rect 14332 19796 14338 19848
rect 14458 19836 14464 19848
rect 14419 19808 14464 19836
rect 14458 19796 14464 19808
rect 14516 19796 14522 19848
rect 14553 19839 14611 19845
rect 14553 19805 14565 19839
rect 14599 19836 14611 19839
rect 15010 19836 15016 19848
rect 14599 19808 15016 19836
rect 14599 19805 14611 19808
rect 14553 19799 14611 19805
rect 15010 19796 15016 19808
rect 15068 19796 15074 19848
rect 15120 19768 15148 19876
rect 15580 19845 15608 19876
rect 15473 19839 15531 19845
rect 15473 19805 15485 19839
rect 15519 19805 15531 19839
rect 15473 19799 15531 19805
rect 15565 19839 15623 19845
rect 15565 19805 15577 19839
rect 15611 19805 15623 19839
rect 15565 19799 15623 19805
rect 13832 19740 15148 19768
rect 15488 19768 15516 19799
rect 15654 19796 15660 19848
rect 15712 19836 15718 19848
rect 15856 19845 15884 19876
rect 18046 19864 18052 19916
rect 18104 19864 18110 19916
rect 18509 19907 18567 19913
rect 18509 19873 18521 19907
rect 18555 19904 18567 19907
rect 19702 19904 19708 19916
rect 18555 19876 19708 19904
rect 18555 19873 18567 19876
rect 18509 19867 18567 19873
rect 19702 19864 19708 19876
rect 19760 19864 19766 19916
rect 15841 19839 15899 19845
rect 15712 19808 15757 19836
rect 15712 19796 15718 19808
rect 15841 19805 15853 19839
rect 15887 19805 15899 19839
rect 16298 19836 16304 19848
rect 16259 19808 16304 19836
rect 15841 19799 15899 19805
rect 16298 19796 16304 19808
rect 16356 19796 16362 19848
rect 16574 19845 16580 19848
rect 16568 19836 16580 19845
rect 16535 19808 16580 19836
rect 16568 19799 16580 19808
rect 16574 19796 16580 19799
rect 16632 19796 16638 19848
rect 17034 19796 17040 19848
rect 17092 19836 17098 19848
rect 18322 19836 18328 19848
rect 17092 19808 17816 19836
rect 18283 19808 18328 19836
rect 17092 19796 17098 19808
rect 16482 19768 16488 19780
rect 15488 19740 16488 19768
rect 15856 19712 15884 19740
rect 16482 19728 16488 19740
rect 16540 19728 16546 19780
rect 14642 19700 14648 19712
rect 13004 19672 14648 19700
rect 14642 19660 14648 19672
rect 14700 19660 14706 19712
rect 15102 19660 15108 19712
rect 15160 19700 15166 19712
rect 15286 19700 15292 19712
rect 15160 19672 15292 19700
rect 15160 19660 15166 19672
rect 15286 19660 15292 19672
rect 15344 19660 15350 19712
rect 15838 19660 15844 19712
rect 15896 19660 15902 19712
rect 16574 19660 16580 19712
rect 16632 19700 16638 19712
rect 16758 19700 16764 19712
rect 16632 19672 16764 19700
rect 16632 19660 16638 19672
rect 16758 19660 16764 19672
rect 16816 19700 16822 19712
rect 17678 19700 17684 19712
rect 16816 19672 17684 19700
rect 16816 19660 16822 19672
rect 17678 19660 17684 19672
rect 17736 19660 17742 19712
rect 17788 19700 17816 19808
rect 18322 19796 18328 19808
rect 18380 19796 18386 19848
rect 18601 19839 18659 19845
rect 18601 19805 18613 19839
rect 18647 19836 18659 19839
rect 19150 19836 19156 19848
rect 18647 19808 19156 19836
rect 18647 19805 18659 19808
rect 18601 19799 18659 19805
rect 19150 19796 19156 19808
rect 19208 19796 19214 19848
rect 19245 19839 19303 19845
rect 19245 19805 19257 19839
rect 19291 19805 19303 19839
rect 19426 19836 19432 19848
rect 19387 19808 19432 19836
rect 19245 19799 19303 19805
rect 19260 19700 19288 19799
rect 19426 19796 19432 19808
rect 19484 19796 19490 19848
rect 19978 19796 19984 19848
rect 20036 19836 20042 19848
rect 20272 19845 20300 19944
rect 22554 19932 22560 19984
rect 22612 19932 22618 19984
rect 25976 19972 26004 20012
rect 26326 20000 26332 20012
rect 26384 20000 26390 20052
rect 23492 19944 26004 19972
rect 22094 19864 22100 19916
rect 22152 19904 22158 19916
rect 22152 19876 22416 19904
rect 22152 19864 22158 19876
rect 20165 19839 20223 19845
rect 20165 19836 20177 19839
rect 20036 19808 20177 19836
rect 20036 19796 20042 19808
rect 20165 19805 20177 19808
rect 20211 19805 20223 19839
rect 20165 19799 20223 19805
rect 20257 19839 20315 19845
rect 20257 19805 20269 19839
rect 20303 19805 20315 19839
rect 20257 19799 20315 19805
rect 20346 19796 20352 19848
rect 20404 19836 20410 19848
rect 20533 19839 20591 19845
rect 20404 19808 20449 19836
rect 20404 19796 20410 19808
rect 20533 19805 20545 19839
rect 20579 19836 20591 19839
rect 22278 19836 22284 19848
rect 20579 19808 22284 19836
rect 20579 19805 20591 19808
rect 20533 19799 20591 19805
rect 22278 19796 22284 19808
rect 22336 19796 22342 19848
rect 22388 19836 22416 19876
rect 22572 19845 22600 19932
rect 23106 19864 23112 19916
rect 23164 19904 23170 19916
rect 23492 19913 23520 19944
rect 23477 19907 23535 19913
rect 23477 19904 23489 19907
rect 23164 19876 23489 19904
rect 23164 19864 23170 19876
rect 23477 19873 23489 19876
rect 23523 19873 23535 19907
rect 23477 19867 23535 19873
rect 23566 19864 23572 19916
rect 23624 19904 23630 19916
rect 24762 19904 24768 19916
rect 23624 19876 24768 19904
rect 23624 19864 23630 19876
rect 24762 19864 24768 19876
rect 24820 19864 24826 19916
rect 25222 19864 25228 19916
rect 25280 19904 25286 19916
rect 25317 19907 25375 19913
rect 25317 19904 25329 19907
rect 25280 19876 25329 19904
rect 25280 19864 25286 19876
rect 25317 19873 25329 19876
rect 25363 19873 25375 19907
rect 25958 19904 25964 19916
rect 25919 19876 25964 19904
rect 25317 19867 25375 19873
rect 25958 19864 25964 19876
rect 26016 19864 26022 19916
rect 22465 19839 22523 19845
rect 22465 19836 22477 19839
rect 22388 19808 22477 19836
rect 22465 19805 22477 19808
rect 22511 19805 22523 19839
rect 22465 19799 22523 19805
rect 22557 19839 22615 19845
rect 22557 19805 22569 19839
rect 22603 19805 22615 19839
rect 22557 19799 22615 19805
rect 22646 19796 22652 19848
rect 22704 19836 22710 19848
rect 22833 19839 22891 19845
rect 22704 19808 22749 19836
rect 22704 19796 22710 19808
rect 22833 19805 22845 19839
rect 22879 19805 22891 19839
rect 22833 19799 22891 19805
rect 23661 19839 23719 19845
rect 23661 19805 23673 19839
rect 23707 19836 23719 19839
rect 24210 19836 24216 19848
rect 23707 19808 24216 19836
rect 23707 19805 23719 19808
rect 23661 19799 23719 19805
rect 21177 19771 21235 19777
rect 21177 19737 21189 19771
rect 21223 19768 21235 19771
rect 22186 19768 22192 19780
rect 21223 19740 22192 19768
rect 21223 19737 21235 19740
rect 21177 19731 21235 19737
rect 22186 19728 22192 19740
rect 22244 19728 22250 19780
rect 22296 19768 22324 19796
rect 22848 19768 22876 19799
rect 24210 19796 24216 19808
rect 24268 19796 24274 19848
rect 24302 19796 24308 19848
rect 24360 19836 24366 19848
rect 24486 19836 24492 19848
rect 24360 19808 24492 19836
rect 24360 19796 24366 19808
rect 24486 19796 24492 19808
rect 24544 19796 24550 19848
rect 26228 19839 26286 19845
rect 26228 19805 26240 19839
rect 26274 19836 26286 19839
rect 27246 19836 27252 19848
rect 26274 19808 27252 19836
rect 26274 19805 26286 19808
rect 26228 19799 26286 19805
rect 27246 19796 27252 19808
rect 27304 19796 27310 19848
rect 25866 19768 25872 19780
rect 22296 19740 22876 19768
rect 25240 19740 25872 19768
rect 25240 19712 25268 19740
rect 25866 19728 25872 19740
rect 25924 19728 25930 19780
rect 17788 19672 19288 19700
rect 19429 19703 19487 19709
rect 19429 19669 19441 19703
rect 19475 19700 19487 19703
rect 19794 19700 19800 19712
rect 19475 19672 19800 19700
rect 19475 19669 19487 19672
rect 19429 19663 19487 19669
rect 19794 19660 19800 19672
rect 19852 19660 19858 19712
rect 20622 19660 20628 19712
rect 20680 19700 20686 19712
rect 21377 19703 21435 19709
rect 21377 19700 21389 19703
rect 20680 19672 21389 19700
rect 20680 19660 20686 19672
rect 21377 19669 21389 19672
rect 21423 19669 21435 19703
rect 21377 19663 21435 19669
rect 21545 19703 21603 19709
rect 21545 19669 21557 19703
rect 21591 19700 21603 19703
rect 23290 19700 23296 19712
rect 21591 19672 23296 19700
rect 21591 19669 21603 19672
rect 21545 19663 21603 19669
rect 23290 19660 23296 19672
rect 23348 19660 23354 19712
rect 24762 19700 24768 19712
rect 24723 19672 24768 19700
rect 24762 19660 24768 19672
rect 24820 19660 24826 19712
rect 25038 19660 25044 19712
rect 25096 19700 25102 19712
rect 25133 19703 25191 19709
rect 25133 19700 25145 19703
rect 25096 19672 25145 19700
rect 25096 19660 25102 19672
rect 25133 19669 25145 19672
rect 25179 19669 25191 19703
rect 25133 19663 25191 19669
rect 25222 19660 25228 19712
rect 25280 19700 25286 19712
rect 25280 19672 25325 19700
rect 25280 19660 25286 19672
rect 25590 19660 25596 19712
rect 25648 19700 25654 19712
rect 27341 19703 27399 19709
rect 27341 19700 27353 19703
rect 25648 19672 27353 19700
rect 25648 19660 25654 19672
rect 27341 19669 27353 19672
rect 27387 19669 27399 19703
rect 27341 19663 27399 19669
rect 1104 19610 28060 19632
rect 1104 19558 9935 19610
rect 9987 19558 9999 19610
rect 10051 19558 10063 19610
rect 10115 19558 10127 19610
rect 10179 19558 10191 19610
rect 10243 19558 18920 19610
rect 18972 19558 18984 19610
rect 19036 19558 19048 19610
rect 19100 19558 19112 19610
rect 19164 19558 19176 19610
rect 19228 19558 28060 19610
rect 1104 19536 28060 19558
rect 1673 19499 1731 19505
rect 1673 19465 1685 19499
rect 1719 19496 1731 19499
rect 1854 19496 1860 19508
rect 1719 19468 1860 19496
rect 1719 19465 1731 19468
rect 1673 19459 1731 19465
rect 1854 19456 1860 19468
rect 1912 19456 1918 19508
rect 3602 19496 3608 19508
rect 2332 19468 3608 19496
rect 2332 19369 2360 19468
rect 3602 19456 3608 19468
rect 3660 19456 3666 19508
rect 4430 19456 4436 19508
rect 4488 19496 4494 19508
rect 4890 19496 4896 19508
rect 4488 19468 4896 19496
rect 4488 19456 4494 19468
rect 4890 19456 4896 19468
rect 4948 19456 4954 19508
rect 4985 19499 5043 19505
rect 4985 19465 4997 19499
rect 5031 19496 5043 19499
rect 6086 19496 6092 19508
rect 5031 19468 6092 19496
rect 5031 19465 5043 19468
rect 4985 19459 5043 19465
rect 6086 19456 6092 19468
rect 6144 19456 6150 19508
rect 6917 19499 6975 19505
rect 6917 19465 6929 19499
rect 6963 19496 6975 19499
rect 7282 19496 7288 19508
rect 6963 19468 7288 19496
rect 6963 19465 6975 19468
rect 6917 19459 6975 19465
rect 7282 19456 7288 19468
rect 7340 19456 7346 19508
rect 8294 19456 8300 19508
rect 8352 19496 8358 19508
rect 13262 19496 13268 19508
rect 8352 19468 13268 19496
rect 8352 19456 8358 19468
rect 13262 19456 13268 19468
rect 13320 19456 13326 19508
rect 13446 19456 13452 19508
rect 13504 19496 13510 19508
rect 13541 19499 13599 19505
rect 13541 19496 13553 19499
rect 13504 19468 13553 19496
rect 13504 19456 13510 19468
rect 13541 19465 13553 19468
rect 13587 19465 13599 19499
rect 13541 19459 13599 19465
rect 13998 19456 14004 19508
rect 14056 19456 14062 19508
rect 14458 19456 14464 19508
rect 14516 19496 14522 19508
rect 15930 19496 15936 19508
rect 14516 19468 15936 19496
rect 14516 19456 14522 19468
rect 15930 19456 15936 19468
rect 15988 19496 15994 19508
rect 16117 19499 16175 19505
rect 16117 19496 16129 19499
rect 15988 19468 16129 19496
rect 15988 19456 15994 19468
rect 16117 19465 16129 19468
rect 16163 19465 16175 19499
rect 16117 19459 16175 19465
rect 16761 19499 16819 19505
rect 16761 19465 16773 19499
rect 16807 19496 16819 19499
rect 17678 19496 17684 19508
rect 16807 19468 17684 19496
rect 16807 19465 16819 19468
rect 16761 19459 16819 19465
rect 17678 19456 17684 19468
rect 17736 19456 17742 19508
rect 18141 19499 18199 19505
rect 18141 19465 18153 19499
rect 18187 19496 18199 19499
rect 18322 19496 18328 19508
rect 18187 19468 18328 19496
rect 18187 19465 18199 19468
rect 18141 19459 18199 19465
rect 18322 19456 18328 19468
rect 18380 19456 18386 19508
rect 18616 19468 18920 19496
rect 3872 19431 3930 19437
rect 2424 19400 3832 19428
rect 1857 19363 1915 19369
rect 1857 19329 1869 19363
rect 1903 19360 1915 19363
rect 2317 19363 2375 19369
rect 1903 19332 2268 19360
rect 1903 19329 1915 19332
rect 1857 19323 1915 19329
rect 2240 19292 2268 19332
rect 2317 19329 2329 19363
rect 2363 19329 2375 19363
rect 2317 19323 2375 19329
rect 2424 19292 2452 19400
rect 2498 19320 2504 19372
rect 2556 19360 2562 19372
rect 2961 19363 3019 19369
rect 2961 19360 2973 19363
rect 2556 19332 2601 19360
rect 2746 19332 2973 19360
rect 2556 19320 2562 19332
rect 2240 19264 2452 19292
rect 2746 19236 2774 19332
rect 2961 19329 2973 19332
rect 3007 19329 3019 19363
rect 3142 19360 3148 19372
rect 3103 19332 3148 19360
rect 2961 19323 3019 19329
rect 3142 19320 3148 19332
rect 3200 19320 3206 19372
rect 3602 19360 3608 19372
rect 3563 19332 3608 19360
rect 3602 19320 3608 19332
rect 3660 19320 3666 19372
rect 3804 19360 3832 19400
rect 3872 19397 3884 19431
rect 3918 19428 3930 19431
rect 3918 19400 7787 19428
rect 3918 19397 3930 19400
rect 3872 19391 3930 19397
rect 5537 19363 5595 19369
rect 3804 19332 5488 19360
rect 5460 19292 5488 19332
rect 5537 19329 5549 19363
rect 5583 19360 5595 19363
rect 5583 19332 6040 19360
rect 5583 19329 5595 19332
rect 5537 19323 5595 19329
rect 6012 19292 6040 19332
rect 6086 19320 6092 19372
rect 6144 19360 6150 19372
rect 6825 19363 6883 19369
rect 6825 19360 6837 19363
rect 6144 19332 6837 19360
rect 6144 19320 6150 19332
rect 6825 19329 6837 19332
rect 6871 19329 6883 19363
rect 6825 19323 6883 19329
rect 7558 19292 7564 19304
rect 5460 19264 5580 19292
rect 6012 19264 7564 19292
rect 2682 19184 2688 19236
rect 2740 19196 2774 19236
rect 2740 19184 2746 19196
rect 5258 19184 5264 19236
rect 5316 19184 5322 19236
rect 5552 19224 5580 19264
rect 7558 19252 7564 19264
rect 7616 19252 7622 19304
rect 7282 19224 7288 19236
rect 5552 19196 7288 19224
rect 7282 19184 7288 19196
rect 7340 19184 7346 19236
rect 2409 19159 2467 19165
rect 2409 19125 2421 19159
rect 2455 19156 2467 19159
rect 2590 19156 2596 19168
rect 2455 19128 2596 19156
rect 2455 19125 2467 19128
rect 2409 19119 2467 19125
rect 2590 19116 2596 19128
rect 2648 19116 2654 19168
rect 2961 19159 3019 19165
rect 2961 19125 2973 19159
rect 3007 19156 3019 19159
rect 4614 19156 4620 19168
rect 3007 19128 4620 19156
rect 3007 19125 3019 19128
rect 2961 19119 3019 19125
rect 4614 19116 4620 19128
rect 4672 19116 4678 19168
rect 5276 19156 5304 19184
rect 5629 19159 5687 19165
rect 5629 19156 5641 19159
rect 5276 19128 5641 19156
rect 5629 19125 5641 19128
rect 5675 19156 5687 19159
rect 6914 19156 6920 19168
rect 5675 19128 6920 19156
rect 5675 19125 5687 19128
rect 5629 19119 5687 19125
rect 6914 19116 6920 19128
rect 6972 19116 6978 19168
rect 7006 19116 7012 19168
rect 7064 19156 7070 19168
rect 7653 19159 7711 19165
rect 7653 19156 7665 19159
rect 7064 19128 7665 19156
rect 7064 19116 7070 19128
rect 7653 19125 7665 19128
rect 7699 19125 7711 19159
rect 7759 19156 7787 19400
rect 8772 19400 9168 19428
rect 7834 19320 7840 19372
rect 7892 19350 7898 19372
rect 7929 19363 7987 19369
rect 7929 19350 7941 19363
rect 7892 19329 7941 19350
rect 7975 19329 7987 19363
rect 7892 19323 7987 19329
rect 8021 19363 8079 19369
rect 8021 19329 8033 19363
rect 8067 19329 8079 19363
rect 8021 19323 8079 19329
rect 7892 19322 7972 19323
rect 7892 19320 7898 19322
rect 8036 19292 8064 19323
rect 8110 19320 8116 19372
rect 8168 19360 8174 19372
rect 8772 19369 8800 19400
rect 9030 19369 9036 19372
rect 8297 19363 8355 19369
rect 8168 19332 8213 19360
rect 8168 19320 8174 19332
rect 8297 19329 8309 19363
rect 8343 19360 8355 19363
rect 8757 19363 8815 19369
rect 8343 19332 8432 19360
rect 8343 19329 8355 19332
rect 8297 19323 8355 19329
rect 8404 19304 8432 19332
rect 8757 19329 8769 19363
rect 8803 19329 8815 19363
rect 9024 19360 9036 19369
rect 8991 19332 9036 19360
rect 8757 19323 8815 19329
rect 9024 19323 9036 19332
rect 9030 19320 9036 19323
rect 9088 19320 9094 19372
rect 9140 19360 9168 19400
rect 9582 19388 9588 19440
rect 9640 19428 9646 19440
rect 9640 19400 10640 19428
rect 9640 19388 9646 19400
rect 10226 19360 10232 19372
rect 9140 19332 10232 19360
rect 10226 19320 10232 19332
rect 10284 19320 10290 19372
rect 8036 19264 8294 19292
rect 8266 19224 8294 19264
rect 8386 19252 8392 19304
rect 8444 19252 8450 19304
rect 10612 19292 10640 19400
rect 10686 19388 10692 19440
rect 10744 19428 10750 19440
rect 10962 19428 10968 19440
rect 10744 19400 10968 19428
rect 10744 19388 10750 19400
rect 10962 19388 10968 19400
rect 11020 19388 11026 19440
rect 12986 19428 12992 19440
rect 12176 19400 12992 19428
rect 11606 19320 11612 19372
rect 11664 19360 11670 19372
rect 11747 19363 11805 19369
rect 11747 19360 11759 19363
rect 11664 19332 11759 19360
rect 11664 19320 11670 19332
rect 11747 19329 11759 19332
rect 11793 19329 11805 19363
rect 11882 19360 11888 19372
rect 11843 19332 11888 19360
rect 11747 19323 11805 19329
rect 11882 19320 11888 19332
rect 11940 19320 11946 19372
rect 11977 19363 12035 19369
rect 11977 19329 11989 19363
rect 12023 19360 12035 19363
rect 12066 19360 12072 19372
rect 12023 19332 12072 19360
rect 12023 19329 12035 19332
rect 11977 19323 12035 19329
rect 12066 19320 12072 19332
rect 12124 19320 12130 19372
rect 12176 19369 12204 19400
rect 12986 19388 12992 19400
rect 13044 19388 13050 19440
rect 12161 19363 12219 19369
rect 12161 19329 12173 19363
rect 12207 19329 12219 19363
rect 12161 19323 12219 19329
rect 12176 19292 12204 19323
rect 12618 19320 12624 19372
rect 12676 19360 12682 19372
rect 12676 19332 12721 19360
rect 12676 19320 12682 19332
rect 12802 19320 12808 19372
rect 12860 19360 12866 19372
rect 13814 19369 13820 19372
rect 13797 19363 13820 19369
rect 12860 19332 12905 19360
rect 12860 19320 12866 19332
rect 13797 19329 13809 19363
rect 13797 19323 13820 19329
rect 13814 19320 13820 19323
rect 13872 19320 13878 19372
rect 14016 19369 14044 19456
rect 16298 19428 16304 19440
rect 14752 19400 16304 19428
rect 13906 19363 13964 19369
rect 13906 19329 13918 19363
rect 13952 19329 13964 19363
rect 13906 19323 13964 19329
rect 14001 19363 14059 19369
rect 14001 19329 14013 19363
rect 14047 19329 14059 19363
rect 14182 19360 14188 19372
rect 14143 19332 14188 19360
rect 14001 19323 14059 19329
rect 10612 19264 12204 19292
rect 12434 19252 12440 19304
rect 12492 19292 12498 19304
rect 12989 19295 13047 19301
rect 12989 19292 13001 19295
rect 12492 19264 13001 19292
rect 12492 19252 12498 19264
rect 12989 19261 13001 19264
rect 13035 19261 13047 19295
rect 13921 19292 13949 19323
rect 14182 19320 14188 19332
rect 14240 19320 14246 19372
rect 14752 19369 14780 19400
rect 16298 19388 16304 19400
rect 16356 19388 16362 19440
rect 18616 19428 18644 19468
rect 16592 19400 18644 19428
rect 18892 19428 18920 19468
rect 19610 19456 19616 19508
rect 19668 19496 19674 19508
rect 20622 19496 20628 19508
rect 19668 19468 20628 19496
rect 19668 19456 19674 19468
rect 20622 19456 20628 19468
rect 20680 19496 20686 19508
rect 22281 19499 22339 19505
rect 20680 19468 22094 19496
rect 20680 19456 20686 19468
rect 20165 19431 20223 19437
rect 20165 19428 20177 19431
rect 18892 19400 20177 19428
rect 14737 19363 14795 19369
rect 14737 19329 14749 19363
rect 14783 19329 14795 19363
rect 14737 19323 14795 19329
rect 14826 19320 14832 19372
rect 14884 19360 14890 19372
rect 14993 19363 15051 19369
rect 14993 19360 15005 19363
rect 14884 19332 15005 19360
rect 14884 19320 14890 19332
rect 14993 19329 15005 19332
rect 15039 19329 15051 19363
rect 14993 19323 15051 19329
rect 15746 19294 15752 19346
rect 15804 19334 15810 19346
rect 15804 19306 15900 19334
rect 16114 19320 16120 19372
rect 16172 19360 16178 19372
rect 16592 19360 16620 19400
rect 20165 19397 20177 19400
rect 20211 19428 20223 19431
rect 21085 19431 21143 19437
rect 21085 19428 21097 19431
rect 20211 19400 21097 19428
rect 20211 19397 20223 19400
rect 20165 19391 20223 19397
rect 21085 19397 21097 19400
rect 21131 19397 21143 19431
rect 21085 19391 21143 19397
rect 16172 19332 16620 19360
rect 16669 19363 16727 19369
rect 16172 19320 16178 19332
rect 16669 19329 16681 19363
rect 16715 19360 16727 19363
rect 16758 19360 16764 19372
rect 16715 19332 16764 19360
rect 16715 19329 16727 19332
rect 16669 19323 16727 19329
rect 16758 19320 16764 19332
rect 16816 19320 16822 19372
rect 17402 19360 17408 19372
rect 17363 19332 17408 19360
rect 17402 19320 17408 19332
rect 17460 19320 17466 19372
rect 17589 19363 17647 19369
rect 17589 19329 17601 19363
rect 17635 19360 17647 19363
rect 17862 19360 17868 19372
rect 17635 19332 17868 19360
rect 17635 19329 17647 19332
rect 17589 19323 17647 19329
rect 17862 19320 17868 19332
rect 17920 19320 17926 19372
rect 17957 19363 18015 19369
rect 17957 19329 17969 19363
rect 18003 19360 18015 19363
rect 18690 19360 18696 19372
rect 18003 19332 18696 19360
rect 18003 19329 18015 19332
rect 17957 19323 18015 19329
rect 18690 19320 18696 19332
rect 18748 19320 18754 19372
rect 18874 19360 18880 19372
rect 18835 19332 18880 19360
rect 18874 19320 18880 19332
rect 18932 19320 18938 19372
rect 19061 19363 19119 19369
rect 19061 19329 19073 19363
rect 19107 19329 19119 19363
rect 19061 19323 19119 19329
rect 19245 19363 19303 19369
rect 19245 19329 19257 19363
rect 19291 19360 19303 19363
rect 19429 19363 19487 19369
rect 19291 19332 19380 19360
rect 19291 19329 19303 19332
rect 19245 19323 19303 19329
rect 15804 19294 15810 19306
rect 12989 19255 13047 19261
rect 13740 19264 13949 19292
rect 15872 19292 15900 19306
rect 16482 19292 16488 19304
rect 15872 19264 16488 19292
rect 13740 19236 13768 19264
rect 16482 19252 16488 19264
rect 16540 19252 16546 19304
rect 17218 19252 17224 19304
rect 17276 19292 17282 19304
rect 17681 19295 17739 19301
rect 17681 19292 17693 19295
rect 17276 19264 17693 19292
rect 17276 19252 17282 19264
rect 17681 19261 17693 19264
rect 17727 19261 17739 19295
rect 17681 19255 17739 19261
rect 17773 19295 17831 19301
rect 17773 19261 17785 19295
rect 17819 19292 17831 19295
rect 18322 19292 18328 19304
rect 17819 19264 18328 19292
rect 17819 19261 17831 19264
rect 17773 19255 17831 19261
rect 18322 19252 18328 19264
rect 18380 19252 18386 19304
rect 19076 19292 19104 19323
rect 18524 19264 19104 19292
rect 19153 19295 19211 19301
rect 8570 19224 8576 19236
rect 8266 19196 8576 19224
rect 8570 19184 8576 19196
rect 8628 19184 8634 19236
rect 10318 19224 10324 19236
rect 10152 19196 10324 19224
rect 8110 19156 8116 19168
rect 7759 19128 8116 19156
rect 7653 19119 7711 19125
rect 8110 19116 8116 19128
rect 8168 19116 8174 19168
rect 9950 19116 9956 19168
rect 10008 19156 10014 19168
rect 10152 19165 10180 19196
rect 10318 19184 10324 19196
rect 10376 19184 10382 19236
rect 12526 19224 12532 19236
rect 12176 19196 12532 19224
rect 10137 19159 10195 19165
rect 10137 19156 10149 19159
rect 10008 19128 10149 19156
rect 10008 19116 10014 19128
rect 10137 19125 10149 19128
rect 10183 19125 10195 19159
rect 10137 19119 10195 19125
rect 10226 19116 10232 19168
rect 10284 19156 10290 19168
rect 10778 19156 10784 19168
rect 10284 19128 10784 19156
rect 10284 19116 10290 19128
rect 10778 19116 10784 19128
rect 10836 19116 10842 19168
rect 11514 19156 11520 19168
rect 11475 19128 11520 19156
rect 11514 19116 11520 19128
rect 11572 19116 11578 19168
rect 11882 19116 11888 19168
rect 11940 19156 11946 19168
rect 12176 19156 12204 19196
rect 12526 19184 12532 19196
rect 12584 19184 12590 19236
rect 13722 19184 13728 19236
rect 13780 19184 13786 19236
rect 14458 19224 14464 19236
rect 14005 19196 14464 19224
rect 11940 19128 12204 19156
rect 11940 19116 11946 19128
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 13078 19156 13084 19168
rect 12492 19128 13084 19156
rect 12492 19116 12498 19128
rect 13078 19116 13084 19128
rect 13136 19116 13142 19168
rect 13354 19116 13360 19168
rect 13412 19156 13418 19168
rect 14005 19156 14033 19196
rect 14458 19184 14464 19196
rect 14516 19184 14522 19236
rect 17862 19184 17868 19236
rect 17920 19224 17926 19236
rect 18524 19224 18552 19264
rect 19153 19261 19165 19295
rect 19199 19261 19211 19295
rect 19153 19255 19211 19261
rect 17920 19196 18552 19224
rect 17920 19184 17926 19196
rect 19058 19184 19064 19236
rect 19116 19224 19122 19236
rect 19168 19224 19196 19255
rect 19116 19196 19196 19224
rect 19116 19184 19122 19196
rect 13412 19128 14033 19156
rect 13412 19116 13418 19128
rect 14090 19116 14096 19168
rect 14148 19156 14154 19168
rect 16482 19156 16488 19168
rect 14148 19128 16488 19156
rect 14148 19116 14154 19128
rect 16482 19116 16488 19128
rect 16540 19116 16546 19168
rect 18322 19116 18328 19168
rect 18380 19156 18386 19168
rect 19352 19156 19380 19332
rect 19429 19329 19441 19363
rect 19475 19360 19487 19363
rect 20070 19360 20076 19372
rect 19475 19332 20076 19360
rect 19475 19329 19487 19332
rect 19429 19323 19487 19329
rect 20070 19320 20076 19332
rect 20128 19320 20134 19372
rect 22066 19360 22094 19468
rect 22281 19465 22293 19499
rect 22327 19496 22339 19499
rect 22370 19496 22376 19508
rect 22327 19468 22376 19496
rect 22327 19465 22339 19468
rect 22281 19459 22339 19465
rect 22370 19456 22376 19468
rect 22428 19456 22434 19508
rect 23014 19456 23020 19508
rect 23072 19496 23078 19508
rect 23293 19499 23351 19505
rect 23293 19496 23305 19499
rect 23072 19468 23305 19496
rect 23072 19456 23078 19468
rect 23293 19465 23305 19468
rect 23339 19465 23351 19499
rect 25685 19499 25743 19505
rect 23293 19459 23351 19465
rect 23952 19468 24624 19496
rect 22186 19388 22192 19440
rect 22244 19428 22250 19440
rect 22244 19400 22600 19428
rect 22244 19388 22250 19400
rect 22572 19369 22600 19400
rect 23198 19388 23204 19440
rect 23256 19428 23262 19440
rect 23256 19400 23520 19428
rect 23256 19388 23262 19400
rect 22465 19363 22523 19369
rect 22465 19360 22477 19363
rect 22066 19332 22477 19360
rect 22465 19329 22477 19332
rect 22511 19329 22523 19363
rect 22465 19323 22523 19329
rect 22557 19363 22615 19369
rect 22557 19329 22569 19363
rect 22603 19329 22615 19363
rect 22557 19323 22615 19329
rect 22646 19320 22652 19372
rect 22704 19350 22710 19372
rect 22741 19363 22799 19369
rect 22741 19350 22753 19363
rect 22704 19329 22753 19350
rect 22787 19329 22799 19363
rect 22704 19323 22799 19329
rect 22833 19364 22891 19369
rect 22833 19363 23060 19364
rect 22833 19329 22845 19363
rect 22879 19360 23060 19363
rect 23290 19360 23296 19372
rect 22879 19336 23296 19360
rect 22879 19329 22891 19336
rect 23032 19332 23296 19336
rect 22833 19323 22891 19329
rect 22704 19322 22784 19323
rect 22704 19320 22710 19322
rect 23290 19320 23296 19332
rect 23348 19320 23354 19372
rect 23492 19369 23520 19400
rect 23477 19363 23535 19369
rect 23477 19329 23489 19363
rect 23523 19329 23535 19363
rect 23477 19323 23535 19329
rect 23842 19320 23848 19372
rect 23900 19360 23906 19372
rect 23952 19369 23980 19468
rect 24118 19428 24124 19440
rect 24079 19400 24124 19428
rect 24118 19388 24124 19400
rect 24176 19388 24182 19440
rect 24486 19428 24492 19440
rect 24320 19400 24492 19428
rect 24320 19369 24348 19400
rect 24486 19388 24492 19400
rect 24544 19388 24550 19440
rect 23937 19363 23995 19369
rect 23937 19360 23949 19363
rect 23900 19332 23949 19360
rect 23900 19320 23906 19332
rect 23937 19329 23949 19332
rect 23983 19329 23995 19363
rect 24213 19363 24271 19369
rect 24213 19360 24225 19363
rect 23937 19323 23995 19329
rect 24136 19329 24225 19360
rect 24259 19329 24271 19363
rect 24136 19323 24271 19329
rect 24305 19363 24363 19369
rect 24305 19329 24317 19363
rect 24351 19329 24363 19363
rect 24596 19358 24624 19468
rect 25685 19465 25697 19499
rect 25731 19465 25743 19499
rect 25685 19459 25743 19465
rect 26237 19499 26295 19505
rect 26237 19465 26249 19499
rect 26283 19496 26295 19499
rect 26418 19496 26424 19508
rect 26283 19468 26424 19496
rect 26283 19465 26295 19468
rect 26237 19459 26295 19465
rect 24762 19388 24768 19440
rect 24820 19428 24826 19440
rect 25317 19431 25375 19437
rect 25317 19428 25329 19431
rect 24820 19400 25329 19428
rect 24820 19388 24826 19400
rect 25317 19397 25329 19400
rect 25363 19397 25375 19431
rect 25700 19428 25728 19459
rect 26418 19456 26424 19468
rect 26476 19456 26482 19508
rect 26878 19456 26884 19508
rect 26936 19496 26942 19508
rect 27341 19499 27399 19505
rect 27341 19496 27353 19499
rect 26936 19468 27353 19496
rect 26936 19456 26942 19468
rect 27341 19465 27353 19468
rect 27387 19465 27399 19499
rect 27341 19459 27399 19465
rect 25700 19400 27200 19428
rect 25317 19391 25375 19397
rect 25133 19363 25191 19369
rect 25133 19360 25145 19363
rect 24657 19358 25145 19360
rect 24596 19332 25145 19358
rect 24596 19330 24685 19332
rect 24305 19323 24363 19329
rect 25133 19329 25145 19332
rect 25179 19329 25191 19363
rect 25409 19363 25467 19369
rect 25409 19360 25421 19363
rect 25133 19323 25191 19329
rect 25332 19332 25421 19360
rect 24136 19306 24256 19323
rect 21269 19295 21327 19301
rect 21269 19261 21281 19295
rect 21315 19292 21327 19295
rect 23658 19292 23664 19304
rect 21315 19264 23664 19292
rect 21315 19261 21327 19264
rect 21269 19255 21327 19261
rect 23658 19252 23664 19264
rect 23716 19252 23722 19304
rect 22646 19184 22652 19236
rect 22704 19224 22710 19236
rect 23106 19224 23112 19236
rect 22704 19196 23112 19224
rect 22704 19184 22710 19196
rect 23106 19184 23112 19196
rect 23164 19184 23170 19236
rect 23566 19184 23572 19236
rect 23624 19224 23630 19236
rect 23842 19224 23848 19236
rect 23624 19196 23848 19224
rect 23624 19184 23630 19196
rect 23842 19184 23848 19196
rect 23900 19184 23906 19236
rect 24228 19224 24256 19306
rect 25332 19304 25360 19332
rect 25409 19329 25421 19332
rect 25455 19329 25467 19363
rect 25409 19323 25467 19329
rect 25501 19363 25559 19369
rect 25501 19329 25513 19363
rect 25547 19360 25559 19363
rect 25774 19360 25780 19372
rect 25547 19332 25780 19360
rect 25547 19329 25559 19332
rect 25501 19323 25559 19329
rect 25774 19320 25780 19332
rect 25832 19320 25838 19372
rect 26050 19320 26056 19372
rect 26108 19360 26114 19372
rect 27172 19369 27200 19400
rect 26421 19363 26479 19369
rect 26421 19360 26433 19363
rect 26108 19332 26433 19360
rect 26108 19320 26114 19332
rect 26421 19329 26433 19332
rect 26467 19329 26479 19363
rect 26421 19323 26479 19329
rect 27157 19363 27215 19369
rect 27157 19329 27169 19363
rect 27203 19329 27215 19363
rect 27157 19323 27215 19329
rect 25314 19252 25320 19304
rect 25372 19252 25378 19304
rect 26326 19252 26332 19304
rect 26384 19292 26390 19304
rect 26973 19295 27031 19301
rect 26973 19292 26985 19295
rect 26384 19264 26985 19292
rect 26384 19252 26390 19264
rect 26973 19261 26985 19264
rect 27019 19261 27031 19295
rect 26973 19255 27031 19261
rect 24228 19196 24624 19224
rect 19610 19156 19616 19168
rect 18380 19128 19380 19156
rect 19571 19128 19616 19156
rect 18380 19116 18386 19128
rect 19610 19116 19616 19128
rect 19668 19116 19674 19168
rect 20070 19116 20076 19168
rect 20128 19156 20134 19168
rect 20257 19159 20315 19165
rect 20257 19156 20269 19159
rect 20128 19128 20269 19156
rect 20128 19116 20134 19128
rect 20257 19125 20269 19128
rect 20303 19125 20315 19159
rect 20257 19119 20315 19125
rect 22278 19116 22284 19168
rect 22336 19156 22342 19168
rect 24026 19156 24032 19168
rect 22336 19128 24032 19156
rect 22336 19116 22342 19128
rect 24026 19116 24032 19128
rect 24084 19116 24090 19168
rect 24210 19116 24216 19168
rect 24268 19156 24274 19168
rect 24489 19159 24547 19165
rect 24489 19156 24501 19159
rect 24268 19128 24501 19156
rect 24268 19116 24274 19128
rect 24489 19125 24501 19128
rect 24535 19125 24547 19159
rect 24596 19156 24624 19196
rect 24946 19156 24952 19168
rect 24596 19128 24952 19156
rect 24489 19119 24547 19125
rect 24946 19116 24952 19128
rect 25004 19116 25010 19168
rect 25038 19116 25044 19168
rect 25096 19156 25102 19168
rect 25314 19156 25320 19168
rect 25096 19128 25320 19156
rect 25096 19116 25102 19128
rect 25314 19116 25320 19128
rect 25372 19116 25378 19168
rect 1104 19066 28060 19088
rect 1104 19014 5442 19066
rect 5494 19014 5506 19066
rect 5558 19014 5570 19066
rect 5622 19014 5634 19066
rect 5686 19014 5698 19066
rect 5750 19014 14428 19066
rect 14480 19014 14492 19066
rect 14544 19014 14556 19066
rect 14608 19014 14620 19066
rect 14672 19014 14684 19066
rect 14736 19014 23413 19066
rect 23465 19014 23477 19066
rect 23529 19014 23541 19066
rect 23593 19014 23605 19066
rect 23657 19014 23669 19066
rect 23721 19014 28060 19066
rect 1104 18992 28060 19014
rect 1581 18955 1639 18961
rect 1581 18921 1593 18955
rect 1627 18952 1639 18955
rect 1627 18924 3556 18952
rect 1627 18921 1639 18924
rect 1581 18915 1639 18921
rect 2409 18887 2467 18893
rect 2409 18853 2421 18887
rect 2455 18884 2467 18887
rect 3528 18884 3556 18924
rect 3602 18912 3608 18964
rect 3660 18952 3666 18964
rect 4893 18955 4951 18961
rect 4893 18952 4905 18955
rect 3660 18924 4905 18952
rect 3660 18912 3666 18924
rect 4893 18921 4905 18924
rect 4939 18921 4951 18955
rect 8478 18952 8484 18964
rect 4893 18915 4951 18921
rect 5000 18924 8484 18952
rect 5000 18884 5028 18924
rect 8478 18912 8484 18924
rect 8536 18912 8542 18964
rect 9030 18912 9036 18964
rect 9088 18952 9094 18964
rect 9769 18955 9827 18961
rect 9769 18952 9781 18955
rect 9088 18924 9781 18952
rect 9088 18912 9094 18924
rect 9769 18921 9781 18924
rect 9815 18921 9827 18955
rect 11882 18952 11888 18964
rect 9769 18915 9827 18921
rect 9876 18924 11888 18952
rect 6822 18884 6828 18896
rect 2455 18856 3464 18884
rect 3528 18856 5028 18884
rect 6783 18856 6828 18884
rect 2455 18853 2467 18856
rect 2409 18847 2467 18853
rect 3142 18776 3148 18828
rect 3200 18816 3206 18828
rect 3436 18816 3464 18856
rect 6822 18844 6828 18856
rect 6880 18844 6886 18896
rect 6914 18844 6920 18896
rect 6972 18884 6978 18896
rect 9876 18884 9904 18924
rect 11882 18912 11888 18924
rect 11940 18912 11946 18964
rect 13541 18955 13599 18961
rect 13541 18921 13553 18955
rect 13587 18952 13599 18955
rect 13998 18952 14004 18964
rect 13587 18924 14004 18952
rect 13587 18921 13599 18924
rect 13541 18915 13599 18921
rect 13998 18912 14004 18924
rect 14056 18912 14062 18964
rect 14090 18912 14096 18964
rect 14148 18952 14154 18964
rect 14148 18924 16160 18952
rect 14148 18912 14154 18924
rect 10686 18884 10692 18896
rect 6972 18856 9904 18884
rect 9968 18856 10692 18884
rect 6972 18844 6978 18856
rect 7558 18816 7564 18828
rect 3200 18788 3372 18816
rect 3436 18788 5396 18816
rect 7519 18788 7564 18816
rect 3200 18776 3206 18788
rect 1394 18708 1400 18760
rect 1452 18748 1458 18760
rect 1581 18751 1639 18757
rect 1581 18748 1593 18751
rect 1452 18720 1593 18748
rect 1452 18708 1458 18720
rect 1581 18717 1593 18720
rect 1627 18717 1639 18751
rect 1581 18711 1639 18717
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18748 1823 18751
rect 1854 18748 1860 18760
rect 1811 18720 1860 18748
rect 1811 18717 1823 18720
rect 1765 18711 1823 18717
rect 1596 18680 1624 18711
rect 1854 18708 1860 18720
rect 1912 18708 1918 18760
rect 2133 18751 2191 18757
rect 2133 18717 2145 18751
rect 2179 18748 2191 18751
rect 2593 18751 2651 18757
rect 2593 18748 2605 18751
rect 2179 18720 2605 18748
rect 2179 18717 2191 18720
rect 2133 18711 2191 18717
rect 2593 18717 2605 18720
rect 2639 18748 2651 18751
rect 2682 18748 2688 18760
rect 2639 18720 2688 18748
rect 2639 18717 2651 18720
rect 2593 18711 2651 18717
rect 2682 18708 2688 18720
rect 2740 18708 2746 18760
rect 3237 18751 3295 18757
rect 3237 18717 3249 18751
rect 3283 18744 3295 18751
rect 3344 18744 3372 18788
rect 5368 18760 5396 18788
rect 7558 18776 7564 18788
rect 7616 18776 7622 18828
rect 9309 18819 9367 18825
rect 9309 18785 9321 18819
rect 9355 18816 9367 18819
rect 9968 18816 9996 18856
rect 10686 18844 10692 18856
rect 10744 18844 10750 18896
rect 10870 18844 10876 18896
rect 10928 18884 10934 18896
rect 12250 18884 12256 18896
rect 10928 18856 10973 18884
rect 11164 18856 12256 18884
rect 10928 18844 10934 18856
rect 9355 18788 9996 18816
rect 10152 18788 10916 18816
rect 9355 18785 9367 18788
rect 9309 18779 9367 18785
rect 3283 18717 3372 18744
rect 3237 18716 3372 18717
rect 4249 18751 4307 18757
rect 4249 18717 4261 18751
rect 4295 18744 4307 18751
rect 4801 18751 4859 18757
rect 4295 18717 4375 18744
rect 4249 18716 4375 18717
rect 3237 18711 3295 18716
rect 4249 18711 4307 18716
rect 4347 18680 4375 18716
rect 4801 18717 4813 18751
rect 4847 18748 4859 18751
rect 4890 18748 4896 18760
rect 4847 18720 4896 18748
rect 4847 18717 4859 18720
rect 4801 18711 4859 18717
rect 4890 18708 4896 18720
rect 4948 18708 4954 18760
rect 5350 18708 5356 18760
rect 5408 18708 5414 18760
rect 5445 18751 5503 18757
rect 5445 18717 5457 18751
rect 5491 18748 5503 18751
rect 6546 18748 6552 18760
rect 5491 18720 6552 18748
rect 5491 18717 5503 18720
rect 5445 18711 5503 18717
rect 6546 18708 6552 18720
rect 6604 18708 6610 18760
rect 7006 18748 7012 18760
rect 6656 18720 7012 18748
rect 5534 18680 5540 18692
rect 1596 18652 2360 18680
rect 1854 18572 1860 18624
rect 1912 18612 1918 18624
rect 2222 18612 2228 18624
rect 1912 18584 2228 18612
rect 1912 18572 1918 18584
rect 2222 18572 2228 18584
rect 2280 18572 2286 18624
rect 2332 18612 2360 18652
rect 3344 18652 4200 18680
rect 4347 18652 4752 18680
rect 2869 18615 2927 18621
rect 2869 18612 2881 18615
rect 2332 18584 2881 18612
rect 2869 18581 2881 18584
rect 2915 18581 2927 18615
rect 2869 18575 2927 18581
rect 3053 18615 3111 18621
rect 3053 18581 3065 18615
rect 3099 18612 3111 18615
rect 3344 18612 3372 18652
rect 3099 18584 3372 18612
rect 3099 18581 3111 18584
rect 3053 18575 3111 18581
rect 3418 18572 3424 18624
rect 3476 18612 3482 18624
rect 4065 18615 4123 18621
rect 4065 18612 4077 18615
rect 3476 18584 4077 18612
rect 3476 18572 3482 18584
rect 4065 18581 4077 18584
rect 4111 18581 4123 18615
rect 4172 18612 4200 18652
rect 4430 18612 4436 18624
rect 4172 18584 4436 18612
rect 4065 18575 4123 18581
rect 4430 18572 4436 18584
rect 4488 18572 4494 18624
rect 4724 18612 4752 18652
rect 5210 18652 5540 18680
rect 5210 18612 5238 18652
rect 5534 18640 5540 18652
rect 5592 18640 5598 18692
rect 5712 18683 5770 18689
rect 5712 18649 5724 18683
rect 5758 18680 5770 18683
rect 6656 18680 6684 18720
rect 7006 18708 7012 18720
rect 7064 18708 7070 18760
rect 7282 18748 7288 18760
rect 7243 18720 7288 18748
rect 7282 18708 7288 18720
rect 7340 18708 7346 18760
rect 9950 18708 9956 18760
rect 10008 18757 10014 18760
rect 10152 18757 10180 18788
rect 10008 18751 10057 18757
rect 10008 18717 10011 18751
rect 10045 18717 10057 18751
rect 10008 18711 10057 18717
rect 10134 18751 10192 18757
rect 10134 18717 10146 18751
rect 10180 18717 10192 18751
rect 10134 18711 10192 18717
rect 10229 18751 10287 18757
rect 10229 18717 10241 18751
rect 10275 18745 10287 18751
rect 10413 18751 10471 18757
rect 10275 18717 10364 18745
rect 10229 18711 10287 18717
rect 10008 18708 10014 18711
rect 5758 18652 6684 18680
rect 5758 18649 5770 18652
rect 5712 18643 5770 18649
rect 6914 18640 6920 18692
rect 6972 18680 6978 18692
rect 9125 18683 9183 18689
rect 9125 18680 9137 18683
rect 6972 18652 9137 18680
rect 6972 18640 6978 18652
rect 9125 18649 9137 18652
rect 9171 18649 9183 18683
rect 10336 18680 10364 18717
rect 10413 18717 10425 18751
rect 10459 18748 10471 18751
rect 10686 18748 10692 18760
rect 10459 18720 10692 18748
rect 10459 18717 10471 18720
rect 10413 18711 10471 18717
rect 10686 18708 10692 18720
rect 10744 18708 10750 18760
rect 10888 18692 10916 18788
rect 11164 18757 11192 18856
rect 12250 18844 12256 18856
rect 12308 18844 12314 18896
rect 12360 18856 14044 18884
rect 11606 18816 11612 18828
rect 11519 18788 11612 18816
rect 11532 18757 11560 18788
rect 11606 18776 11612 18788
rect 11664 18816 11670 18828
rect 12360 18816 12388 18856
rect 14016 18828 14044 18856
rect 14182 18844 14188 18896
rect 14240 18884 14246 18896
rect 15749 18887 15807 18893
rect 15749 18884 15761 18887
rect 14240 18856 15761 18884
rect 14240 18844 14246 18856
rect 15749 18853 15761 18856
rect 15795 18853 15807 18887
rect 15749 18847 15807 18853
rect 11664 18788 12388 18816
rect 12437 18819 12495 18825
rect 11664 18776 11670 18788
rect 12437 18785 12449 18819
rect 12483 18816 12495 18819
rect 13078 18816 13084 18828
rect 12483 18788 13084 18816
rect 12483 18785 12495 18788
rect 12437 18779 12495 18785
rect 13078 18776 13084 18788
rect 13136 18776 13142 18828
rect 13998 18776 14004 18828
rect 14056 18776 14062 18828
rect 14274 18776 14280 18828
rect 14332 18816 14338 18828
rect 14369 18819 14427 18825
rect 14369 18816 14381 18819
rect 14332 18788 14381 18816
rect 14332 18776 14338 18788
rect 14369 18785 14381 18788
rect 14415 18785 14427 18819
rect 14369 18779 14427 18785
rect 15657 18819 15715 18825
rect 15657 18785 15669 18819
rect 15703 18816 15715 18819
rect 16132 18816 16160 18924
rect 16482 18912 16488 18964
rect 16540 18952 16546 18964
rect 21910 18952 21916 18964
rect 16540 18924 20208 18952
rect 21871 18924 21916 18952
rect 16540 18912 16546 18924
rect 16206 18844 16212 18896
rect 16264 18884 16270 18896
rect 16264 18856 18092 18884
rect 16264 18844 16270 18856
rect 18064 18825 18092 18856
rect 18322 18844 18328 18896
rect 18380 18844 18386 18896
rect 18509 18887 18567 18893
rect 18509 18853 18521 18887
rect 18555 18884 18567 18887
rect 18874 18884 18880 18896
rect 18555 18856 18880 18884
rect 18555 18853 18567 18856
rect 18509 18847 18567 18853
rect 18874 18844 18880 18856
rect 18932 18844 18938 18896
rect 20180 18884 20208 18924
rect 21910 18912 21916 18924
rect 21968 18912 21974 18964
rect 26786 18952 26792 18964
rect 22066 18924 26792 18952
rect 22066 18884 22094 18924
rect 26786 18912 26792 18924
rect 26844 18912 26850 18964
rect 27246 18952 27252 18964
rect 27207 18924 27252 18952
rect 27246 18912 27252 18924
rect 27304 18912 27310 18964
rect 20180 18856 22094 18884
rect 18049 18819 18107 18825
rect 15703 18788 16084 18816
rect 16132 18788 16804 18816
rect 15703 18785 15715 18788
rect 15657 18779 15715 18785
rect 11149 18751 11207 18757
rect 11149 18717 11161 18751
rect 11195 18717 11207 18751
rect 11149 18711 11207 18717
rect 11238 18748 11296 18754
rect 11354 18751 11412 18757
rect 11238 18714 11250 18748
rect 11284 18714 11297 18748
rect 11238 18708 11297 18714
rect 11354 18717 11366 18751
rect 11400 18748 11412 18751
rect 11517 18751 11575 18757
rect 11400 18720 11468 18748
rect 11400 18717 11412 18720
rect 11354 18711 11412 18717
rect 10594 18680 10600 18692
rect 10336 18652 10600 18680
rect 9125 18643 9183 18649
rect 10594 18640 10600 18652
rect 10652 18640 10658 18692
rect 10870 18640 10876 18692
rect 10928 18680 10934 18692
rect 11269 18680 11297 18708
rect 10928 18652 11297 18680
rect 11440 18680 11468 18720
rect 11517 18717 11529 18751
rect 11563 18717 11575 18751
rect 11517 18711 11575 18717
rect 11977 18751 12035 18757
rect 11977 18717 11989 18751
rect 12023 18748 12035 18751
rect 12066 18748 12072 18760
rect 12023 18720 12072 18748
rect 12023 18717 12035 18720
rect 11977 18711 12035 18717
rect 12066 18708 12072 18720
rect 12124 18708 12130 18760
rect 12158 18708 12164 18760
rect 12216 18748 12222 18760
rect 12526 18748 12532 18760
rect 12216 18720 12261 18748
rect 12487 18720 12532 18748
rect 12216 18708 12222 18720
rect 12526 18708 12532 18720
rect 12584 18708 12590 18760
rect 13173 18751 13231 18757
rect 13173 18748 13185 18751
rect 12912 18720 13185 18748
rect 11606 18680 11612 18692
rect 11440 18652 11612 18680
rect 10928 18640 10934 18652
rect 11606 18640 11612 18652
rect 11664 18640 11670 18692
rect 4724 18584 5238 18612
rect 6086 18572 6092 18624
rect 6144 18612 6150 18624
rect 6362 18612 6368 18624
rect 6144 18584 6368 18612
rect 6144 18572 6150 18584
rect 6362 18572 6368 18584
rect 6420 18572 6426 18624
rect 9490 18572 9496 18624
rect 9548 18612 9554 18624
rect 12618 18612 12624 18624
rect 9548 18584 12624 18612
rect 9548 18572 9554 18584
rect 12618 18572 12624 18584
rect 12676 18612 12682 18624
rect 12912 18612 12940 18720
rect 13173 18717 13185 18720
rect 13219 18748 13231 18751
rect 13814 18748 13820 18760
rect 13219 18720 13820 18748
rect 13219 18717 13231 18720
rect 13173 18711 13231 18717
rect 13814 18708 13820 18720
rect 13872 18708 13878 18760
rect 14090 18748 14096 18760
rect 14051 18720 14096 18748
rect 14090 18708 14096 18720
rect 14148 18708 14154 18760
rect 15010 18708 15016 18760
rect 15068 18748 15074 18760
rect 15565 18751 15623 18757
rect 15565 18748 15577 18751
rect 15068 18720 15577 18748
rect 15068 18708 15074 18720
rect 15565 18717 15577 18720
rect 15611 18717 15623 18751
rect 15565 18711 15623 18717
rect 15841 18751 15899 18757
rect 15841 18717 15853 18751
rect 15887 18748 15899 18751
rect 15930 18748 15936 18760
rect 15887 18720 15936 18748
rect 15887 18717 15899 18720
rect 15841 18711 15899 18717
rect 15930 18708 15936 18720
rect 15988 18708 15994 18760
rect 12986 18640 12992 18692
rect 13044 18680 13050 18692
rect 13357 18683 13415 18689
rect 13357 18680 13369 18683
rect 13044 18652 13369 18680
rect 13044 18640 13050 18652
rect 13357 18649 13369 18652
rect 13403 18649 13415 18683
rect 13357 18643 13415 18649
rect 12676 18584 12940 18612
rect 12676 18572 12682 18584
rect 15194 18572 15200 18624
rect 15252 18612 15258 18624
rect 15381 18615 15439 18621
rect 15381 18612 15393 18615
rect 15252 18584 15393 18612
rect 15252 18572 15258 18584
rect 15381 18581 15393 18584
rect 15427 18581 15439 18615
rect 16056 18612 16084 18788
rect 16482 18748 16488 18760
rect 16443 18720 16488 18748
rect 16482 18708 16488 18720
rect 16540 18708 16546 18760
rect 16776 18757 16804 18788
rect 18049 18785 18061 18819
rect 18095 18785 18107 18819
rect 18049 18779 18107 18785
rect 18141 18819 18199 18825
rect 18141 18785 18153 18819
rect 18187 18816 18199 18819
rect 18340 18816 18368 18844
rect 18187 18788 18368 18816
rect 18187 18785 18199 18788
rect 18141 18779 18199 18785
rect 22094 18776 22100 18828
rect 22152 18816 22158 18828
rect 22465 18819 22523 18825
rect 22465 18816 22477 18819
rect 22152 18788 22477 18816
rect 22152 18776 22158 18788
rect 22465 18785 22477 18788
rect 22511 18785 22523 18819
rect 22465 18779 22523 18785
rect 23198 18776 23204 18828
rect 23256 18816 23262 18828
rect 23569 18819 23627 18825
rect 23569 18816 23581 18819
rect 23256 18788 23581 18816
rect 23256 18776 23262 18788
rect 23569 18785 23581 18788
rect 23615 18785 23627 18819
rect 23569 18779 23627 18785
rect 16761 18751 16819 18757
rect 16761 18717 16773 18751
rect 16807 18748 16819 18751
rect 17402 18748 17408 18760
rect 16807 18720 17408 18748
rect 16807 18717 16819 18720
rect 16761 18711 16819 18717
rect 17402 18708 17408 18720
rect 17460 18748 17466 18760
rect 17770 18748 17776 18760
rect 17460 18720 17776 18748
rect 17460 18708 17466 18720
rect 17770 18708 17776 18720
rect 17828 18708 17834 18760
rect 17862 18708 17868 18760
rect 17920 18748 17926 18760
rect 17957 18751 18015 18757
rect 17957 18748 17969 18751
rect 17920 18720 17969 18748
rect 17920 18708 17926 18720
rect 17957 18717 17969 18720
rect 18003 18717 18015 18751
rect 17957 18711 18015 18717
rect 18325 18751 18383 18757
rect 18325 18717 18337 18751
rect 18371 18748 18383 18751
rect 18414 18748 18420 18760
rect 18371 18720 18420 18748
rect 18371 18717 18383 18720
rect 18325 18711 18383 18717
rect 18414 18708 18420 18720
rect 18472 18708 18478 18760
rect 18782 18708 18788 18760
rect 18840 18748 18846 18760
rect 19245 18751 19303 18757
rect 19245 18748 19257 18751
rect 18840 18720 19257 18748
rect 18840 18708 18846 18720
rect 19245 18717 19257 18720
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 19501 18751 19559 18757
rect 19501 18717 19513 18751
rect 19547 18736 19559 18751
rect 21269 18751 21327 18757
rect 21269 18748 21281 18751
rect 19812 18744 19932 18748
rect 20272 18744 21281 18748
rect 19501 18711 19515 18717
rect 19509 18684 19515 18711
rect 19567 18684 19573 18736
rect 19812 18720 21281 18744
rect 17034 18612 17040 18624
rect 16056 18584 17040 18612
rect 15381 18575 15439 18581
rect 17034 18572 17040 18584
rect 17092 18572 17098 18624
rect 17218 18572 17224 18624
rect 17276 18612 17282 18624
rect 19812 18612 19840 18720
rect 19904 18716 20300 18720
rect 21269 18717 21281 18720
rect 21315 18717 21327 18751
rect 21269 18711 21327 18717
rect 22002 18708 22008 18760
rect 22060 18748 22066 18760
rect 23293 18751 23351 18757
rect 23293 18748 23305 18751
rect 22060 18720 23305 18748
rect 22060 18708 22066 18720
rect 23293 18717 23305 18720
rect 23339 18717 23351 18751
rect 23293 18711 23351 18717
rect 23477 18751 23535 18757
rect 23477 18717 23489 18751
rect 23523 18748 23535 18751
rect 24302 18748 24308 18760
rect 23523 18720 24308 18748
rect 23523 18717 23535 18720
rect 23477 18711 23535 18717
rect 24302 18708 24308 18720
rect 24360 18708 24366 18760
rect 24765 18751 24823 18757
rect 24765 18717 24777 18751
rect 24811 18748 24823 18751
rect 24854 18748 24860 18760
rect 24811 18720 24860 18748
rect 24811 18717 24823 18720
rect 24765 18711 24823 18717
rect 24854 18708 24860 18720
rect 24912 18708 24918 18760
rect 27065 18751 27123 18757
rect 27065 18748 27077 18751
rect 24964 18720 27077 18748
rect 20898 18640 20904 18692
rect 20956 18680 20962 18692
rect 24964 18680 24992 18720
rect 27065 18717 27077 18720
rect 27111 18717 27123 18751
rect 27065 18711 27123 18717
rect 20956 18652 24992 18680
rect 25032 18683 25090 18689
rect 20956 18640 20962 18652
rect 25032 18649 25044 18683
rect 25078 18680 25090 18683
rect 25130 18680 25136 18692
rect 25078 18652 25136 18680
rect 25078 18649 25090 18652
rect 25032 18643 25090 18649
rect 25130 18640 25136 18652
rect 25188 18640 25194 18692
rect 17276 18584 19840 18612
rect 17276 18572 17282 18584
rect 19886 18572 19892 18624
rect 19944 18612 19950 18624
rect 20625 18615 20683 18621
rect 20625 18612 20637 18615
rect 19944 18584 20637 18612
rect 19944 18572 19950 18584
rect 20625 18581 20637 18584
rect 20671 18581 20683 18615
rect 20625 18575 20683 18581
rect 21085 18615 21143 18621
rect 21085 18581 21097 18615
rect 21131 18612 21143 18615
rect 21358 18612 21364 18624
rect 21131 18584 21364 18612
rect 21131 18581 21143 18584
rect 21085 18575 21143 18581
rect 21358 18572 21364 18584
rect 21416 18572 21422 18624
rect 22278 18612 22284 18624
rect 22239 18584 22284 18612
rect 22278 18572 22284 18584
rect 22336 18572 22342 18624
rect 22370 18572 22376 18624
rect 22428 18612 22434 18624
rect 23106 18612 23112 18624
rect 22428 18584 22473 18612
rect 23067 18584 23112 18612
rect 22428 18572 22434 18584
rect 23106 18572 23112 18584
rect 23164 18572 23170 18624
rect 24946 18572 24952 18624
rect 25004 18612 25010 18624
rect 26145 18615 26203 18621
rect 26145 18612 26157 18615
rect 25004 18584 26157 18612
rect 25004 18572 25010 18584
rect 26145 18581 26157 18584
rect 26191 18581 26203 18615
rect 26145 18575 26203 18581
rect 1104 18522 28060 18544
rect 1104 18470 9935 18522
rect 9987 18470 9999 18522
rect 10051 18470 10063 18522
rect 10115 18470 10127 18522
rect 10179 18470 10191 18522
rect 10243 18470 18920 18522
rect 18972 18470 18984 18522
rect 19036 18470 19048 18522
rect 19100 18470 19112 18522
rect 19164 18470 19176 18522
rect 19228 18470 28060 18522
rect 1104 18448 28060 18470
rect 1946 18368 1952 18420
rect 2004 18408 2010 18420
rect 2222 18408 2228 18420
rect 2004 18380 2228 18408
rect 2004 18368 2010 18380
rect 2222 18368 2228 18380
rect 2280 18368 2286 18420
rect 5350 18368 5356 18420
rect 5408 18408 5414 18420
rect 5408 18380 6960 18408
rect 5408 18368 5414 18380
rect 3602 18340 3608 18352
rect 1964 18312 3608 18340
rect 1964 18216 1992 18312
rect 3602 18300 3608 18312
rect 3660 18300 3666 18352
rect 4893 18343 4951 18349
rect 4893 18309 4905 18343
rect 4939 18340 4951 18343
rect 4939 18312 5488 18340
rect 4939 18309 4951 18312
rect 4893 18303 4951 18309
rect 2216 18275 2274 18281
rect 2216 18241 2228 18275
rect 2262 18272 2274 18275
rect 2498 18272 2504 18284
rect 2262 18244 2504 18272
rect 2262 18241 2274 18244
rect 2216 18235 2274 18241
rect 2498 18232 2504 18244
rect 2556 18232 2562 18284
rect 4065 18275 4123 18281
rect 4065 18241 4077 18275
rect 4111 18241 4123 18275
rect 4065 18235 4123 18241
rect 1946 18204 1952 18216
rect 1907 18176 1952 18204
rect 1946 18164 1952 18176
rect 2004 18164 2010 18216
rect 4080 18204 4108 18235
rect 4154 18232 4160 18284
rect 4212 18272 4218 18284
rect 4525 18275 4583 18281
rect 4525 18272 4537 18275
rect 4212 18244 4537 18272
rect 4212 18232 4218 18244
rect 4525 18241 4537 18244
rect 4571 18241 4583 18275
rect 4525 18235 4583 18241
rect 4614 18232 4620 18284
rect 4672 18272 4678 18284
rect 4709 18275 4767 18281
rect 4709 18272 4721 18275
rect 4672 18244 4721 18272
rect 4672 18232 4678 18244
rect 4709 18241 4721 18244
rect 4755 18241 4767 18275
rect 5350 18272 5356 18284
rect 5311 18244 5356 18272
rect 4709 18235 4767 18241
rect 5350 18232 5356 18244
rect 5408 18232 5414 18284
rect 5460 18272 5488 18312
rect 5534 18300 5540 18352
rect 5592 18340 5598 18352
rect 5592 18312 5637 18340
rect 5592 18300 5598 18312
rect 5902 18300 5908 18352
rect 5960 18340 5966 18352
rect 6822 18340 6828 18352
rect 5960 18312 6828 18340
rect 5960 18300 5966 18312
rect 6822 18300 6828 18312
rect 6880 18300 6886 18352
rect 6932 18340 6960 18380
rect 7282 18368 7288 18420
rect 7340 18408 7346 18420
rect 7745 18411 7803 18417
rect 7745 18408 7757 18411
rect 7340 18380 7757 18408
rect 7340 18368 7346 18380
rect 7745 18377 7757 18380
rect 7791 18377 7803 18411
rect 7745 18371 7803 18377
rect 6932 18312 7420 18340
rect 5718 18272 5724 18284
rect 5460 18244 5724 18272
rect 5718 18232 5724 18244
rect 5776 18232 5782 18284
rect 6454 18232 6460 18284
rect 6512 18272 6518 18284
rect 6621 18275 6679 18281
rect 6621 18272 6633 18275
rect 6512 18244 6633 18272
rect 6512 18232 6518 18244
rect 6621 18241 6633 18244
rect 6667 18241 6679 18275
rect 6621 18235 6679 18241
rect 4890 18204 4896 18216
rect 4080 18176 4896 18204
rect 4890 18164 4896 18176
rect 4948 18164 4954 18216
rect 6362 18204 6368 18216
rect 6323 18176 6368 18204
rect 6362 18164 6368 18176
rect 6420 18164 6426 18216
rect 3329 18139 3387 18145
rect 3329 18105 3341 18139
rect 3375 18136 3387 18139
rect 5902 18136 5908 18148
rect 3375 18108 5908 18136
rect 3375 18105 3387 18108
rect 3329 18099 3387 18105
rect 5902 18096 5908 18108
rect 5960 18096 5966 18148
rect 7392 18136 7420 18312
rect 7760 18272 7788 18371
rect 7926 18368 7932 18420
rect 7984 18408 7990 18420
rect 8297 18411 8355 18417
rect 8297 18408 8309 18411
rect 7984 18380 8309 18408
rect 7984 18368 7990 18380
rect 8297 18377 8309 18380
rect 8343 18377 8355 18411
rect 8297 18371 8355 18377
rect 10318 18368 10324 18420
rect 10376 18368 10382 18420
rect 10870 18368 10876 18420
rect 10928 18408 10934 18420
rect 11977 18411 12035 18417
rect 11977 18408 11989 18411
rect 10928 18380 11989 18408
rect 10928 18368 10934 18380
rect 11977 18377 11989 18380
rect 12023 18377 12035 18411
rect 13262 18408 13268 18420
rect 11977 18371 12035 18377
rect 12176 18380 13268 18408
rect 10336 18340 10364 18368
rect 12066 18340 12072 18352
rect 12124 18349 12130 18352
rect 12124 18343 12137 18349
rect 10336 18312 12072 18340
rect 8205 18275 8263 18281
rect 8205 18272 8217 18275
rect 7760 18244 8217 18272
rect 8205 18241 8217 18244
rect 8251 18241 8263 18275
rect 9490 18272 9496 18284
rect 9451 18244 9496 18272
rect 8205 18235 8263 18241
rect 9490 18232 9496 18244
rect 9548 18232 9554 18284
rect 9582 18232 9588 18284
rect 9640 18272 9646 18284
rect 10134 18272 10140 18284
rect 9640 18244 10140 18272
rect 9640 18232 9646 18244
rect 10134 18232 10140 18244
rect 10192 18232 10198 18284
rect 10689 18275 10747 18281
rect 10689 18272 10701 18275
rect 10336 18244 10701 18272
rect 9214 18204 9220 18216
rect 9175 18176 9220 18204
rect 9214 18164 9220 18176
rect 9272 18164 9278 18216
rect 10042 18136 10048 18148
rect 7392 18108 10048 18136
rect 10042 18096 10048 18108
rect 10100 18096 10106 18148
rect 3878 18068 3884 18080
rect 3839 18040 3884 18068
rect 3878 18028 3884 18040
rect 3936 18028 3942 18080
rect 4246 18028 4252 18080
rect 4304 18068 4310 18080
rect 5721 18071 5779 18077
rect 5721 18068 5733 18071
rect 4304 18040 5733 18068
rect 4304 18028 4310 18040
rect 5721 18037 5733 18040
rect 5767 18037 5779 18071
rect 5721 18031 5779 18037
rect 8754 18028 8760 18080
rect 8812 18068 8818 18080
rect 10134 18068 10140 18080
rect 8812 18040 10140 18068
rect 8812 18028 8818 18040
rect 10134 18028 10140 18040
rect 10192 18028 10198 18080
rect 10336 18068 10364 18244
rect 10689 18241 10701 18244
rect 10735 18241 10747 18275
rect 10870 18272 10876 18284
rect 10831 18244 10876 18272
rect 10689 18235 10747 18241
rect 10870 18232 10876 18244
rect 10928 18232 10934 18284
rect 10980 18281 11008 18312
rect 12066 18300 12072 18312
rect 12125 18340 12137 18343
rect 12176 18340 12204 18380
rect 13262 18368 13268 18380
rect 13320 18368 13326 18420
rect 14737 18411 14795 18417
rect 14737 18377 14749 18411
rect 14783 18408 14795 18411
rect 14826 18408 14832 18420
rect 14783 18380 14832 18408
rect 14783 18377 14795 18380
rect 14737 18371 14795 18377
rect 14826 18368 14832 18380
rect 14884 18368 14890 18420
rect 15746 18368 15752 18420
rect 15804 18408 15810 18420
rect 16025 18411 16083 18417
rect 16025 18408 16037 18411
rect 15804 18380 16037 18408
rect 15804 18368 15810 18380
rect 16025 18377 16037 18380
rect 16071 18377 16083 18411
rect 16025 18371 16083 18377
rect 16482 18368 16488 18420
rect 16540 18408 16546 18420
rect 17402 18408 17408 18420
rect 16540 18380 17408 18408
rect 16540 18368 16546 18380
rect 17402 18368 17408 18380
rect 17460 18368 17466 18420
rect 18598 18408 18604 18420
rect 18529 18380 18604 18408
rect 13998 18340 14004 18352
rect 12125 18312 12204 18340
rect 12728 18312 14004 18340
rect 12125 18309 12137 18312
rect 12124 18303 12137 18309
rect 12124 18300 12130 18303
rect 10965 18275 11023 18281
rect 10965 18241 10977 18275
rect 11011 18241 11023 18275
rect 11790 18272 11796 18284
rect 11751 18244 11796 18272
rect 10965 18235 11023 18241
rect 11790 18232 11796 18244
rect 11848 18232 11854 18284
rect 12728 18281 12756 18312
rect 13998 18300 14004 18312
rect 14056 18340 14062 18352
rect 14056 18312 14320 18340
rect 14056 18300 14062 18312
rect 12713 18275 12771 18281
rect 12713 18241 12725 18275
rect 12759 18241 12771 18275
rect 12894 18272 12900 18284
rect 12855 18244 12900 18272
rect 12713 18235 12771 18241
rect 12894 18232 12900 18244
rect 12952 18232 12958 18284
rect 14090 18272 14096 18284
rect 14051 18244 14096 18272
rect 14090 18232 14096 18244
rect 14148 18232 14154 18284
rect 14292 18281 14320 18312
rect 14277 18275 14335 18281
rect 14277 18241 14289 18275
rect 14323 18272 14335 18275
rect 14921 18275 14979 18281
rect 14921 18272 14933 18275
rect 14323 18244 14933 18272
rect 14323 18241 14335 18244
rect 14277 18235 14335 18241
rect 14921 18241 14933 18244
rect 14967 18241 14979 18275
rect 15102 18272 15108 18284
rect 15063 18244 15108 18272
rect 14921 18235 14979 18241
rect 15102 18232 15108 18244
rect 15160 18232 15166 18284
rect 15194 18232 15200 18284
rect 15252 18272 15258 18284
rect 15657 18275 15715 18281
rect 15252 18244 15297 18272
rect 15252 18232 15258 18244
rect 15657 18241 15669 18275
rect 15703 18241 15715 18275
rect 15657 18235 15715 18241
rect 15841 18275 15899 18281
rect 15841 18241 15853 18275
rect 15887 18272 15899 18275
rect 15930 18272 15936 18284
rect 15887 18244 15936 18272
rect 15887 18241 15899 18244
rect 15841 18235 15899 18241
rect 11698 18164 11704 18216
rect 11756 18204 11762 18216
rect 12066 18204 12072 18216
rect 11756 18176 12072 18204
rect 11756 18164 11762 18176
rect 12066 18164 12072 18176
rect 12124 18164 12130 18216
rect 12989 18207 13047 18213
rect 12989 18204 13001 18207
rect 12406 18176 13001 18204
rect 10689 18139 10747 18145
rect 10689 18105 10701 18139
rect 10735 18136 10747 18139
rect 12406 18136 12434 18176
rect 12989 18173 13001 18176
rect 13035 18204 13047 18207
rect 13078 18204 13084 18216
rect 13035 18176 13084 18204
rect 13035 18173 13047 18176
rect 12989 18167 13047 18173
rect 13078 18164 13084 18176
rect 13136 18164 13142 18216
rect 13814 18164 13820 18216
rect 13872 18204 13878 18216
rect 15010 18204 15016 18216
rect 13872 18176 15016 18204
rect 13872 18164 13878 18176
rect 15010 18164 15016 18176
rect 15068 18204 15074 18216
rect 15672 18204 15700 18235
rect 15930 18232 15936 18244
rect 15988 18232 15994 18284
rect 17770 18232 17776 18284
rect 17828 18272 17834 18284
rect 17957 18275 18015 18281
rect 17957 18272 17969 18275
rect 17828 18244 17969 18272
rect 17828 18232 17834 18244
rect 17957 18241 17969 18244
rect 18003 18241 18015 18275
rect 17957 18235 18015 18241
rect 18141 18275 18199 18281
rect 18141 18241 18153 18275
rect 18187 18241 18199 18275
rect 18322 18272 18328 18284
rect 18283 18244 18328 18272
rect 18141 18235 18199 18241
rect 15068 18176 15700 18204
rect 15068 18164 15074 18176
rect 16482 18164 16488 18216
rect 16540 18204 16546 18216
rect 16669 18207 16727 18213
rect 16669 18204 16681 18207
rect 16540 18176 16681 18204
rect 16540 18164 16546 18176
rect 16669 18173 16681 18176
rect 16715 18173 16727 18207
rect 16669 18167 16727 18173
rect 16945 18207 17003 18213
rect 16945 18173 16957 18207
rect 16991 18204 17003 18207
rect 17862 18204 17868 18216
rect 16991 18176 17868 18204
rect 16991 18173 17003 18176
rect 16945 18167 17003 18173
rect 17862 18164 17868 18176
rect 17920 18204 17926 18216
rect 18156 18204 18184 18235
rect 18322 18232 18328 18244
rect 18380 18232 18386 18284
rect 18529 18281 18557 18380
rect 18598 18368 18604 18380
rect 18656 18368 18662 18420
rect 19429 18411 19487 18417
rect 18892 18380 19380 18408
rect 18892 18352 18920 18380
rect 18874 18300 18880 18352
rect 18932 18300 18938 18352
rect 19352 18340 19380 18380
rect 19429 18377 19441 18411
rect 19475 18408 19487 18411
rect 19518 18408 19524 18420
rect 19475 18380 19524 18408
rect 19475 18377 19487 18380
rect 19429 18371 19487 18377
rect 19518 18368 19524 18380
rect 19576 18368 19582 18420
rect 20530 18408 20536 18420
rect 20491 18380 20536 18408
rect 20530 18368 20536 18380
rect 20588 18368 20594 18420
rect 20898 18408 20904 18420
rect 20640 18380 20904 18408
rect 20640 18340 20668 18380
rect 20898 18368 20904 18380
rect 20956 18368 20962 18420
rect 20993 18411 21051 18417
rect 20993 18377 21005 18411
rect 21039 18408 21051 18411
rect 21821 18411 21879 18417
rect 21821 18408 21833 18411
rect 21039 18380 21833 18408
rect 21039 18377 21051 18380
rect 20993 18371 21051 18377
rect 21821 18377 21833 18380
rect 21867 18377 21879 18411
rect 21821 18371 21879 18377
rect 22094 18368 22100 18420
rect 22152 18408 22158 18420
rect 22189 18411 22247 18417
rect 22189 18408 22201 18411
rect 22152 18380 22201 18408
rect 22152 18368 22158 18380
rect 22189 18377 22201 18380
rect 22235 18408 22247 18411
rect 24670 18408 24676 18420
rect 22235 18380 24676 18408
rect 22235 18377 22247 18380
rect 22189 18371 22247 18377
rect 24670 18368 24676 18380
rect 24728 18368 24734 18420
rect 19352 18312 20668 18340
rect 20806 18300 20812 18352
rect 20864 18340 20870 18352
rect 23284 18343 23342 18349
rect 20864 18312 22232 18340
rect 20864 18300 20870 18312
rect 22204 18284 22232 18312
rect 23284 18309 23296 18343
rect 23330 18340 23342 18343
rect 23934 18340 23940 18352
rect 23330 18312 23940 18340
rect 23330 18309 23342 18312
rect 23284 18303 23342 18309
rect 23934 18300 23940 18312
rect 23992 18300 23998 18352
rect 25308 18343 25366 18349
rect 25308 18309 25320 18343
rect 25354 18340 25366 18343
rect 26510 18340 26516 18352
rect 25354 18312 26516 18340
rect 25354 18309 25366 18312
rect 25308 18303 25366 18309
rect 26510 18300 26516 18312
rect 26568 18300 26574 18352
rect 18520 18275 18578 18281
rect 18520 18241 18532 18275
rect 18566 18241 18578 18275
rect 18520 18235 18578 18241
rect 18966 18232 18972 18284
rect 19024 18272 19030 18284
rect 19426 18272 19432 18284
rect 19024 18244 19432 18272
rect 19024 18232 19030 18244
rect 19426 18232 19432 18244
rect 19484 18232 19490 18284
rect 19610 18272 19616 18284
rect 19571 18244 19616 18272
rect 19610 18232 19616 18244
rect 19668 18232 19674 18284
rect 19702 18232 19708 18284
rect 19760 18272 19766 18284
rect 19797 18275 19855 18281
rect 19797 18272 19809 18275
rect 19760 18244 19809 18272
rect 19760 18232 19766 18244
rect 19797 18241 19809 18244
rect 19843 18241 19855 18275
rect 20898 18272 20904 18284
rect 20859 18244 20904 18272
rect 19797 18235 19855 18241
rect 20898 18232 20904 18244
rect 20956 18232 20962 18284
rect 22186 18232 22192 18284
rect 22244 18272 22250 18284
rect 26970 18272 26976 18284
rect 22244 18244 22416 18272
rect 26883 18244 26976 18272
rect 22244 18232 22250 18244
rect 17920 18176 18184 18204
rect 18233 18207 18291 18213
rect 17920 18164 17926 18176
rect 18233 18173 18245 18207
rect 18279 18173 18291 18207
rect 18340 18204 18368 18232
rect 18874 18204 18880 18216
rect 18340 18176 18880 18204
rect 18233 18167 18291 18173
rect 10735 18108 12434 18136
rect 10735 18105 10747 18108
rect 10689 18099 10747 18105
rect 12618 18096 12624 18148
rect 12676 18136 12682 18148
rect 18248 18136 18276 18167
rect 18874 18164 18880 18176
rect 18932 18164 18938 18216
rect 19886 18204 19892 18216
rect 19847 18176 19892 18204
rect 19886 18164 19892 18176
rect 19944 18164 19950 18216
rect 19978 18164 19984 18216
rect 20036 18204 20042 18216
rect 21085 18207 21143 18213
rect 21085 18204 21097 18207
rect 20036 18176 21097 18204
rect 20036 18164 20042 18176
rect 21085 18173 21097 18176
rect 21131 18173 21143 18207
rect 21085 18167 21143 18173
rect 21818 18164 21824 18216
rect 21876 18204 21882 18216
rect 22388 18213 22416 18244
rect 26970 18232 26976 18244
rect 27028 18232 27034 18284
rect 27157 18275 27215 18281
rect 27157 18241 27169 18275
rect 27203 18272 27215 18275
rect 27338 18272 27344 18284
rect 27203 18244 27344 18272
rect 27203 18241 27215 18244
rect 27157 18235 27215 18241
rect 27338 18232 27344 18244
rect 27396 18232 27402 18284
rect 22281 18207 22339 18213
rect 22281 18204 22293 18207
rect 21876 18176 22293 18204
rect 21876 18164 21882 18176
rect 22281 18173 22293 18176
rect 22327 18173 22339 18207
rect 22281 18167 22339 18173
rect 22373 18207 22431 18213
rect 22373 18173 22385 18207
rect 22419 18173 22431 18207
rect 22373 18167 22431 18173
rect 23017 18207 23075 18213
rect 23017 18173 23029 18207
rect 23063 18173 23075 18207
rect 23017 18167 23075 18173
rect 12676 18108 18276 18136
rect 12676 18096 12682 18108
rect 20806 18096 20812 18148
rect 20864 18136 20870 18148
rect 21174 18136 21180 18148
rect 20864 18108 21180 18136
rect 20864 18096 20870 18108
rect 21174 18096 21180 18108
rect 21232 18096 21238 18148
rect 21910 18096 21916 18148
rect 21968 18136 21974 18148
rect 23032 18136 23060 18167
rect 24854 18164 24860 18216
rect 24912 18204 24918 18216
rect 25038 18204 25044 18216
rect 24912 18176 25044 18204
rect 24912 18164 24918 18176
rect 25038 18164 25044 18176
rect 25096 18164 25102 18216
rect 26988 18204 27016 18232
rect 27246 18204 27252 18216
rect 26988 18176 27252 18204
rect 27246 18164 27252 18176
rect 27304 18164 27310 18216
rect 21968 18108 23060 18136
rect 21968 18096 21974 18108
rect 11146 18068 11152 18080
rect 10336 18040 11152 18068
rect 11146 18028 11152 18040
rect 11204 18028 11210 18080
rect 11609 18071 11667 18077
rect 11609 18037 11621 18071
rect 11655 18068 11667 18071
rect 11790 18068 11796 18080
rect 11655 18040 11796 18068
rect 11655 18037 11667 18040
rect 11609 18031 11667 18037
rect 11790 18028 11796 18040
rect 11848 18028 11854 18080
rect 12526 18068 12532 18080
rect 12487 18040 12532 18068
rect 12526 18028 12532 18040
rect 12584 18028 12590 18080
rect 13262 18028 13268 18080
rect 13320 18068 13326 18080
rect 15194 18068 15200 18080
rect 13320 18040 15200 18068
rect 13320 18028 13326 18040
rect 15194 18028 15200 18040
rect 15252 18028 15258 18080
rect 17862 18028 17868 18080
rect 17920 18068 17926 18080
rect 18693 18071 18751 18077
rect 18693 18068 18705 18071
rect 17920 18040 18705 18068
rect 17920 18028 17926 18040
rect 18693 18037 18705 18040
rect 18739 18037 18751 18071
rect 18693 18031 18751 18037
rect 19978 18028 19984 18080
rect 20036 18068 20042 18080
rect 21082 18068 21088 18080
rect 20036 18040 21088 18068
rect 20036 18028 20042 18040
rect 21082 18028 21088 18040
rect 21140 18028 21146 18080
rect 23934 18028 23940 18080
rect 23992 18068 23998 18080
rect 24397 18071 24455 18077
rect 24397 18068 24409 18071
rect 23992 18040 24409 18068
rect 23992 18028 23998 18040
rect 24397 18037 24409 18040
rect 24443 18037 24455 18071
rect 24397 18031 24455 18037
rect 25314 18028 25320 18080
rect 25372 18068 25378 18080
rect 26421 18071 26479 18077
rect 26421 18068 26433 18071
rect 25372 18040 26433 18068
rect 25372 18028 25378 18040
rect 26421 18037 26433 18040
rect 26467 18037 26479 18071
rect 26421 18031 26479 18037
rect 26973 18071 27031 18077
rect 26973 18037 26985 18071
rect 27019 18068 27031 18071
rect 27154 18068 27160 18080
rect 27019 18040 27160 18068
rect 27019 18037 27031 18040
rect 26973 18031 27031 18037
rect 27154 18028 27160 18040
rect 27212 18028 27218 18080
rect 1104 17978 28060 18000
rect 1104 17926 5442 17978
rect 5494 17926 5506 17978
rect 5558 17926 5570 17978
rect 5622 17926 5634 17978
rect 5686 17926 5698 17978
rect 5750 17926 14428 17978
rect 14480 17926 14492 17978
rect 14544 17926 14556 17978
rect 14608 17926 14620 17978
rect 14672 17926 14684 17978
rect 14736 17926 23413 17978
rect 23465 17926 23477 17978
rect 23529 17926 23541 17978
rect 23593 17926 23605 17978
rect 23657 17926 23669 17978
rect 23721 17926 28060 17978
rect 1104 17904 28060 17926
rect 2590 17824 2596 17876
rect 2648 17864 2654 17876
rect 6454 17864 6460 17876
rect 2648 17836 5939 17864
rect 6415 17836 6460 17864
rect 2648 17824 2654 17836
rect 3602 17688 3608 17740
rect 3660 17728 3666 17740
rect 3789 17731 3847 17737
rect 3789 17728 3801 17731
rect 3660 17700 3801 17728
rect 3660 17688 3666 17700
rect 3789 17697 3801 17700
rect 3835 17697 3847 17731
rect 3789 17691 3847 17697
rect 4890 17688 4896 17740
rect 4948 17728 4954 17740
rect 5626 17728 5632 17740
rect 4948 17700 5632 17728
rect 4948 17688 4954 17700
rect 5626 17688 5632 17700
rect 5684 17688 5690 17740
rect 5911 17728 5939 17836
rect 6454 17824 6460 17836
rect 6512 17824 6518 17876
rect 8294 17864 8300 17876
rect 7116 17836 8300 17864
rect 5911 17700 6960 17728
rect 1857 17663 1915 17669
rect 1857 17629 1869 17663
rect 1903 17660 1915 17663
rect 1946 17660 1952 17672
rect 1903 17632 1952 17660
rect 1903 17629 1915 17632
rect 1857 17623 1915 17629
rect 1946 17620 1952 17632
rect 2004 17620 2010 17672
rect 3878 17620 3884 17672
rect 3936 17660 3942 17672
rect 4045 17663 4103 17669
rect 4045 17660 4057 17663
rect 3936 17632 4057 17660
rect 3936 17620 3942 17632
rect 4045 17629 4057 17632
rect 4091 17629 4103 17663
rect 4045 17623 4103 17629
rect 5813 17663 5871 17669
rect 5813 17629 5825 17663
rect 5859 17660 5871 17663
rect 5902 17660 5908 17672
rect 5859 17632 5908 17660
rect 5859 17629 5871 17632
rect 5813 17623 5871 17629
rect 5902 17620 5908 17632
rect 5960 17620 5966 17672
rect 6638 17620 6644 17672
rect 6696 17660 6702 17672
rect 6932 17669 6960 17700
rect 7116 17669 7144 17836
rect 8294 17824 8300 17836
rect 8352 17824 8358 17876
rect 9398 17824 9404 17876
rect 9456 17864 9462 17876
rect 11514 17864 11520 17876
rect 9456 17836 11520 17864
rect 9456 17824 9462 17836
rect 11514 17824 11520 17836
rect 11572 17824 11578 17876
rect 12989 17867 13047 17873
rect 12989 17833 13001 17867
rect 13035 17864 13047 17867
rect 13170 17864 13176 17876
rect 13035 17836 13176 17864
rect 13035 17833 13047 17836
rect 12989 17827 13047 17833
rect 13170 17824 13176 17836
rect 13228 17824 13234 17876
rect 13262 17824 13268 17876
rect 13320 17864 13326 17876
rect 13722 17864 13728 17876
rect 13320 17836 13728 17864
rect 13320 17824 13326 17836
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 14826 17824 14832 17876
rect 14884 17864 14890 17876
rect 14884 17836 15148 17864
rect 14884 17824 14890 17836
rect 15120 17808 15148 17836
rect 15654 17824 15660 17876
rect 15712 17864 15718 17876
rect 15930 17864 15936 17876
rect 15712 17836 15936 17864
rect 15712 17824 15718 17836
rect 15930 17824 15936 17836
rect 15988 17824 15994 17876
rect 16301 17867 16359 17873
rect 16301 17833 16313 17867
rect 16347 17864 16359 17867
rect 16390 17864 16396 17876
rect 16347 17836 16396 17864
rect 16347 17833 16359 17836
rect 16301 17827 16359 17833
rect 16390 17824 16396 17836
rect 16448 17824 16454 17876
rect 17218 17824 17224 17876
rect 17276 17864 17282 17876
rect 21818 17864 21824 17876
rect 17276 17836 21824 17864
rect 17276 17824 17282 17836
rect 21818 17824 21824 17836
rect 21876 17864 21882 17876
rect 23198 17864 23204 17876
rect 21876 17836 23204 17864
rect 21876 17824 21882 17836
rect 23198 17824 23204 17836
rect 23256 17864 23262 17876
rect 23385 17867 23443 17873
rect 23385 17864 23397 17867
rect 23256 17836 23397 17864
rect 23256 17824 23262 17836
rect 23385 17833 23397 17836
rect 23431 17833 23443 17867
rect 23385 17827 23443 17833
rect 24026 17824 24032 17876
rect 24084 17864 24090 17876
rect 24084 17836 26740 17864
rect 24084 17824 24090 17836
rect 15102 17756 15108 17808
rect 15160 17796 15166 17808
rect 15473 17799 15531 17805
rect 15473 17796 15485 17799
rect 15160 17768 15485 17796
rect 15160 17756 15166 17768
rect 15473 17765 15485 17768
rect 15519 17765 15531 17799
rect 15473 17759 15531 17765
rect 19058 17756 19064 17808
rect 19116 17796 19122 17808
rect 20070 17796 20076 17808
rect 19116 17768 20076 17796
rect 19116 17756 19122 17768
rect 20070 17756 20076 17768
rect 20128 17756 20134 17808
rect 20714 17756 20720 17808
rect 20772 17796 20778 17808
rect 20772 17768 21680 17796
rect 20772 17756 20778 17768
rect 7561 17731 7619 17737
rect 7561 17697 7573 17731
rect 7607 17728 7619 17731
rect 8294 17728 8300 17740
rect 7607 17700 8300 17728
rect 7607 17697 7619 17700
rect 7561 17691 7619 17697
rect 8294 17688 8300 17700
rect 8352 17688 8358 17740
rect 18874 17688 18880 17740
rect 18932 17728 18938 17740
rect 19705 17731 19763 17737
rect 19705 17728 19717 17731
rect 18932 17700 19717 17728
rect 18932 17688 18938 17700
rect 19705 17697 19717 17700
rect 19751 17728 19763 17731
rect 19978 17728 19984 17740
rect 19751 17700 19984 17728
rect 19751 17697 19763 17700
rect 19705 17691 19763 17697
rect 19978 17688 19984 17700
rect 20036 17688 20042 17740
rect 20993 17731 21051 17737
rect 20993 17697 21005 17731
rect 21039 17728 21051 17731
rect 21542 17728 21548 17740
rect 21039 17700 21548 17728
rect 21039 17697 21051 17700
rect 20993 17691 21051 17697
rect 21542 17688 21548 17700
rect 21600 17688 21606 17740
rect 6733 17663 6791 17669
rect 6733 17660 6745 17663
rect 6696 17632 6745 17660
rect 6696 17620 6702 17632
rect 6733 17629 6745 17632
rect 6779 17629 6791 17663
rect 6733 17623 6791 17629
rect 6825 17663 6883 17669
rect 6825 17629 6837 17663
rect 6871 17629 6883 17663
rect 6825 17623 6883 17629
rect 6917 17663 6975 17669
rect 6917 17629 6929 17663
rect 6963 17629 6975 17663
rect 6917 17623 6975 17629
rect 7101 17663 7159 17669
rect 7101 17629 7113 17663
rect 7147 17629 7159 17663
rect 7101 17623 7159 17629
rect 7837 17663 7895 17669
rect 7837 17629 7849 17663
rect 7883 17660 7895 17663
rect 8662 17660 8668 17672
rect 7883 17632 8668 17660
rect 7883 17629 7895 17632
rect 7837 17623 7895 17629
rect 2124 17595 2182 17601
rect 2124 17561 2136 17595
rect 2170 17592 2182 17595
rect 3602 17592 3608 17604
rect 2170 17564 3608 17592
rect 2170 17561 2182 17564
rect 2124 17555 2182 17561
rect 3602 17552 3608 17564
rect 3660 17552 3666 17604
rect 5350 17552 5356 17604
rect 5408 17592 5414 17604
rect 5629 17595 5687 17601
rect 5629 17592 5641 17595
rect 5408 17564 5641 17592
rect 5408 17552 5414 17564
rect 5629 17561 5641 17564
rect 5675 17561 5687 17595
rect 6840 17592 6868 17623
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 8938 17620 8944 17672
rect 8996 17660 9002 17672
rect 9493 17663 9551 17669
rect 9493 17660 9505 17663
rect 8996 17632 9505 17660
rect 8996 17620 9002 17632
rect 9493 17629 9505 17632
rect 9539 17660 9551 17663
rect 10778 17660 10784 17672
rect 9539 17632 10784 17660
rect 9539 17629 9551 17632
rect 9493 17623 9551 17629
rect 10778 17620 10784 17632
rect 10836 17660 10842 17672
rect 11609 17663 11667 17669
rect 11609 17660 11621 17663
rect 10836 17632 11621 17660
rect 10836 17620 10842 17632
rect 11609 17629 11621 17632
rect 11655 17660 11667 17663
rect 14093 17663 14151 17669
rect 14093 17660 14105 17663
rect 11655 17632 14105 17660
rect 11655 17629 11667 17632
rect 11609 17623 11667 17629
rect 14093 17629 14105 17632
rect 14139 17629 14151 17663
rect 14093 17623 14151 17629
rect 17313 17663 17371 17669
rect 17313 17629 17325 17663
rect 17359 17660 17371 17663
rect 17954 17660 17960 17672
rect 17359 17632 17960 17660
rect 17359 17629 17371 17632
rect 17313 17623 17371 17629
rect 17954 17620 17960 17632
rect 18012 17660 18018 17672
rect 18782 17660 18788 17672
rect 18012 17632 18788 17660
rect 18012 17620 18018 17632
rect 18782 17620 18788 17632
rect 18840 17620 18846 17672
rect 19429 17663 19487 17669
rect 19429 17629 19441 17663
rect 19475 17629 19487 17663
rect 20806 17660 20812 17672
rect 20732 17647 20812 17660
rect 19429 17623 19487 17629
rect 20717 17641 20812 17647
rect 8570 17592 8576 17604
rect 6840 17564 8576 17592
rect 5629 17555 5687 17561
rect 8570 17552 8576 17564
rect 8628 17552 8634 17604
rect 9582 17552 9588 17604
rect 9640 17592 9646 17604
rect 9738 17595 9796 17601
rect 9738 17592 9750 17595
rect 9640 17564 9750 17592
rect 9640 17552 9646 17564
rect 9738 17561 9750 17564
rect 9784 17561 9796 17595
rect 9738 17555 9796 17561
rect 11876 17595 11934 17601
rect 11876 17561 11888 17595
rect 11922 17592 11934 17595
rect 12526 17592 12532 17604
rect 11922 17564 12532 17592
rect 11922 17561 11934 17564
rect 11876 17555 11934 17561
rect 12526 17552 12532 17564
rect 12584 17552 12590 17604
rect 13722 17552 13728 17604
rect 13780 17592 13786 17604
rect 14338 17595 14396 17601
rect 14338 17592 14350 17595
rect 13780 17564 14350 17592
rect 13780 17552 13786 17564
rect 14338 17561 14350 17564
rect 14384 17561 14396 17595
rect 14338 17555 14396 17561
rect 15010 17552 15016 17604
rect 15068 17592 15074 17604
rect 15933 17595 15991 17601
rect 15933 17592 15945 17595
rect 15068 17564 15945 17592
rect 15068 17552 15074 17564
rect 15933 17561 15945 17564
rect 15979 17561 15991 17595
rect 15933 17555 15991 17561
rect 16117 17595 16175 17601
rect 16117 17561 16129 17595
rect 16163 17592 16175 17595
rect 16482 17592 16488 17604
rect 16163 17564 16488 17592
rect 16163 17561 16175 17564
rect 16117 17555 16175 17561
rect 16482 17552 16488 17564
rect 16540 17552 16546 17604
rect 17586 17601 17592 17604
rect 17580 17592 17592 17601
rect 17547 17564 17592 17592
rect 17580 17555 17592 17564
rect 17586 17552 17592 17555
rect 17644 17552 17650 17604
rect 19444 17592 19472 17623
rect 20717 17607 20729 17641
rect 20763 17632 20812 17641
rect 20763 17607 20775 17632
rect 20806 17620 20812 17632
rect 20864 17620 20870 17672
rect 20901 17663 20959 17669
rect 20901 17629 20913 17663
rect 20947 17629 20959 17663
rect 20901 17623 20959 17629
rect 20622 17592 20628 17604
rect 17696 17564 20628 17592
rect 3237 17527 3295 17533
rect 3237 17493 3249 17527
rect 3283 17524 3295 17527
rect 4890 17524 4896 17536
rect 3283 17496 4896 17524
rect 3283 17493 3295 17496
rect 3237 17487 3295 17493
rect 4890 17484 4896 17496
rect 4948 17484 4954 17536
rect 5169 17527 5227 17533
rect 5169 17493 5181 17527
rect 5215 17524 5227 17527
rect 5534 17524 5540 17536
rect 5215 17496 5540 17524
rect 5215 17493 5227 17496
rect 5169 17487 5227 17493
rect 5534 17484 5540 17496
rect 5592 17484 5598 17536
rect 5718 17484 5724 17536
rect 5776 17524 5782 17536
rect 5997 17527 6055 17533
rect 5997 17524 6009 17527
rect 5776 17496 6009 17524
rect 5776 17484 5782 17496
rect 5997 17493 6009 17496
rect 6043 17493 6055 17527
rect 5997 17487 6055 17493
rect 10502 17484 10508 17536
rect 10560 17524 10566 17536
rect 10870 17524 10876 17536
rect 10560 17496 10876 17524
rect 10560 17484 10566 17496
rect 10870 17484 10876 17496
rect 10928 17484 10934 17536
rect 11514 17484 11520 17536
rect 11572 17524 11578 17536
rect 11790 17524 11796 17536
rect 11572 17496 11796 17524
rect 11572 17484 11578 17496
rect 11790 17484 11796 17496
rect 11848 17524 11854 17536
rect 17696 17524 17724 17564
rect 20622 17552 20628 17564
rect 20680 17552 20686 17604
rect 20717 17601 20775 17607
rect 20916 17592 20944 17623
rect 21082 17620 21088 17672
rect 21140 17660 21146 17672
rect 21269 17663 21327 17669
rect 21140 17632 21185 17660
rect 21140 17620 21146 17632
rect 21269 17629 21281 17663
rect 21315 17660 21327 17663
rect 21652 17660 21680 17768
rect 26712 17737 26740 17836
rect 26697 17731 26755 17737
rect 26697 17697 26709 17731
rect 26743 17728 26755 17731
rect 26878 17728 26884 17740
rect 26743 17700 26884 17728
rect 26743 17697 26755 17700
rect 26697 17691 26755 17697
rect 26878 17688 26884 17700
rect 26936 17688 26942 17740
rect 21315 17632 21680 17660
rect 21315 17629 21327 17632
rect 21269 17623 21327 17629
rect 21910 17620 21916 17672
rect 21968 17660 21974 17672
rect 22005 17663 22063 17669
rect 22005 17660 22017 17663
rect 21968 17632 22017 17660
rect 21968 17620 21974 17632
rect 22005 17629 22017 17632
rect 22051 17660 22063 17663
rect 24397 17663 24455 17669
rect 24397 17660 24409 17663
rect 22051 17632 24409 17660
rect 22051 17629 22063 17632
rect 22005 17623 22063 17629
rect 24397 17629 24409 17632
rect 24443 17660 24455 17663
rect 25038 17660 25044 17672
rect 24443 17632 25044 17660
rect 24443 17629 24455 17632
rect 24397 17623 24455 17629
rect 25038 17620 25044 17632
rect 25096 17620 25102 17672
rect 25774 17620 25780 17672
rect 25832 17660 25838 17672
rect 26421 17663 26479 17669
rect 26421 17660 26433 17663
rect 25832 17632 26433 17660
rect 25832 17620 25838 17632
rect 26421 17629 26433 17632
rect 26467 17629 26479 17663
rect 26421 17623 26479 17629
rect 26510 17620 26516 17672
rect 26568 17660 26574 17672
rect 26605 17663 26663 17669
rect 26605 17660 26617 17663
rect 26568 17632 26617 17660
rect 26568 17620 26574 17632
rect 26605 17629 26617 17632
rect 26651 17629 26663 17663
rect 26605 17623 26663 17629
rect 27341 17663 27399 17669
rect 27341 17629 27353 17663
rect 27387 17629 27399 17663
rect 27341 17623 27399 17629
rect 22094 17592 22100 17604
rect 20916 17564 22100 17592
rect 22094 17552 22100 17564
rect 22152 17552 22158 17604
rect 22272 17595 22330 17601
rect 22272 17561 22284 17595
rect 22318 17592 22330 17595
rect 23106 17592 23112 17604
rect 22318 17564 23112 17592
rect 22318 17561 22330 17564
rect 22272 17555 22330 17561
rect 23106 17552 23112 17564
rect 23164 17552 23170 17604
rect 24210 17552 24216 17604
rect 24268 17592 24274 17604
rect 24642 17595 24700 17601
rect 24642 17592 24654 17595
rect 24268 17564 24654 17592
rect 24268 17552 24274 17564
rect 24642 17561 24654 17564
rect 24688 17561 24700 17595
rect 27356 17592 27384 17623
rect 24642 17555 24700 17561
rect 24780 17564 27384 17592
rect 11848 17496 17724 17524
rect 11848 17484 11854 17496
rect 17770 17484 17776 17536
rect 17828 17524 17834 17536
rect 18693 17527 18751 17533
rect 18693 17524 18705 17527
rect 17828 17496 18705 17524
rect 17828 17484 17834 17496
rect 18693 17493 18705 17496
rect 18739 17493 18751 17527
rect 18693 17487 18751 17493
rect 21082 17484 21088 17536
rect 21140 17524 21146 17536
rect 21453 17527 21511 17533
rect 21453 17524 21465 17527
rect 21140 17496 21465 17524
rect 21140 17484 21146 17496
rect 21453 17493 21465 17496
rect 21499 17493 21511 17527
rect 21453 17487 21511 17493
rect 23290 17484 23296 17536
rect 23348 17524 23354 17536
rect 24780 17524 24808 17564
rect 23348 17496 24808 17524
rect 23348 17484 23354 17496
rect 24854 17484 24860 17536
rect 24912 17524 24918 17536
rect 25777 17527 25835 17533
rect 25777 17524 25789 17527
rect 24912 17496 25789 17524
rect 24912 17484 24918 17496
rect 25777 17493 25789 17496
rect 25823 17493 25835 17527
rect 25777 17487 25835 17493
rect 26237 17527 26295 17533
rect 26237 17493 26249 17527
rect 26283 17524 26295 17527
rect 26326 17524 26332 17536
rect 26283 17496 26332 17524
rect 26283 17493 26295 17496
rect 26237 17487 26295 17493
rect 26326 17484 26332 17496
rect 26384 17484 26390 17536
rect 26786 17484 26792 17536
rect 26844 17524 26850 17536
rect 27157 17527 27215 17533
rect 27157 17524 27169 17527
rect 26844 17496 27169 17524
rect 26844 17484 26850 17496
rect 27157 17493 27169 17496
rect 27203 17493 27215 17527
rect 27157 17487 27215 17493
rect 1104 17434 28060 17456
rect 1104 17382 9935 17434
rect 9987 17382 9999 17434
rect 10051 17382 10063 17434
rect 10115 17382 10127 17434
rect 10179 17382 10191 17434
rect 10243 17382 18920 17434
rect 18972 17382 18984 17434
rect 19036 17382 19048 17434
rect 19100 17382 19112 17434
rect 19164 17382 19176 17434
rect 19228 17382 28060 17434
rect 1104 17360 28060 17382
rect 2498 17280 2504 17332
rect 2556 17320 2562 17332
rect 3881 17323 3939 17329
rect 3881 17320 3893 17323
rect 2556 17292 3893 17320
rect 2556 17280 2562 17292
rect 3881 17289 3893 17292
rect 3927 17289 3939 17323
rect 5718 17320 5724 17332
rect 3881 17283 3939 17289
rect 4448 17292 5724 17320
rect 2216 17255 2274 17261
rect 2216 17221 2228 17255
rect 2262 17252 2274 17255
rect 3418 17252 3424 17264
rect 2262 17224 3424 17252
rect 2262 17221 2274 17224
rect 2216 17215 2274 17221
rect 3418 17212 3424 17224
rect 3476 17212 3482 17264
rect 4065 17187 4123 17193
rect 4065 17153 4077 17187
rect 4111 17184 4123 17187
rect 4448 17184 4476 17292
rect 5718 17280 5724 17292
rect 5776 17280 5782 17332
rect 9582 17320 9588 17332
rect 9543 17292 9588 17320
rect 9582 17280 9588 17292
rect 9640 17280 9646 17332
rect 10873 17323 10931 17329
rect 10873 17289 10885 17323
rect 10919 17320 10931 17323
rect 12158 17320 12164 17332
rect 10919 17292 12164 17320
rect 10919 17289 10931 17292
rect 10873 17283 10931 17289
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 12989 17323 13047 17329
rect 12989 17289 13001 17323
rect 13035 17320 13047 17323
rect 13170 17320 13176 17332
rect 13035 17292 13176 17320
rect 13035 17289 13047 17292
rect 12989 17283 13047 17289
rect 13170 17280 13176 17292
rect 13228 17280 13234 17332
rect 13722 17320 13728 17332
rect 13683 17292 13728 17320
rect 13722 17280 13728 17292
rect 13780 17280 13786 17332
rect 16758 17320 16764 17332
rect 13832 17292 16764 17320
rect 4709 17255 4767 17261
rect 4709 17221 4721 17255
rect 4755 17252 4767 17255
rect 4890 17252 4896 17264
rect 4755 17224 4896 17252
rect 4755 17221 4767 17224
rect 4709 17215 4767 17221
rect 4890 17212 4896 17224
rect 4948 17212 4954 17264
rect 5534 17252 5540 17264
rect 5495 17224 5540 17252
rect 5534 17212 5540 17224
rect 5592 17212 5598 17264
rect 11330 17252 11336 17264
rect 9876 17224 11336 17252
rect 4111 17156 4476 17184
rect 4525 17187 4583 17193
rect 4111 17153 4123 17156
rect 4065 17147 4123 17153
rect 4525 17153 4537 17187
rect 4571 17184 4583 17187
rect 5350 17184 5356 17196
rect 4571 17156 5356 17184
rect 4571 17153 4583 17156
rect 4525 17147 4583 17153
rect 1946 17116 1952 17128
rect 1907 17088 1952 17116
rect 1946 17076 1952 17088
rect 2004 17076 2010 17128
rect 4154 17076 4160 17128
rect 4212 17116 4218 17128
rect 4540 17116 4568 17147
rect 5350 17144 5356 17156
rect 5408 17144 5414 17196
rect 5626 17144 5632 17196
rect 5684 17184 5690 17196
rect 5721 17187 5779 17193
rect 5721 17184 5733 17187
rect 5684 17156 5733 17184
rect 5684 17144 5690 17156
rect 5721 17153 5733 17156
rect 5767 17153 5779 17187
rect 5721 17147 5779 17153
rect 6270 17144 6276 17196
rect 6328 17184 6334 17196
rect 6621 17187 6679 17193
rect 6621 17184 6633 17187
rect 6328 17156 6633 17184
rect 6328 17144 6334 17156
rect 6621 17153 6633 17156
rect 6667 17153 6679 17187
rect 8294 17184 8300 17196
rect 8207 17156 8300 17184
rect 6621 17147 6679 17153
rect 8294 17144 8300 17156
rect 8352 17184 8358 17196
rect 9214 17184 9220 17196
rect 8352 17156 9220 17184
rect 8352 17144 8358 17156
rect 9214 17144 9220 17156
rect 9272 17144 9278 17196
rect 9876 17193 9904 17224
rect 11330 17212 11336 17224
rect 11388 17212 11394 17264
rect 11790 17212 11796 17264
rect 11848 17252 11854 17264
rect 13832 17252 13860 17292
rect 16758 17280 16764 17292
rect 16816 17280 16822 17332
rect 17586 17320 17592 17332
rect 17547 17292 17592 17320
rect 17586 17280 17592 17292
rect 17644 17280 17650 17332
rect 19518 17320 19524 17332
rect 17696 17292 19524 17320
rect 14826 17252 14832 17264
rect 11848 17224 13860 17252
rect 14005 17224 14832 17252
rect 11848 17212 11854 17224
rect 9861 17187 9919 17193
rect 9861 17153 9873 17187
rect 9907 17153 9919 17187
rect 9861 17147 9919 17153
rect 9953 17187 10011 17193
rect 9953 17153 9965 17187
rect 9999 17153 10011 17187
rect 9953 17147 10011 17153
rect 10045 17187 10103 17193
rect 10045 17153 10057 17187
rect 10091 17153 10103 17187
rect 10045 17147 10103 17153
rect 10229 17187 10287 17193
rect 10229 17153 10241 17187
rect 10275 17153 10287 17187
rect 10229 17147 10287 17153
rect 4212 17088 4568 17116
rect 4212 17076 4218 17088
rect 5810 17076 5816 17128
rect 5868 17116 5874 17128
rect 6362 17116 6368 17128
rect 5868 17088 6368 17116
rect 5868 17076 5874 17088
rect 6362 17076 6368 17088
rect 6420 17076 6426 17128
rect 8570 17116 8576 17128
rect 8483 17088 8576 17116
rect 8570 17076 8576 17088
rect 8628 17076 8634 17128
rect 3329 17051 3387 17057
rect 3329 17017 3341 17051
rect 3375 17048 3387 17051
rect 4614 17048 4620 17060
rect 3375 17020 4620 17048
rect 3375 17017 3387 17020
rect 3329 17011 3387 17017
rect 4614 17008 4620 17020
rect 4672 17008 4678 17060
rect 8588 17048 8616 17076
rect 9968 17048 9996 17147
rect 8588 17020 9996 17048
rect 4522 16940 4528 16992
rect 4580 16980 4586 16992
rect 4706 16980 4712 16992
rect 4580 16952 4712 16980
rect 4580 16940 4586 16952
rect 4706 16940 4712 16952
rect 4764 16940 4770 16992
rect 4893 16983 4951 16989
rect 4893 16949 4905 16983
rect 4939 16980 4951 16983
rect 4982 16980 4988 16992
rect 4939 16952 4988 16980
rect 4939 16949 4951 16952
rect 4893 16943 4951 16949
rect 4982 16940 4988 16952
rect 5040 16940 5046 16992
rect 7374 16940 7380 16992
rect 7432 16980 7438 16992
rect 7745 16983 7803 16989
rect 7745 16980 7757 16983
rect 7432 16952 7757 16980
rect 7432 16940 7438 16952
rect 7745 16949 7757 16952
rect 7791 16949 7803 16983
rect 7745 16943 7803 16949
rect 9674 16940 9680 16992
rect 9732 16980 9738 16992
rect 10060 16980 10088 17147
rect 10244 17116 10272 17147
rect 10502 17144 10508 17196
rect 10560 17184 10566 17196
rect 10781 17187 10839 17193
rect 10781 17184 10793 17187
rect 10560 17156 10793 17184
rect 10560 17144 10566 17156
rect 10781 17153 10793 17156
rect 10827 17153 10839 17187
rect 11698 17184 11704 17196
rect 11659 17156 11704 17184
rect 10781 17147 10839 17153
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 11977 17187 12035 17193
rect 11977 17153 11989 17187
rect 12023 17153 12035 17187
rect 12158 17184 12164 17196
rect 12119 17156 12164 17184
rect 11977 17147 12035 17153
rect 10962 17116 10968 17128
rect 10244 17088 10968 17116
rect 10962 17076 10968 17088
rect 11020 17076 11026 17128
rect 11992 17116 12020 17147
rect 12158 17144 12164 17156
rect 12216 17144 12222 17196
rect 12802 17184 12808 17196
rect 12763 17156 12808 17184
rect 12802 17144 12808 17156
rect 12860 17144 12866 17196
rect 13078 17144 13084 17196
rect 13136 17184 13142 17196
rect 13136 17156 13181 17184
rect 13136 17144 13142 17156
rect 13538 17144 13544 17196
rect 13596 17184 13602 17196
rect 13722 17184 13728 17196
rect 13596 17156 13728 17184
rect 13596 17144 13602 17156
rect 13722 17144 13728 17156
rect 13780 17144 13786 17196
rect 14005 17193 14033 17224
rect 14826 17212 14832 17224
rect 14884 17212 14890 17264
rect 14921 17255 14979 17261
rect 14921 17221 14933 17255
rect 14967 17252 14979 17255
rect 15010 17252 15016 17264
rect 14967 17224 15016 17252
rect 14967 17221 14979 17224
rect 14921 17215 14979 17221
rect 15010 17212 15016 17224
rect 15068 17212 15074 17264
rect 17696 17252 17724 17292
rect 19518 17280 19524 17292
rect 19576 17280 19582 17332
rect 20806 17280 20812 17332
rect 20864 17320 20870 17332
rect 24210 17320 24216 17332
rect 20864 17292 23336 17320
rect 24171 17292 24216 17320
rect 20864 17280 20870 17292
rect 18782 17252 18788 17264
rect 15856 17224 17724 17252
rect 18743 17224 18788 17252
rect 13981 17187 14039 17193
rect 13981 17153 13993 17187
rect 14027 17153 14039 17187
rect 13981 17147 14039 17153
rect 14093 17187 14151 17193
rect 14093 17153 14105 17187
rect 14139 17153 14151 17187
rect 14093 17147 14151 17153
rect 14185 17187 14243 17193
rect 14185 17153 14197 17187
rect 14231 17153 14243 17187
rect 14366 17184 14372 17196
rect 14327 17156 14372 17184
rect 14185 17147 14243 17153
rect 12621 17119 12679 17125
rect 12621 17116 12633 17119
rect 11992 17088 12633 17116
rect 12621 17085 12633 17088
rect 12667 17085 12679 17119
rect 12621 17079 12679 17085
rect 13262 17076 13268 17128
rect 13320 17116 13326 17128
rect 14108 17116 14136 17147
rect 13320 17088 14136 17116
rect 14200 17116 14228 17147
rect 14366 17144 14372 17156
rect 14424 17144 14430 17196
rect 15856 17193 15884 17224
rect 18782 17212 18788 17224
rect 18840 17212 18846 17264
rect 19702 17212 19708 17264
rect 19760 17252 19766 17264
rect 20162 17252 20168 17264
rect 19760 17224 20168 17252
rect 19760 17212 19766 17224
rect 20162 17212 20168 17224
rect 20220 17212 20226 17264
rect 22094 17252 22100 17264
rect 22007 17224 22100 17252
rect 15105 17187 15163 17193
rect 15105 17153 15117 17187
rect 15151 17184 15163 17187
rect 15841 17187 15899 17193
rect 15151 17156 15792 17184
rect 15151 17153 15163 17156
rect 15105 17147 15163 17153
rect 15289 17119 15347 17125
rect 15289 17116 15301 17119
rect 14200 17088 15301 17116
rect 13320 17076 13326 17088
rect 15289 17085 15301 17088
rect 15335 17085 15347 17119
rect 15764 17116 15792 17156
rect 15841 17153 15853 17187
rect 15887 17153 15899 17187
rect 15841 17147 15899 17153
rect 15930 17144 15936 17196
rect 15988 17184 15994 17196
rect 16853 17187 16911 17193
rect 16853 17184 16865 17187
rect 15988 17156 16865 17184
rect 15988 17144 15994 17156
rect 16853 17153 16865 17156
rect 16899 17153 16911 17187
rect 16853 17147 16911 17153
rect 17310 17144 17316 17196
rect 17368 17144 17374 17196
rect 17773 17187 17831 17193
rect 17773 17153 17785 17187
rect 17819 17184 17831 17187
rect 18506 17184 18512 17196
rect 17819 17156 18512 17184
rect 17819 17153 17831 17156
rect 17773 17147 17831 17153
rect 18506 17144 18512 17156
rect 18564 17144 18570 17196
rect 18601 17187 18659 17193
rect 18601 17153 18613 17187
rect 18647 17184 18659 17187
rect 18690 17184 18696 17196
rect 18647 17156 18696 17184
rect 18647 17153 18659 17156
rect 18601 17147 18659 17153
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 19613 17187 19671 17193
rect 19613 17184 19625 17187
rect 18800 17156 19625 17184
rect 16390 17116 16396 17128
rect 15764 17088 16396 17116
rect 15289 17079 15347 17085
rect 16390 17076 16396 17088
rect 16448 17076 16454 17128
rect 16669 17119 16727 17125
rect 16669 17085 16681 17119
rect 16715 17116 16727 17119
rect 17218 17116 17224 17128
rect 16715 17088 17224 17116
rect 16715 17085 16727 17088
rect 16669 17079 16727 17085
rect 17218 17076 17224 17088
rect 17276 17076 17282 17128
rect 17328 17116 17356 17144
rect 17678 17116 17684 17128
rect 17328 17088 17684 17116
rect 17678 17076 17684 17088
rect 17736 17076 17742 17128
rect 18049 17119 18107 17125
rect 18049 17085 18061 17119
rect 18095 17116 18107 17119
rect 18800 17116 18828 17156
rect 19613 17153 19625 17156
rect 19659 17153 19671 17187
rect 20530 17184 20536 17196
rect 19613 17147 19671 17153
rect 19904 17156 20536 17184
rect 18095 17088 18828 17116
rect 18095 17085 18107 17088
rect 18049 17079 18107 17085
rect 11793 17051 11851 17057
rect 11793 17017 11805 17051
rect 11839 17017 11851 17051
rect 11793 17011 11851 17017
rect 11885 17051 11943 17057
rect 11885 17017 11897 17051
rect 11931 17048 11943 17051
rect 12158 17048 12164 17060
rect 11931 17020 12164 17048
rect 11931 17017 11943 17020
rect 11885 17011 11943 17017
rect 9732 16952 10088 16980
rect 9732 16940 9738 16952
rect 10962 16940 10968 16992
rect 11020 16980 11026 16992
rect 11517 16983 11575 16989
rect 11517 16980 11529 16983
rect 11020 16952 11529 16980
rect 11020 16940 11026 16952
rect 11517 16949 11529 16952
rect 11563 16949 11575 16983
rect 11808 16980 11836 17011
rect 12158 17008 12164 17020
rect 12216 17008 12222 17060
rect 16482 17008 16488 17060
rect 16540 17048 16546 17060
rect 17037 17051 17095 17057
rect 17037 17048 17049 17051
rect 16540 17020 17049 17048
rect 16540 17008 16546 17020
rect 17037 17017 17049 17020
rect 17083 17017 17095 17051
rect 17037 17011 17095 17017
rect 17770 17008 17776 17060
rect 17828 17048 17834 17060
rect 18064 17048 18092 17079
rect 19334 17076 19340 17128
rect 19392 17116 19398 17128
rect 19904 17125 19932 17156
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 21174 17144 21180 17196
rect 21232 17184 21238 17196
rect 22020 17193 22048 17224
rect 22094 17212 22100 17224
rect 22152 17252 22158 17264
rect 22152 17224 23244 17252
rect 22152 17212 22158 17224
rect 23216 17196 23244 17224
rect 21825 17187 21883 17193
rect 21825 17186 21837 17187
rect 21744 17184 21837 17186
rect 21232 17158 21837 17184
rect 21232 17156 21772 17158
rect 21232 17144 21238 17156
rect 21825 17153 21837 17158
rect 21871 17153 21883 17187
rect 21825 17147 21883 17153
rect 22005 17187 22063 17193
rect 22005 17153 22017 17187
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 22189 17187 22247 17193
rect 22189 17153 22201 17187
rect 22235 17184 22247 17187
rect 22373 17187 22431 17193
rect 22235 17156 22327 17184
rect 22235 17153 22247 17156
rect 22189 17147 22247 17153
rect 19705 17119 19763 17125
rect 19705 17116 19717 17119
rect 19392 17088 19717 17116
rect 19392 17076 19398 17088
rect 19705 17085 19717 17088
rect 19751 17085 19763 17119
rect 19705 17079 19763 17085
rect 19889 17119 19947 17125
rect 19889 17085 19901 17119
rect 19935 17085 19947 17119
rect 19889 17079 19947 17085
rect 20070 17076 20076 17128
rect 20128 17116 20134 17128
rect 20441 17119 20499 17125
rect 20441 17116 20453 17119
rect 20128 17088 20453 17116
rect 20128 17076 20134 17088
rect 20441 17085 20453 17088
rect 20487 17116 20499 17119
rect 21082 17116 21088 17128
rect 20487 17088 21088 17116
rect 20487 17085 20499 17088
rect 20441 17079 20499 17085
rect 21082 17076 21088 17088
rect 21140 17076 21146 17128
rect 22020 17116 22048 17147
rect 21928 17088 22048 17116
rect 17828 17020 18092 17048
rect 17828 17008 17834 17020
rect 18966 17008 18972 17060
rect 19024 17048 19030 17060
rect 20806 17048 20812 17060
rect 19024 17020 20812 17048
rect 19024 17008 19030 17020
rect 20806 17008 20812 17020
rect 20864 17008 20870 17060
rect 12526 16980 12532 16992
rect 11808 16952 12532 16980
rect 11517 16943 11575 16949
rect 12526 16940 12532 16952
rect 12584 16940 12590 16992
rect 16117 16983 16175 16989
rect 16117 16949 16129 16983
rect 16163 16980 16175 16983
rect 16850 16980 16856 16992
rect 16163 16952 16856 16980
rect 16163 16949 16175 16952
rect 16117 16943 16175 16949
rect 16850 16940 16856 16952
rect 16908 16940 16914 16992
rect 17310 16940 17316 16992
rect 17368 16980 17374 16992
rect 17957 16983 18015 16989
rect 17957 16980 17969 16983
rect 17368 16952 17969 16980
rect 17368 16940 17374 16952
rect 17957 16949 17969 16952
rect 18003 16949 18015 16983
rect 17957 16943 18015 16949
rect 18046 16940 18052 16992
rect 18104 16980 18110 16992
rect 19245 16983 19303 16989
rect 19245 16980 19257 16983
rect 18104 16952 19257 16980
rect 18104 16940 18110 16952
rect 19245 16949 19257 16952
rect 19291 16949 19303 16983
rect 19245 16943 19303 16949
rect 20671 16983 20729 16989
rect 20671 16949 20683 16983
rect 20717 16980 20729 16983
rect 21928 16980 21956 17088
rect 22094 17076 22100 17128
rect 22152 17116 22158 17128
rect 22299 17116 22327 17156
rect 22373 17153 22385 17187
rect 22419 17184 22431 17187
rect 22646 17184 22652 17196
rect 22419 17156 22652 17184
rect 22419 17153 22431 17156
rect 22373 17147 22431 17153
rect 22646 17144 22652 17156
rect 22704 17144 22710 17196
rect 23014 17184 23020 17196
rect 22975 17156 23020 17184
rect 23014 17144 23020 17156
rect 23072 17144 23078 17196
rect 23198 17184 23204 17196
rect 23159 17156 23204 17184
rect 23198 17144 23204 17156
rect 23256 17144 23262 17196
rect 23308 17193 23336 17292
rect 24210 17280 24216 17292
rect 24268 17280 24274 17332
rect 26234 17280 26240 17332
rect 26292 17320 26298 17332
rect 26292 17292 26372 17320
rect 26292 17280 26298 17292
rect 25685 17255 25743 17261
rect 25685 17221 25697 17255
rect 25731 17252 25743 17255
rect 26344 17252 26372 17292
rect 26694 17280 26700 17332
rect 26752 17320 26758 17332
rect 26970 17320 26976 17332
rect 26752 17292 26976 17320
rect 26752 17280 26758 17292
rect 26970 17280 26976 17292
rect 27028 17280 27034 17332
rect 27065 17255 27123 17261
rect 27065 17252 27077 17255
rect 25731 17224 26271 17252
rect 26344 17224 27077 17252
rect 25731 17221 25743 17224
rect 25685 17215 25743 17221
rect 23293 17187 23351 17193
rect 23293 17153 23305 17187
rect 23339 17153 23351 17187
rect 23293 17147 23351 17153
rect 23569 17187 23627 17193
rect 23569 17153 23581 17187
rect 23615 17184 23627 17187
rect 23658 17184 23664 17196
rect 23615 17156 23664 17184
rect 23615 17153 23627 17156
rect 23569 17147 23627 17153
rect 23658 17144 23664 17156
rect 23716 17144 23722 17196
rect 23753 17187 23811 17193
rect 23753 17153 23765 17187
rect 23799 17184 23811 17187
rect 24397 17187 24455 17193
rect 24397 17184 24409 17187
rect 23799 17156 24409 17184
rect 23799 17153 23811 17156
rect 23753 17147 23811 17153
rect 24397 17153 24409 17156
rect 24443 17153 24455 17187
rect 24670 17184 24676 17196
rect 24631 17156 24676 17184
rect 24397 17147 24455 17153
rect 24670 17144 24676 17156
rect 24728 17184 24734 17196
rect 24854 17184 24860 17196
rect 24728 17156 24860 17184
rect 24728 17144 24734 17156
rect 24854 17144 24860 17156
rect 24912 17144 24918 17196
rect 25130 17144 25136 17196
rect 25188 17184 25194 17196
rect 25869 17187 25927 17193
rect 25869 17184 25881 17187
rect 25188 17156 25881 17184
rect 25188 17144 25194 17156
rect 25869 17153 25881 17156
rect 25915 17153 25927 17187
rect 25869 17147 25927 17153
rect 25958 17144 25964 17196
rect 26016 17184 26022 17196
rect 26016 17156 26188 17184
rect 26016 17144 26022 17156
rect 23385 17119 23443 17125
rect 23385 17116 23397 17119
rect 22152 17088 22197 17116
rect 22299 17088 23397 17116
rect 22152 17076 22158 17088
rect 23385 17085 23397 17088
rect 23431 17116 23443 17119
rect 24026 17116 24032 17128
rect 23431 17088 24032 17116
rect 23431 17085 23443 17088
rect 23385 17079 23443 17085
rect 24026 17076 24032 17088
rect 24084 17076 24090 17128
rect 24302 17076 24308 17128
rect 24360 17116 24366 17128
rect 26160 17125 26188 17156
rect 26243 17128 26271 17224
rect 27065 17221 27077 17224
rect 27111 17221 27123 17255
rect 27065 17215 27123 17221
rect 24581 17119 24639 17125
rect 24581 17116 24593 17119
rect 24360 17088 24593 17116
rect 24360 17076 24366 17088
rect 24581 17085 24593 17088
rect 24627 17116 24639 17119
rect 26053 17119 26111 17125
rect 26053 17116 26065 17119
rect 24627 17088 26065 17116
rect 24627 17085 24639 17088
rect 24581 17079 24639 17085
rect 20717 16952 21956 16980
rect 22557 16983 22615 16989
rect 20717 16949 20729 16952
rect 20671 16943 20729 16949
rect 22557 16949 22569 16983
rect 22603 16980 22615 16983
rect 23290 16980 23296 16992
rect 22603 16952 23296 16980
rect 22603 16949 22615 16952
rect 22557 16943 22615 16949
rect 23290 16940 23296 16952
rect 23348 16940 23354 16992
rect 25884 16980 25912 17088
rect 26053 17085 26065 17088
rect 26099 17085 26111 17119
rect 26053 17079 26111 17085
rect 26145 17119 26203 17125
rect 26145 17085 26157 17119
rect 26191 17085 26203 17119
rect 26145 17079 26203 17085
rect 26234 17076 26240 17128
rect 26292 17076 26298 17128
rect 25958 17008 25964 17060
rect 26016 17048 26022 17060
rect 27249 17051 27307 17057
rect 27249 17048 27261 17051
rect 26016 17020 27261 17048
rect 26016 17008 26022 17020
rect 27249 17017 27261 17020
rect 27295 17017 27307 17051
rect 27249 17011 27307 17017
rect 26510 16980 26516 16992
rect 25884 16952 26516 16980
rect 26510 16940 26516 16952
rect 26568 16940 26574 16992
rect 1104 16890 28060 16912
rect 1104 16838 5442 16890
rect 5494 16838 5506 16890
rect 5558 16838 5570 16890
rect 5622 16838 5634 16890
rect 5686 16838 5698 16890
rect 5750 16838 14428 16890
rect 14480 16838 14492 16890
rect 14544 16838 14556 16890
rect 14608 16838 14620 16890
rect 14672 16838 14684 16890
rect 14736 16838 23413 16890
rect 23465 16838 23477 16890
rect 23529 16838 23541 16890
rect 23593 16838 23605 16890
rect 23657 16838 23669 16890
rect 23721 16838 28060 16890
rect 1104 16816 28060 16838
rect 3602 16736 3608 16788
rect 3660 16776 3666 16788
rect 4801 16779 4859 16785
rect 4801 16776 4813 16779
rect 3660 16748 4813 16776
rect 3660 16736 3666 16748
rect 4801 16745 4813 16748
rect 4847 16745 4859 16779
rect 6270 16776 6276 16788
rect 6231 16748 6276 16776
rect 4801 16739 4859 16745
rect 6270 16736 6276 16748
rect 6328 16736 6334 16788
rect 10137 16779 10195 16785
rect 10137 16745 10149 16779
rect 10183 16776 10195 16779
rect 11606 16776 11612 16788
rect 10183 16748 11612 16776
rect 10183 16745 10195 16748
rect 10137 16739 10195 16745
rect 11606 16736 11612 16748
rect 11664 16736 11670 16788
rect 11977 16779 12035 16785
rect 11977 16745 11989 16779
rect 12023 16776 12035 16779
rect 12802 16776 12808 16788
rect 12023 16748 12808 16776
rect 12023 16745 12035 16748
rect 11977 16739 12035 16745
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 15930 16736 15936 16788
rect 15988 16776 15994 16788
rect 15988 16748 16528 16776
rect 15988 16736 15994 16748
rect 1026 16668 1032 16720
rect 1084 16708 1090 16720
rect 1394 16708 1400 16720
rect 1084 16680 1400 16708
rect 1084 16668 1090 16680
rect 1394 16668 1400 16680
rect 1452 16668 1458 16720
rect 13449 16711 13507 16717
rect 11624 16680 12940 16708
rect 2866 16600 2872 16652
rect 2924 16640 2930 16652
rect 3602 16640 3608 16652
rect 2924 16612 3608 16640
rect 2924 16600 2930 16612
rect 3602 16600 3608 16612
rect 3660 16600 3666 16652
rect 5810 16600 5816 16652
rect 5868 16640 5874 16652
rect 7009 16643 7067 16649
rect 7009 16640 7021 16643
rect 5868 16612 7021 16640
rect 5868 16600 5874 16612
rect 7009 16609 7021 16612
rect 7055 16609 7067 16643
rect 7009 16603 7067 16609
rect 8938 16600 8944 16652
rect 8996 16640 9002 16652
rect 10597 16643 10655 16649
rect 10597 16640 10609 16643
rect 8996 16612 10609 16640
rect 8996 16600 9002 16612
rect 10597 16609 10609 16612
rect 10643 16609 10655 16643
rect 10597 16603 10655 16609
rect 1394 16532 1400 16584
rect 1452 16572 1458 16584
rect 1857 16575 1915 16581
rect 1857 16572 1869 16575
rect 1452 16544 1869 16572
rect 1452 16532 1458 16544
rect 1857 16541 1869 16544
rect 1903 16572 1915 16575
rect 1946 16572 1952 16584
rect 1903 16544 1952 16572
rect 1903 16541 1915 16544
rect 1857 16535 1915 16541
rect 1946 16532 1952 16544
rect 2004 16532 2010 16584
rect 4246 16532 4252 16584
rect 4304 16572 4310 16584
rect 4341 16575 4399 16581
rect 4341 16572 4353 16575
rect 4304 16544 4353 16572
rect 4304 16532 4310 16544
rect 4341 16541 4353 16544
rect 4387 16541 4399 16575
rect 4982 16572 4988 16584
rect 4943 16544 4988 16572
rect 4341 16535 4399 16541
rect 4982 16532 4988 16544
rect 5040 16532 5046 16584
rect 5166 16532 5172 16584
rect 5224 16572 5230 16584
rect 5629 16575 5687 16581
rect 5629 16572 5641 16575
rect 5224 16544 5641 16572
rect 5224 16532 5230 16544
rect 5629 16541 5641 16544
rect 5675 16541 5687 16575
rect 5629 16535 5687 16541
rect 6457 16575 6515 16581
rect 6457 16541 6469 16575
rect 6503 16572 6515 16575
rect 7558 16572 7564 16584
rect 6503 16544 7564 16572
rect 6503 16541 6515 16544
rect 6457 16535 6515 16541
rect 7558 16532 7564 16544
rect 7616 16532 7622 16584
rect 8386 16532 8392 16584
rect 8444 16572 8450 16584
rect 9125 16575 9183 16581
rect 9125 16572 9137 16575
rect 8444 16544 9137 16572
rect 8444 16532 8450 16544
rect 9125 16541 9137 16544
rect 9171 16541 9183 16575
rect 9125 16535 9183 16541
rect 9674 16532 9680 16584
rect 9732 16572 9738 16584
rect 11624 16572 11652 16680
rect 9732 16544 11652 16572
rect 12621 16575 12679 16581
rect 9732 16532 9738 16544
rect 12621 16541 12633 16575
rect 12667 16572 12679 16575
rect 12912 16572 12940 16680
rect 13449 16677 13461 16711
rect 13495 16708 13507 16711
rect 13538 16708 13544 16720
rect 13495 16680 13544 16708
rect 13495 16677 13507 16680
rect 13449 16671 13507 16677
rect 13538 16668 13544 16680
rect 13596 16668 13602 16720
rect 13998 16668 14004 16720
rect 14056 16708 14062 16720
rect 14737 16711 14795 16717
rect 14737 16708 14749 16711
rect 14056 16680 14749 16708
rect 14056 16668 14062 16680
rect 14737 16677 14749 16680
rect 14783 16677 14795 16711
rect 14737 16671 14795 16677
rect 15841 16711 15899 16717
rect 15841 16677 15853 16711
rect 15887 16708 15899 16711
rect 16206 16708 16212 16720
rect 15887 16680 16212 16708
rect 15887 16677 15899 16680
rect 15841 16671 15899 16677
rect 16206 16668 16212 16680
rect 16264 16668 16270 16720
rect 15930 16640 15936 16652
rect 13464 16612 15936 16640
rect 12667 16544 12940 16572
rect 13081 16575 13139 16581
rect 12667 16541 12679 16544
rect 12621 16535 12679 16541
rect 13081 16541 13093 16575
rect 13127 16572 13139 16575
rect 13354 16572 13360 16584
rect 13127 16544 13360 16572
rect 13127 16541 13139 16544
rect 13081 16535 13139 16541
rect 13354 16532 13360 16544
rect 13412 16532 13418 16584
rect 2124 16507 2182 16513
rect 2124 16473 2136 16507
rect 2170 16504 2182 16507
rect 7276 16507 7334 16513
rect 2170 16476 4200 16504
rect 2170 16473 2182 16476
rect 2124 16467 2182 16473
rect 3237 16439 3295 16445
rect 3237 16405 3249 16439
rect 3283 16436 3295 16439
rect 4062 16436 4068 16448
rect 3283 16408 4068 16436
rect 3283 16405 3295 16408
rect 3237 16399 3295 16405
rect 4062 16396 4068 16408
rect 4120 16396 4126 16448
rect 4172 16445 4200 16476
rect 7276 16473 7288 16507
rect 7322 16504 7334 16507
rect 7322 16476 8984 16504
rect 7322 16473 7334 16476
rect 7276 16467 7334 16473
rect 4157 16439 4215 16445
rect 4157 16405 4169 16439
rect 4203 16405 4215 16439
rect 5442 16436 5448 16448
rect 5403 16408 5448 16436
rect 4157 16399 4215 16405
rect 5442 16396 5448 16408
rect 5500 16396 5506 16448
rect 6270 16396 6276 16448
rect 6328 16436 6334 16448
rect 6730 16436 6736 16448
rect 6328 16408 6736 16436
rect 6328 16396 6334 16408
rect 6730 16396 6736 16408
rect 6788 16396 6794 16448
rect 8202 16396 8208 16448
rect 8260 16436 8266 16448
rect 8956 16445 8984 16476
rect 9582 16464 9588 16516
rect 9640 16504 9646 16516
rect 9769 16507 9827 16513
rect 9769 16504 9781 16507
rect 9640 16476 9781 16504
rect 9640 16464 9646 16476
rect 9769 16473 9781 16476
rect 9815 16473 9827 16507
rect 9769 16467 9827 16473
rect 9953 16507 10011 16513
rect 9953 16473 9965 16507
rect 9999 16504 10011 16507
rect 10686 16504 10692 16516
rect 9999 16476 10692 16504
rect 9999 16473 10011 16476
rect 9953 16467 10011 16473
rect 10686 16464 10692 16476
rect 10744 16464 10750 16516
rect 10864 16507 10922 16513
rect 10864 16473 10876 16507
rect 10910 16504 10922 16507
rect 10962 16504 10968 16516
rect 10910 16476 10968 16504
rect 10910 16473 10922 16476
rect 10864 16467 10922 16473
rect 10962 16464 10968 16476
rect 11020 16464 11026 16516
rect 12158 16464 12164 16516
rect 12216 16504 12222 16516
rect 13464 16504 13492 16612
rect 14573 16581 14601 16612
rect 15930 16600 15936 16612
rect 15988 16600 15994 16652
rect 16301 16643 16359 16649
rect 16301 16609 16313 16643
rect 16347 16609 16359 16643
rect 16301 16603 16359 16609
rect 14093 16575 14151 16581
rect 14093 16572 14105 16575
rect 12216 16476 13492 16504
rect 13556 16544 14105 16572
rect 12216 16464 12222 16476
rect 8389 16439 8447 16445
rect 8389 16436 8401 16439
rect 8260 16408 8401 16436
rect 8260 16396 8266 16408
rect 8389 16405 8401 16408
rect 8435 16405 8447 16439
rect 8389 16399 8447 16405
rect 8941 16439 8999 16445
rect 8941 16405 8953 16439
rect 8987 16405 8999 16439
rect 8941 16399 8999 16405
rect 12434 16396 12440 16448
rect 12492 16436 12498 16448
rect 13556 16445 13584 16544
rect 14093 16541 14105 16544
rect 14139 16541 14151 16575
rect 14093 16535 14151 16541
rect 14186 16575 14244 16581
rect 14186 16541 14198 16575
rect 14232 16541 14244 16575
rect 14186 16535 14244 16541
rect 14558 16575 14616 16581
rect 14558 16541 14570 16575
rect 14604 16541 14616 16575
rect 14558 16535 14616 16541
rect 13722 16464 13728 16516
rect 13780 16504 13786 16516
rect 14201 16504 14229 16535
rect 14826 16532 14832 16584
rect 14884 16572 14890 16584
rect 15378 16581 15384 16584
rect 15197 16575 15255 16581
rect 15197 16572 15209 16575
rect 14884 16544 15209 16572
rect 14884 16532 14890 16544
rect 15197 16541 15209 16544
rect 15243 16541 15255 16575
rect 15197 16535 15255 16541
rect 15345 16575 15384 16581
rect 15345 16541 15357 16575
rect 15345 16535 15384 16541
rect 15378 16532 15384 16535
rect 15436 16532 15442 16584
rect 15654 16572 15660 16584
rect 15712 16581 15718 16584
rect 15620 16544 15660 16572
rect 15654 16532 15660 16544
rect 15712 16535 15720 16581
rect 15712 16532 15718 16535
rect 14366 16504 14372 16516
rect 13780 16476 14229 16504
rect 14327 16476 14372 16504
rect 13780 16464 13786 16476
rect 14366 16464 14372 16476
rect 14424 16464 14430 16516
rect 14461 16507 14519 16513
rect 14461 16473 14473 16507
rect 14507 16473 14519 16507
rect 14461 16467 14519 16473
rect 13541 16439 13599 16445
rect 12492 16408 12537 16436
rect 12492 16396 12498 16408
rect 13541 16405 13553 16439
rect 13587 16405 13599 16439
rect 14476 16436 14504 16467
rect 15010 16464 15016 16516
rect 15068 16504 15074 16516
rect 15473 16507 15531 16513
rect 15473 16504 15485 16507
rect 15068 16476 15485 16504
rect 15068 16464 15074 16476
rect 15473 16473 15485 16476
rect 15519 16473 15531 16507
rect 15473 16467 15531 16473
rect 15565 16507 15623 16513
rect 15565 16473 15577 16507
rect 15611 16504 15623 16507
rect 15746 16504 15752 16516
rect 15611 16476 15752 16504
rect 15611 16473 15623 16476
rect 15565 16467 15623 16473
rect 15746 16464 15752 16476
rect 15804 16464 15810 16516
rect 15930 16464 15936 16516
rect 15988 16504 15994 16516
rect 16316 16504 16344 16603
rect 16500 16581 16528 16748
rect 17310 16736 17316 16788
rect 17368 16776 17374 16788
rect 18233 16779 18291 16785
rect 18233 16776 18245 16779
rect 17368 16748 18245 16776
rect 17368 16736 17374 16748
rect 18233 16745 18245 16748
rect 18279 16776 18291 16779
rect 19610 16776 19616 16788
rect 18279 16748 19616 16776
rect 18279 16745 18291 16748
rect 18233 16739 18291 16745
rect 19610 16736 19616 16748
rect 19668 16776 19674 16788
rect 19797 16779 19855 16785
rect 19797 16776 19809 16779
rect 19668 16748 19809 16776
rect 19668 16736 19674 16748
rect 19797 16745 19809 16748
rect 19843 16745 19855 16779
rect 19797 16739 19855 16745
rect 21913 16779 21971 16785
rect 21913 16745 21925 16779
rect 21959 16776 21971 16779
rect 22002 16776 22008 16788
rect 21959 16748 22008 16776
rect 21959 16745 21971 16748
rect 21913 16739 21971 16745
rect 22002 16736 22008 16748
rect 22060 16736 22066 16788
rect 25130 16776 25136 16788
rect 25091 16748 25136 16776
rect 25130 16736 25136 16748
rect 25188 16736 25194 16788
rect 17218 16708 17224 16720
rect 16960 16680 17224 16708
rect 16669 16643 16727 16649
rect 16669 16609 16681 16643
rect 16715 16640 16727 16643
rect 16960 16640 16988 16680
rect 17218 16668 17224 16680
rect 17276 16668 17282 16720
rect 17865 16711 17923 16717
rect 17865 16677 17877 16711
rect 17911 16708 17923 16711
rect 18046 16708 18052 16720
rect 17911 16680 18052 16708
rect 17911 16677 17923 16680
rect 17865 16671 17923 16677
rect 18046 16668 18052 16680
rect 18104 16668 18110 16720
rect 18506 16668 18512 16720
rect 18564 16708 18570 16720
rect 18564 16680 19472 16708
rect 18564 16668 18570 16680
rect 17405 16643 17463 16649
rect 17405 16640 17417 16643
rect 16715 16612 16988 16640
rect 17043 16612 17417 16640
rect 16715 16609 16727 16612
rect 16669 16603 16727 16609
rect 16485 16575 16543 16581
rect 16485 16541 16497 16575
rect 16531 16541 16543 16575
rect 16485 16535 16543 16541
rect 16942 16532 16948 16584
rect 17000 16572 17006 16584
rect 17043 16572 17071 16612
rect 17405 16609 17417 16612
rect 17451 16609 17463 16643
rect 17405 16603 17463 16609
rect 18325 16643 18383 16649
rect 18325 16609 18337 16643
rect 18371 16640 18383 16643
rect 19334 16640 19340 16652
rect 18371 16612 19340 16640
rect 18371 16609 18383 16612
rect 18325 16603 18383 16609
rect 18524 16584 18552 16612
rect 19334 16600 19340 16612
rect 19392 16600 19398 16652
rect 19444 16640 19472 16680
rect 20806 16668 20812 16720
rect 20864 16708 20870 16720
rect 21818 16708 21824 16720
rect 20864 16680 21824 16708
rect 20864 16668 20870 16680
rect 21818 16668 21824 16680
rect 21876 16668 21882 16720
rect 22094 16668 22100 16720
rect 22152 16708 22158 16720
rect 22646 16708 22652 16720
rect 22152 16680 22652 16708
rect 22152 16668 22158 16680
rect 22646 16668 22652 16680
rect 22704 16668 22710 16720
rect 24026 16708 24032 16720
rect 22756 16680 24032 16708
rect 21453 16643 21511 16649
rect 21453 16640 21465 16643
rect 19444 16612 21465 16640
rect 21453 16609 21465 16612
rect 21499 16609 21511 16643
rect 21453 16603 21511 16609
rect 21545 16643 21603 16649
rect 21545 16609 21557 16643
rect 21591 16640 21603 16643
rect 22756 16640 22784 16680
rect 24026 16668 24032 16680
rect 24084 16668 24090 16720
rect 21591 16612 22784 16640
rect 22833 16643 22891 16649
rect 21591 16609 21603 16612
rect 21545 16603 21603 16609
rect 22833 16609 22845 16643
rect 22879 16640 22891 16643
rect 22922 16640 22928 16652
rect 22879 16612 22928 16640
rect 22879 16609 22891 16612
rect 22833 16603 22891 16609
rect 22922 16600 22928 16612
rect 22980 16600 22986 16652
rect 23014 16600 23020 16652
rect 23072 16640 23078 16652
rect 23109 16643 23167 16649
rect 23109 16640 23121 16643
rect 23072 16612 23121 16640
rect 23072 16600 23078 16612
rect 23109 16609 23121 16612
rect 23155 16609 23167 16643
rect 23109 16603 23167 16609
rect 24210 16600 24216 16652
rect 24268 16640 24274 16652
rect 24673 16643 24731 16649
rect 24673 16640 24685 16643
rect 24268 16612 24685 16640
rect 24268 16600 24274 16612
rect 24673 16609 24685 16612
rect 24719 16609 24731 16643
rect 24673 16603 24731 16609
rect 25038 16600 25044 16652
rect 25096 16640 25102 16652
rect 25958 16640 25964 16652
rect 25096 16612 25964 16640
rect 25096 16600 25102 16612
rect 25958 16600 25964 16612
rect 26016 16600 26022 16652
rect 17770 16572 17776 16584
rect 17000 16544 17071 16572
rect 17144 16544 17776 16572
rect 17000 16532 17006 16544
rect 15988 16476 16344 16504
rect 15988 16464 15994 16476
rect 17144 16436 17172 16544
rect 17770 16532 17776 16544
rect 17828 16532 17834 16584
rect 18049 16575 18107 16581
rect 18049 16541 18061 16575
rect 18095 16572 18107 16575
rect 18138 16572 18144 16584
rect 18095 16544 18144 16572
rect 18095 16541 18107 16544
rect 18049 16535 18107 16541
rect 18138 16532 18144 16544
rect 18196 16532 18202 16584
rect 18506 16532 18512 16584
rect 18564 16532 18570 16584
rect 19426 16532 19432 16584
rect 19484 16572 19490 16584
rect 20533 16575 20591 16581
rect 20533 16572 20545 16575
rect 19484 16544 20545 16572
rect 19484 16532 19490 16544
rect 20533 16541 20545 16544
rect 20579 16541 20591 16575
rect 21174 16572 21180 16584
rect 21135 16544 21180 16572
rect 20533 16535 20591 16541
rect 21174 16532 21180 16544
rect 21232 16532 21238 16584
rect 21361 16575 21419 16581
rect 21361 16541 21373 16575
rect 21407 16541 21419 16575
rect 21361 16535 21419 16541
rect 21729 16575 21787 16581
rect 21729 16541 21741 16575
rect 21775 16572 21787 16575
rect 22002 16572 22008 16584
rect 21775 16544 22008 16572
rect 21775 16541 21787 16544
rect 21729 16535 21787 16541
rect 17221 16507 17279 16513
rect 17221 16473 17233 16507
rect 17267 16473 17279 16507
rect 17221 16467 17279 16473
rect 14476 16408 17172 16436
rect 17236 16436 17264 16467
rect 18782 16464 18788 16516
rect 18840 16504 18846 16516
rect 19705 16507 19763 16513
rect 19705 16504 19717 16507
rect 18840 16476 19717 16504
rect 18840 16464 18846 16476
rect 19705 16473 19717 16476
rect 19751 16473 19763 16507
rect 21376 16504 21404 16535
rect 22002 16532 22008 16544
rect 22060 16532 22066 16584
rect 24394 16572 24400 16584
rect 24355 16544 24400 16572
rect 24394 16532 24400 16544
rect 24452 16532 24458 16584
rect 26234 16581 26240 16584
rect 24581 16575 24639 16581
rect 24581 16541 24593 16575
rect 24627 16541 24639 16575
rect 24581 16535 24639 16541
rect 24765 16575 24823 16581
rect 24765 16541 24777 16575
rect 24811 16541 24823 16575
rect 24765 16535 24823 16541
rect 24949 16575 25007 16581
rect 24949 16541 24961 16575
rect 24995 16541 25007 16575
rect 26228 16572 26240 16581
rect 26195 16544 26240 16572
rect 24949 16535 25007 16541
rect 26228 16535 26240 16544
rect 23198 16504 23204 16516
rect 21376 16476 23204 16504
rect 19705 16467 19763 16473
rect 23198 16464 23204 16476
rect 23256 16504 23262 16516
rect 24596 16504 24624 16535
rect 23256 16476 24624 16504
rect 23256 16464 23262 16476
rect 24670 16464 24676 16516
rect 24728 16504 24734 16516
rect 24780 16504 24808 16535
rect 24728 16476 24808 16504
rect 24728 16464 24734 16476
rect 17402 16436 17408 16448
rect 17236 16408 17408 16436
rect 13541 16399 13599 16405
rect 17402 16396 17408 16408
rect 17460 16436 17466 16448
rect 17770 16436 17776 16448
rect 17460 16408 17776 16436
rect 17460 16396 17466 16408
rect 17770 16396 17776 16408
rect 17828 16396 17834 16448
rect 17862 16396 17868 16448
rect 17920 16436 17926 16448
rect 18138 16436 18144 16448
rect 17920 16408 18144 16436
rect 17920 16396 17926 16408
rect 18138 16396 18144 16408
rect 18196 16396 18202 16448
rect 20162 16396 20168 16448
rect 20220 16436 20226 16448
rect 20349 16439 20407 16445
rect 20349 16436 20361 16439
rect 20220 16408 20361 16436
rect 20220 16396 20226 16408
rect 20349 16405 20361 16408
rect 20395 16405 20407 16439
rect 20349 16399 20407 16405
rect 21082 16396 21088 16448
rect 21140 16436 21146 16448
rect 22002 16436 22008 16448
rect 21140 16408 22008 16436
rect 21140 16396 21146 16408
rect 22002 16396 22008 16408
rect 22060 16396 22066 16448
rect 24118 16396 24124 16448
rect 24176 16436 24182 16448
rect 24964 16436 24992 16535
rect 26234 16532 26240 16535
rect 26292 16532 26298 16584
rect 24176 16408 24992 16436
rect 24176 16396 24182 16408
rect 25222 16396 25228 16448
rect 25280 16436 25286 16448
rect 25866 16436 25872 16448
rect 25280 16408 25872 16436
rect 25280 16396 25286 16408
rect 25866 16396 25872 16408
rect 25924 16436 25930 16448
rect 27341 16439 27399 16445
rect 27341 16436 27353 16439
rect 25924 16408 27353 16436
rect 25924 16396 25930 16408
rect 27341 16405 27353 16408
rect 27387 16405 27399 16439
rect 27341 16399 27399 16405
rect 1104 16346 28060 16368
rect 1104 16294 9935 16346
rect 9987 16294 9999 16346
rect 10051 16294 10063 16346
rect 10115 16294 10127 16346
rect 10179 16294 10191 16346
rect 10243 16294 18920 16346
rect 18972 16294 18984 16346
rect 19036 16294 19048 16346
rect 19100 16294 19112 16346
rect 19164 16294 19176 16346
rect 19228 16294 28060 16346
rect 1104 16272 28060 16294
rect 4982 16192 4988 16244
rect 5040 16232 5046 16244
rect 5445 16235 5503 16241
rect 5445 16232 5457 16235
rect 5040 16204 5457 16232
rect 5040 16192 5046 16204
rect 5445 16201 5457 16204
rect 5491 16201 5503 16235
rect 7558 16232 7564 16244
rect 7519 16204 7564 16232
rect 5445 16195 5503 16201
rect 7558 16192 7564 16204
rect 7616 16192 7622 16244
rect 8386 16232 8392 16244
rect 7852 16204 8156 16232
rect 8347 16204 8392 16232
rect 1946 16124 1952 16176
rect 2004 16164 2010 16176
rect 5810 16164 5816 16176
rect 2004 16136 5816 16164
rect 2004 16124 2010 16136
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16065 2099 16099
rect 2498 16096 2504 16108
rect 2459 16068 2504 16096
rect 2041 16059 2099 16065
rect 2056 15960 2084 16059
rect 2498 16056 2504 16068
rect 2556 16056 2562 16108
rect 2685 16099 2743 16105
rect 2685 16065 2697 16099
rect 2731 16096 2743 16099
rect 2774 16096 2780 16108
rect 2731 16068 2780 16096
rect 2731 16065 2743 16068
rect 2685 16059 2743 16065
rect 2774 16056 2780 16068
rect 2832 16056 2838 16108
rect 3510 16096 3516 16108
rect 3471 16068 3516 16096
rect 3510 16056 3516 16068
rect 3568 16056 3574 16108
rect 4080 16105 4108 16136
rect 5810 16124 5816 16136
rect 5868 16124 5874 16176
rect 7193 16167 7251 16173
rect 7193 16133 7205 16167
rect 7239 16133 7251 16167
rect 7193 16127 7251 16133
rect 7409 16167 7467 16173
rect 7409 16133 7421 16167
rect 7455 16164 7467 16167
rect 7852 16164 7880 16204
rect 7455 16136 7880 16164
rect 7455 16133 7467 16136
rect 7409 16127 7467 16133
rect 4065 16099 4123 16105
rect 4065 16065 4077 16099
rect 4111 16065 4123 16099
rect 4065 16059 4123 16065
rect 4332 16099 4390 16105
rect 4332 16065 4344 16099
rect 4378 16096 4390 16099
rect 5442 16096 5448 16108
rect 4378 16068 5448 16096
rect 4378 16065 4390 16068
rect 4332 16059 4390 16065
rect 5442 16056 5448 16068
rect 5500 16056 5506 16108
rect 6549 16099 6607 16105
rect 6549 16065 6561 16099
rect 6595 16096 6607 16099
rect 6730 16096 6736 16108
rect 6595 16068 6736 16096
rect 6595 16065 6607 16068
rect 6549 16059 6607 16065
rect 6730 16056 6736 16068
rect 6788 16056 6794 16108
rect 7208 16096 7236 16127
rect 7926 16124 7932 16176
rect 7984 16164 7990 16176
rect 8021 16167 8079 16173
rect 8021 16164 8033 16167
rect 7984 16136 8033 16164
rect 7984 16124 7990 16136
rect 8021 16133 8033 16136
rect 8067 16133 8079 16167
rect 8128 16164 8156 16204
rect 8386 16192 8392 16204
rect 8444 16192 8450 16244
rect 12250 16192 12256 16244
rect 12308 16232 12314 16244
rect 12308 16204 13676 16232
rect 12308 16192 12314 16204
rect 8237 16167 8295 16173
rect 8237 16164 8249 16167
rect 8128 16136 8249 16164
rect 8021 16127 8079 16133
rect 8237 16133 8249 16136
rect 8283 16164 8295 16167
rect 8662 16164 8668 16176
rect 8283 16136 8668 16164
rect 8283 16133 8295 16136
rect 8237 16127 8295 16133
rect 8662 16124 8668 16136
rect 8720 16124 8726 16176
rect 9208 16167 9266 16173
rect 9208 16133 9220 16167
rect 9254 16164 9266 16167
rect 9398 16164 9404 16176
rect 9254 16136 9404 16164
rect 9254 16133 9266 16136
rect 9208 16127 9266 16133
rect 9398 16124 9404 16136
rect 9456 16124 9462 16176
rect 13648 16173 13676 16204
rect 13722 16192 13728 16244
rect 13780 16232 13786 16244
rect 14366 16232 14372 16244
rect 13780 16204 14372 16232
rect 13780 16192 13786 16204
rect 14366 16192 14372 16204
rect 14424 16192 14430 16244
rect 21818 16232 21824 16244
rect 15120 16204 21824 16232
rect 13633 16167 13691 16173
rect 13633 16133 13645 16167
rect 13679 16133 13691 16167
rect 13633 16127 13691 16133
rect 7944 16096 7972 16124
rect 8938 16096 8944 16108
rect 7208 16068 7972 16096
rect 8899 16068 8944 16096
rect 8938 16056 8944 16068
rect 8996 16056 9002 16108
rect 10778 16096 10784 16108
rect 10739 16068 10784 16096
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 10965 16099 11023 16105
rect 10965 16065 10977 16099
rect 11011 16096 11023 16099
rect 11606 16096 11612 16108
rect 11011 16068 11612 16096
rect 11011 16065 11023 16068
rect 10965 16059 11023 16065
rect 11606 16056 11612 16068
rect 11664 16056 11670 16108
rect 12158 16096 12164 16108
rect 12119 16068 12164 16096
rect 12158 16056 12164 16068
rect 12216 16056 12222 16108
rect 13078 16056 13084 16108
rect 13136 16096 13142 16108
rect 13265 16099 13323 16105
rect 13265 16096 13277 16099
rect 13136 16068 13277 16096
rect 13136 16056 13142 16068
rect 13265 16065 13277 16068
rect 13311 16065 13323 16099
rect 13265 16059 13323 16065
rect 13358 16099 13416 16105
rect 13358 16065 13370 16099
rect 13404 16065 13416 16099
rect 13538 16096 13544 16108
rect 13499 16068 13544 16096
rect 13358 16059 13416 16065
rect 10796 16028 10824 16056
rect 11885 16031 11943 16037
rect 11885 16028 11897 16031
rect 10796 16000 11897 16028
rect 11885 15997 11897 16000
rect 11931 15997 11943 16031
rect 11885 15991 11943 15997
rect 13170 15988 13176 16040
rect 13228 16028 13234 16040
rect 13372 16028 13400 16059
rect 13538 16056 13544 16068
rect 13596 16056 13602 16108
rect 13814 16105 13820 16108
rect 13771 16099 13820 16105
rect 13771 16065 13783 16099
rect 13817 16065 13820 16099
rect 13771 16059 13820 16065
rect 13814 16056 13820 16059
rect 13872 16056 13878 16108
rect 14366 16096 14372 16108
rect 14327 16068 14372 16096
rect 14366 16056 14372 16068
rect 14424 16056 14430 16108
rect 13228 16000 13400 16028
rect 13556 16028 13584 16056
rect 15010 16028 15016 16040
rect 13556 16000 15016 16028
rect 13228 15988 13234 16000
rect 15010 15988 15016 16000
rect 15068 15988 15074 16040
rect 2056 15932 4108 15960
rect 1857 15895 1915 15901
rect 1857 15861 1869 15895
rect 1903 15892 1915 15895
rect 2406 15892 2412 15904
rect 1903 15864 2412 15892
rect 1903 15861 1915 15864
rect 1857 15855 1915 15861
rect 2406 15852 2412 15864
rect 2464 15852 2470 15904
rect 2866 15892 2872 15904
rect 2827 15864 2872 15892
rect 2866 15852 2872 15864
rect 2924 15852 2930 15904
rect 3329 15895 3387 15901
rect 3329 15861 3341 15895
rect 3375 15892 3387 15895
rect 3878 15892 3884 15904
rect 3375 15864 3884 15892
rect 3375 15861 3387 15864
rect 3329 15855 3387 15861
rect 3878 15852 3884 15864
rect 3936 15852 3942 15904
rect 4080 15892 4108 15932
rect 5000 15932 7512 15960
rect 5000 15892 5028 15932
rect 6362 15892 6368 15904
rect 4080 15864 5028 15892
rect 6323 15864 6368 15892
rect 6362 15852 6368 15864
rect 6420 15852 6426 15904
rect 7374 15892 7380 15904
rect 7335 15864 7380 15892
rect 7374 15852 7380 15864
rect 7432 15852 7438 15904
rect 7484 15892 7512 15932
rect 7760 15932 8340 15960
rect 7760 15892 7788 15932
rect 8202 15892 8208 15904
rect 7484 15864 7788 15892
rect 8163 15864 8208 15892
rect 8202 15852 8208 15864
rect 8260 15852 8266 15904
rect 8312 15892 8340 15932
rect 10134 15920 10140 15972
rect 10192 15960 10198 15972
rect 15120 15960 15148 16204
rect 21818 16192 21824 16204
rect 21876 16192 21882 16244
rect 23750 16232 23756 16244
rect 21928 16204 23756 16232
rect 16206 16124 16212 16176
rect 16264 16164 16270 16176
rect 16264 16136 16988 16164
rect 16264 16124 16270 16136
rect 16850 16096 16856 16108
rect 16811 16068 16856 16096
rect 16850 16056 16856 16068
rect 16908 16056 16914 16108
rect 16960 16105 16988 16136
rect 17972 16136 19840 16164
rect 17972 16108 18000 16136
rect 16945 16099 17003 16105
rect 16945 16065 16957 16099
rect 16991 16065 17003 16099
rect 16945 16059 17003 16065
rect 17221 16099 17279 16105
rect 17221 16065 17233 16099
rect 17267 16096 17279 16099
rect 17770 16096 17776 16108
rect 17267 16068 17776 16096
rect 17267 16065 17279 16068
rect 17221 16059 17279 16065
rect 17770 16056 17776 16068
rect 17828 16056 17834 16108
rect 17954 16096 17960 16108
rect 17915 16068 17960 16096
rect 17954 16056 17960 16068
rect 18012 16056 18018 16108
rect 18046 16056 18052 16108
rect 18104 16096 18110 16108
rect 19812 16105 19840 16136
rect 20622 16124 20628 16176
rect 20680 16164 20686 16176
rect 21928 16164 21956 16204
rect 23750 16192 23756 16204
rect 23808 16192 23814 16244
rect 24026 16232 24032 16244
rect 23939 16204 24032 16232
rect 24026 16192 24032 16204
rect 24084 16232 24090 16244
rect 24670 16232 24676 16244
rect 24084 16204 24676 16232
rect 24084 16192 24090 16204
rect 24670 16192 24676 16204
rect 24728 16232 24734 16244
rect 25774 16232 25780 16244
rect 24728 16204 25544 16232
rect 25735 16204 25780 16232
rect 24728 16192 24734 16204
rect 22922 16164 22928 16176
rect 20680 16136 21956 16164
rect 22066 16136 22928 16164
rect 20680 16124 20686 16136
rect 18213 16099 18271 16105
rect 18213 16096 18225 16099
rect 18104 16068 18225 16096
rect 18104 16056 18110 16068
rect 18213 16065 18225 16068
rect 18259 16065 18271 16099
rect 18213 16059 18271 16065
rect 19797 16099 19855 16105
rect 19797 16065 19809 16099
rect 19843 16065 19855 16099
rect 19797 16059 19855 16065
rect 19886 16056 19892 16108
rect 19944 16096 19950 16108
rect 20053 16099 20111 16105
rect 20053 16096 20065 16099
rect 19944 16068 20065 16096
rect 19944 16056 19950 16068
rect 20053 16065 20065 16068
rect 20099 16065 20111 16099
rect 22066 16096 22094 16136
rect 22922 16124 22928 16136
rect 22980 16124 22986 16176
rect 20053 16059 20111 16065
rect 20824 16068 22094 16096
rect 22180 16099 22238 16105
rect 16114 16028 16120 16040
rect 16075 16000 16120 16028
rect 16114 15988 16120 16000
rect 16172 15988 16178 16040
rect 17126 16028 17132 16040
rect 17087 16000 17132 16028
rect 17126 15988 17132 16000
rect 17184 15988 17190 16040
rect 10192 15932 15148 15960
rect 10192 15920 10198 15932
rect 15930 15920 15936 15972
rect 15988 15960 15994 15972
rect 19334 15960 19340 15972
rect 15988 15932 17264 15960
rect 19295 15932 19340 15960
rect 15988 15920 15994 15932
rect 9122 15892 9128 15904
rect 8312 15864 9128 15892
rect 9122 15852 9128 15864
rect 9180 15852 9186 15904
rect 10318 15892 10324 15904
rect 10279 15864 10324 15892
rect 10318 15852 10324 15864
rect 10376 15852 10382 15904
rect 10781 15895 10839 15901
rect 10781 15861 10793 15895
rect 10827 15892 10839 15895
rect 13538 15892 13544 15904
rect 10827 15864 13544 15892
rect 10827 15861 10839 15864
rect 10781 15855 10839 15861
rect 13538 15852 13544 15864
rect 13596 15852 13602 15904
rect 13906 15892 13912 15904
rect 13867 15864 13912 15892
rect 13906 15852 13912 15864
rect 13964 15852 13970 15904
rect 16669 15895 16727 15901
rect 16669 15861 16681 15895
rect 16715 15892 16727 15895
rect 16850 15892 16856 15904
rect 16715 15864 16856 15892
rect 16715 15861 16727 15864
rect 16669 15855 16727 15861
rect 16850 15852 16856 15864
rect 16908 15852 16914 15904
rect 17236 15892 17264 15932
rect 19334 15920 19340 15932
rect 19392 15920 19398 15972
rect 20824 15892 20852 16068
rect 22180 16065 22192 16099
rect 22226 16096 22238 16099
rect 23198 16096 23204 16108
rect 22226 16068 23204 16096
rect 22226 16065 22238 16068
rect 22180 16059 22238 16065
rect 23198 16056 23204 16068
rect 23256 16056 23262 16108
rect 24044 16105 24072 16192
rect 25130 16124 25136 16176
rect 25188 16164 25194 16176
rect 25188 16136 25360 16164
rect 25188 16124 25194 16136
rect 24029 16099 24087 16105
rect 24029 16065 24041 16099
rect 24075 16065 24087 16099
rect 24029 16059 24087 16065
rect 24394 16056 24400 16108
rect 24452 16096 24458 16108
rect 24670 16096 24676 16108
rect 24452 16068 24676 16096
rect 24452 16056 24458 16068
rect 24670 16056 24676 16068
rect 24728 16096 24734 16108
rect 25332 16105 25360 16136
rect 25406 16124 25412 16176
rect 25464 16124 25470 16176
rect 25516 16164 25544 16204
rect 25774 16192 25780 16204
rect 25832 16192 25838 16244
rect 26510 16192 26516 16244
rect 26568 16232 26574 16244
rect 27249 16235 27307 16241
rect 27249 16232 27261 16235
rect 26568 16204 27261 16232
rect 26568 16192 26574 16204
rect 27249 16201 27261 16204
rect 27295 16201 27307 16235
rect 27249 16195 27307 16201
rect 25516 16136 25728 16164
rect 25041 16099 25099 16105
rect 25041 16096 25053 16099
rect 24728 16068 25053 16096
rect 24728 16056 24734 16068
rect 25041 16065 25053 16068
rect 25087 16065 25099 16099
rect 25041 16059 25099 16065
rect 25225 16099 25283 16105
rect 25225 16065 25237 16099
rect 25271 16065 25283 16099
rect 25225 16059 25283 16065
rect 25317 16099 25375 16105
rect 25317 16065 25329 16099
rect 25363 16065 25375 16099
rect 25424 16096 25452 16124
rect 25593 16099 25651 16105
rect 25593 16096 25605 16099
rect 25424 16068 25605 16096
rect 25317 16059 25375 16065
rect 25593 16065 25605 16068
rect 25639 16065 25651 16099
rect 25593 16059 25651 16065
rect 21910 16028 21916 16040
rect 21871 16000 21916 16028
rect 21910 15988 21916 16000
rect 21968 15988 21974 16040
rect 23750 16028 23756 16040
rect 23711 16000 23756 16028
rect 23750 15988 23756 16000
rect 23808 15988 23814 16040
rect 25240 15960 25268 16059
rect 25409 16031 25467 16037
rect 25409 15997 25421 16031
rect 25455 16028 25467 16031
rect 25700 16028 25728 16136
rect 25866 16056 25872 16108
rect 25924 16096 25930 16108
rect 26421 16099 26479 16105
rect 26421 16096 26433 16099
rect 25924 16068 26433 16096
rect 25924 16056 25930 16068
rect 26421 16065 26433 16068
rect 26467 16065 26479 16099
rect 26421 16059 26479 16065
rect 26510 16056 26516 16108
rect 26568 16096 26574 16108
rect 27157 16099 27215 16105
rect 27157 16096 27169 16099
rect 26568 16068 27169 16096
rect 26568 16056 26574 16068
rect 27157 16065 27169 16068
rect 27203 16065 27215 16099
rect 27157 16059 27215 16065
rect 25455 16000 25728 16028
rect 25455 15997 25467 16000
rect 25409 15991 25467 15997
rect 25682 15960 25688 15972
rect 25240 15932 25688 15960
rect 25682 15920 25688 15932
rect 25740 15920 25746 15972
rect 21174 15892 21180 15904
rect 17236 15864 20852 15892
rect 21135 15864 21180 15892
rect 21174 15852 21180 15864
rect 21232 15852 21238 15904
rect 23106 15852 23112 15904
rect 23164 15892 23170 15904
rect 23293 15895 23351 15901
rect 23293 15892 23305 15895
rect 23164 15864 23305 15892
rect 23164 15852 23170 15864
rect 23293 15861 23305 15864
rect 23339 15861 23351 15895
rect 26234 15892 26240 15904
rect 26195 15864 26240 15892
rect 23293 15855 23351 15861
rect 26234 15852 26240 15864
rect 26292 15852 26298 15904
rect 1104 15802 28060 15824
rect 1104 15750 5442 15802
rect 5494 15750 5506 15802
rect 5558 15750 5570 15802
rect 5622 15750 5634 15802
rect 5686 15750 5698 15802
rect 5750 15750 14428 15802
rect 14480 15750 14492 15802
rect 14544 15750 14556 15802
rect 14608 15750 14620 15802
rect 14672 15750 14684 15802
rect 14736 15750 23413 15802
rect 23465 15750 23477 15802
rect 23529 15750 23541 15802
rect 23593 15750 23605 15802
rect 23657 15750 23669 15802
rect 23721 15750 28060 15802
rect 1104 15728 28060 15750
rect 2774 15648 2780 15700
rect 2832 15688 2838 15700
rect 4154 15688 4160 15700
rect 2832 15660 2877 15688
rect 4115 15660 4160 15688
rect 2832 15648 2838 15660
rect 4154 15648 4160 15660
rect 4212 15648 4218 15700
rect 4982 15688 4988 15700
rect 4943 15660 4988 15688
rect 4982 15648 4988 15660
rect 5040 15648 5046 15700
rect 5166 15688 5172 15700
rect 5127 15660 5172 15688
rect 5166 15648 5172 15660
rect 5224 15648 5230 15700
rect 5810 15688 5816 15700
rect 5644 15660 5816 15688
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 2498 15512 2504 15564
rect 2556 15512 2562 15564
rect 5644 15561 5672 15660
rect 5810 15648 5816 15660
rect 5868 15648 5874 15700
rect 7374 15648 7380 15700
rect 7432 15688 7438 15700
rect 7834 15688 7840 15700
rect 7432 15660 7840 15688
rect 7432 15648 7438 15660
rect 7834 15648 7840 15660
rect 7892 15648 7898 15700
rect 7926 15648 7932 15700
rect 7984 15688 7990 15700
rect 8205 15691 8263 15697
rect 8205 15688 8217 15691
rect 7984 15660 8217 15688
rect 7984 15648 7990 15660
rect 8205 15657 8217 15660
rect 8251 15688 8263 15691
rect 10134 15688 10140 15700
rect 8251 15660 10140 15688
rect 8251 15657 8263 15660
rect 8205 15651 8263 15657
rect 10134 15648 10140 15660
rect 10192 15648 10198 15700
rect 10594 15688 10600 15700
rect 10555 15660 10600 15688
rect 10594 15648 10600 15660
rect 10652 15648 10658 15700
rect 11793 15691 11851 15697
rect 11793 15657 11805 15691
rect 11839 15688 11851 15691
rect 13354 15688 13360 15700
rect 11839 15660 13360 15688
rect 11839 15657 11851 15660
rect 11793 15651 11851 15657
rect 13354 15648 13360 15660
rect 13412 15648 13418 15700
rect 13455 15660 15286 15688
rect 7466 15580 7472 15632
rect 7524 15620 7530 15632
rect 7650 15620 7656 15632
rect 7524 15592 7656 15620
rect 7524 15580 7530 15592
rect 7650 15580 7656 15592
rect 7708 15580 7714 15632
rect 9214 15580 9220 15632
rect 9272 15580 9278 15632
rect 10502 15580 10508 15632
rect 10560 15620 10566 15632
rect 12342 15620 12348 15632
rect 10560 15592 12348 15620
rect 10560 15580 10566 15592
rect 12342 15580 12348 15592
rect 12400 15580 12406 15632
rect 13455 15620 13483 15660
rect 12728 15592 13483 15620
rect 14093 15623 14151 15629
rect 5629 15555 5687 15561
rect 5629 15521 5641 15555
rect 5675 15521 5687 15555
rect 5629 15515 5687 15521
rect 7006 15512 7012 15564
rect 7064 15552 7070 15564
rect 7834 15552 7840 15564
rect 7064 15524 7840 15552
rect 7064 15512 7070 15524
rect 7834 15512 7840 15524
rect 7892 15512 7898 15564
rect 8941 15555 8999 15561
rect 8941 15521 8953 15555
rect 8987 15552 8999 15555
rect 9232 15552 9260 15580
rect 8987 15524 9260 15552
rect 8987 15521 8999 15524
rect 8941 15515 8999 15521
rect 10594 15512 10600 15564
rect 10652 15552 10658 15564
rect 10778 15552 10784 15564
rect 10652 15524 10784 15552
rect 10652 15512 10658 15524
rect 10778 15512 10784 15524
rect 10836 15512 10842 15564
rect 11238 15512 11244 15564
rect 11296 15552 11302 15564
rect 11790 15552 11796 15564
rect 11296 15524 11796 15552
rect 11296 15512 11302 15524
rect 11790 15512 11796 15524
rect 11848 15512 11854 15564
rect 12618 15512 12624 15564
rect 12676 15552 12682 15564
rect 12728 15561 12756 15592
rect 14093 15589 14105 15623
rect 14139 15620 14151 15623
rect 15102 15620 15108 15632
rect 14139 15592 15108 15620
rect 14139 15589 14151 15592
rect 14093 15583 14151 15589
rect 15102 15580 15108 15592
rect 15160 15580 15166 15632
rect 12713 15555 12771 15561
rect 12713 15552 12725 15555
rect 12676 15524 12725 15552
rect 12676 15512 12682 15524
rect 12713 15521 12725 15524
rect 12759 15521 12771 15555
rect 12713 15515 12771 15521
rect 12802 15512 12808 15564
rect 12860 15552 12866 15564
rect 12860 15524 14873 15552
rect 12860 15512 12866 15524
rect 2516 15484 2544 15512
rect 4341 15487 4399 15493
rect 4341 15484 4353 15487
rect 2516 15456 4353 15484
rect 4341 15453 4353 15456
rect 4387 15484 4399 15487
rect 5896 15487 5954 15493
rect 4387 15456 5212 15484
rect 4387 15453 4399 15456
rect 4341 15447 4399 15453
rect 1664 15419 1722 15425
rect 1664 15385 1676 15419
rect 1710 15416 1722 15419
rect 1854 15416 1860 15428
rect 1710 15388 1860 15416
rect 1710 15385 1722 15388
rect 1664 15379 1722 15385
rect 1854 15376 1860 15388
rect 1912 15376 1918 15428
rect 4430 15376 4436 15428
rect 4488 15416 4494 15428
rect 4801 15419 4859 15425
rect 4801 15416 4813 15419
rect 4488 15388 4813 15416
rect 4488 15376 4494 15388
rect 4801 15385 4813 15388
rect 4847 15385 4859 15419
rect 5184 15416 5212 15456
rect 5896 15453 5908 15487
rect 5942 15484 5954 15487
rect 6362 15484 6368 15496
rect 5942 15456 6368 15484
rect 5942 15453 5954 15456
rect 5896 15447 5954 15453
rect 6362 15444 6368 15456
rect 6420 15444 6426 15496
rect 6454 15444 6460 15496
rect 6512 15484 6518 15496
rect 9217 15487 9275 15493
rect 9217 15484 9229 15487
rect 6512 15456 9229 15484
rect 6512 15444 6518 15456
rect 9217 15453 9229 15456
rect 9263 15484 9275 15487
rect 9582 15484 9588 15496
rect 9263 15456 9588 15484
rect 9263 15453 9275 15456
rect 9217 15447 9275 15453
rect 9582 15444 9588 15456
rect 9640 15484 9646 15496
rect 10229 15487 10287 15493
rect 10229 15484 10241 15487
rect 9640 15456 10241 15484
rect 9640 15444 9646 15456
rect 10229 15453 10241 15456
rect 10275 15453 10287 15487
rect 10229 15447 10287 15453
rect 10318 15444 10324 15496
rect 10376 15484 10382 15496
rect 11057 15487 11115 15493
rect 11057 15484 11069 15487
rect 10376 15456 11069 15484
rect 10376 15444 10382 15456
rect 11057 15453 11069 15456
rect 11103 15453 11115 15487
rect 11057 15447 11115 15453
rect 11146 15444 11152 15496
rect 11204 15484 11210 15496
rect 11977 15487 12035 15493
rect 11204 15456 11249 15484
rect 11204 15444 11210 15456
rect 11977 15453 11989 15487
rect 12023 15484 12035 15487
rect 12437 15487 12495 15493
rect 12437 15484 12449 15487
rect 12023 15456 12449 15484
rect 12023 15453 12035 15456
rect 11977 15447 12035 15453
rect 12437 15453 12449 15456
rect 12483 15484 12495 15487
rect 13722 15484 13728 15496
rect 12483 15456 13728 15484
rect 12483 15453 12495 15456
rect 12437 15447 12495 15453
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 14182 15444 14188 15496
rect 14240 15484 14246 15496
rect 14277 15487 14335 15493
rect 14277 15484 14289 15487
rect 14240 15456 14289 15484
rect 14240 15444 14246 15456
rect 14277 15453 14289 15456
rect 14323 15453 14335 15487
rect 14277 15447 14335 15453
rect 14366 15444 14372 15496
rect 14424 15484 14430 15496
rect 14734 15484 14740 15496
rect 14424 15456 14740 15484
rect 14424 15444 14430 15456
rect 14734 15444 14740 15456
rect 14792 15444 14798 15496
rect 14845 15493 14873 15524
rect 14830 15487 14888 15493
rect 14830 15453 14842 15487
rect 14876 15453 14888 15487
rect 15010 15484 15016 15496
rect 14971 15456 15016 15484
rect 14830 15447 14888 15453
rect 15010 15444 15016 15456
rect 15068 15444 15074 15496
rect 15258 15493 15286 15660
rect 15838 15648 15844 15700
rect 15896 15648 15902 15700
rect 16022 15688 16028 15700
rect 15983 15660 16028 15688
rect 16022 15648 16028 15660
rect 16080 15648 16086 15700
rect 16206 15648 16212 15700
rect 16264 15688 16270 15700
rect 16942 15688 16948 15700
rect 16264 15660 16948 15688
rect 16264 15648 16270 15660
rect 16942 15648 16948 15660
rect 17000 15648 17006 15700
rect 17770 15648 17776 15700
rect 17828 15688 17834 15700
rect 18141 15691 18199 15697
rect 18141 15688 18153 15691
rect 17828 15660 18153 15688
rect 17828 15648 17834 15660
rect 18141 15657 18153 15660
rect 18187 15657 18199 15691
rect 18141 15651 18199 15657
rect 19705 15691 19763 15697
rect 19705 15657 19717 15691
rect 19751 15688 19763 15691
rect 19886 15688 19892 15700
rect 19751 15660 19892 15688
rect 19751 15657 19763 15660
rect 19705 15651 19763 15657
rect 19886 15648 19892 15660
rect 19944 15648 19950 15700
rect 20809 15691 20867 15697
rect 20809 15657 20821 15691
rect 20855 15688 20867 15691
rect 20898 15688 20904 15700
rect 20855 15660 20904 15688
rect 20855 15657 20867 15660
rect 20809 15651 20867 15657
rect 20898 15648 20904 15660
rect 20956 15648 20962 15700
rect 22002 15648 22008 15700
rect 22060 15688 22066 15700
rect 22186 15688 22192 15700
rect 22060 15660 22192 15688
rect 22060 15648 22066 15660
rect 22186 15648 22192 15660
rect 22244 15648 22250 15700
rect 23198 15688 23204 15700
rect 23159 15660 23204 15688
rect 23198 15648 23204 15660
rect 23256 15648 23262 15700
rect 23569 15691 23627 15697
rect 23569 15657 23581 15691
rect 23615 15688 23627 15691
rect 24302 15688 24308 15700
rect 23615 15660 24308 15688
rect 23615 15657 23627 15660
rect 23569 15651 23627 15657
rect 24302 15648 24308 15660
rect 24360 15648 24366 15700
rect 25222 15648 25228 15700
rect 25280 15688 25286 15700
rect 25406 15688 25412 15700
rect 25280 15660 25412 15688
rect 25280 15648 25286 15660
rect 25406 15648 25412 15660
rect 25464 15648 25470 15700
rect 26878 15648 26884 15700
rect 26936 15688 26942 15700
rect 27341 15691 27399 15697
rect 27341 15688 27353 15691
rect 26936 15660 27353 15688
rect 26936 15648 26942 15660
rect 27341 15657 27353 15660
rect 27387 15657 27399 15691
rect 27341 15651 27399 15657
rect 15378 15620 15384 15632
rect 15339 15592 15384 15620
rect 15378 15580 15384 15592
rect 15436 15580 15442 15632
rect 15856 15620 15884 15648
rect 15764 15592 15884 15620
rect 15243 15487 15301 15493
rect 15243 15453 15255 15487
rect 15289 15484 15301 15487
rect 15654 15484 15660 15496
rect 15289 15456 15660 15484
rect 15289 15453 15301 15456
rect 15243 15447 15301 15453
rect 15654 15444 15660 15456
rect 15712 15444 15718 15496
rect 6822 15416 6828 15428
rect 5184 15388 6828 15416
rect 4801 15379 4859 15385
rect 6822 15376 6828 15388
rect 6880 15376 6886 15428
rect 8113 15419 8171 15425
rect 8113 15385 8125 15419
rect 8159 15385 8171 15419
rect 8113 15379 8171 15385
rect 10413 15419 10471 15425
rect 10413 15385 10425 15419
rect 10459 15416 10471 15419
rect 14550 15416 14556 15428
rect 10459 15388 14556 15416
rect 10459 15385 10471 15388
rect 10413 15379 10471 15385
rect 2314 15308 2320 15360
rect 2372 15348 2378 15360
rect 2590 15348 2596 15360
rect 2372 15320 2596 15348
rect 2372 15308 2378 15320
rect 2590 15308 2596 15320
rect 2648 15308 2654 15360
rect 5011 15351 5069 15357
rect 5011 15317 5023 15351
rect 5057 15348 5069 15351
rect 5166 15348 5172 15360
rect 5057 15320 5172 15348
rect 5057 15317 5069 15320
rect 5011 15311 5069 15317
rect 5166 15308 5172 15320
rect 5224 15308 5230 15360
rect 6362 15308 6368 15360
rect 6420 15348 6426 15360
rect 7009 15351 7067 15357
rect 7009 15348 7021 15351
rect 6420 15320 7021 15348
rect 6420 15308 6426 15320
rect 7009 15317 7021 15320
rect 7055 15317 7067 15351
rect 8128 15348 8156 15379
rect 14550 15376 14556 15388
rect 14608 15376 14614 15428
rect 14642 15376 14648 15428
rect 14700 15416 14706 15428
rect 15105 15419 15163 15425
rect 15105 15416 15117 15419
rect 14700 15388 15117 15416
rect 14700 15376 14706 15388
rect 15105 15385 15117 15388
rect 15151 15385 15163 15419
rect 15764 15416 15792 15592
rect 19610 15580 19616 15632
rect 19668 15620 19674 15632
rect 20073 15623 20131 15629
rect 20073 15620 20085 15623
rect 19668 15592 20085 15620
rect 19668 15580 19674 15592
rect 20073 15589 20085 15592
rect 20119 15589 20131 15623
rect 20073 15583 20131 15589
rect 20622 15580 20628 15632
rect 20680 15620 20686 15632
rect 22094 15620 22100 15632
rect 20680 15592 20852 15620
rect 20680 15580 20686 15592
rect 15838 15512 15844 15564
rect 15896 15512 15902 15564
rect 20714 15552 20720 15564
rect 19904 15524 20720 15552
rect 15856 15484 15884 15512
rect 16761 15487 16819 15493
rect 15856 15459 16084 15484
rect 15856 15456 16129 15459
rect 16056 15453 16129 15456
rect 15841 15419 15899 15425
rect 16056 15422 16083 15453
rect 15841 15416 15853 15419
rect 15764 15388 15853 15416
rect 15105 15379 15163 15385
rect 15841 15385 15853 15388
rect 15887 15385 15899 15419
rect 16071 15419 16083 15422
rect 16117 15419 16129 15453
rect 16761 15453 16773 15487
rect 16807 15484 16819 15487
rect 17954 15484 17960 15496
rect 16807 15456 17960 15484
rect 16807 15453 16819 15456
rect 16761 15447 16819 15453
rect 17954 15444 17960 15456
rect 18012 15444 18018 15496
rect 19904 15493 19932 15524
rect 20714 15512 20720 15524
rect 20772 15512 20778 15564
rect 20824 15552 20852 15592
rect 21468 15592 22100 15620
rect 21468 15561 21496 15592
rect 22094 15580 22100 15592
rect 22152 15620 22158 15632
rect 22152 15592 22508 15620
rect 22152 15580 22158 15592
rect 21453 15555 21511 15561
rect 20824 15524 21404 15552
rect 19889 15487 19947 15493
rect 19889 15453 19901 15487
rect 19935 15453 19947 15487
rect 19889 15447 19947 15453
rect 20070 15444 20076 15496
rect 20128 15484 20134 15496
rect 20165 15487 20223 15493
rect 20165 15484 20177 15487
rect 20128 15456 20177 15484
rect 20128 15444 20134 15456
rect 20165 15453 20177 15456
rect 20211 15484 20223 15487
rect 21174 15484 21180 15496
rect 20211 15456 21180 15484
rect 20211 15453 20223 15456
rect 20165 15447 20223 15453
rect 21174 15444 21180 15456
rect 21232 15484 21238 15496
rect 21269 15487 21327 15493
rect 21269 15484 21281 15487
rect 21232 15456 21281 15484
rect 21232 15444 21238 15456
rect 21269 15453 21281 15456
rect 21315 15453 21327 15487
rect 21376 15484 21404 15524
rect 21453 15521 21465 15555
rect 21499 15521 21511 15555
rect 22373 15555 22431 15561
rect 22373 15552 22385 15555
rect 21453 15515 21511 15521
rect 21652 15524 22385 15552
rect 21652 15484 21680 15524
rect 22373 15521 22385 15524
rect 22419 15521 22431 15555
rect 22480 15552 22508 15592
rect 22922 15580 22928 15632
rect 22980 15620 22986 15632
rect 22980 15592 24440 15620
rect 22980 15580 22986 15592
rect 23198 15552 23204 15564
rect 22480 15524 23204 15552
rect 22373 15515 22431 15521
rect 23198 15512 23204 15524
rect 23256 15512 23262 15564
rect 23658 15552 23664 15564
rect 23619 15524 23664 15552
rect 23658 15512 23664 15524
rect 23716 15512 23722 15564
rect 24412 15561 24440 15592
rect 24397 15555 24455 15561
rect 24397 15521 24409 15555
rect 24443 15521 24455 15555
rect 24670 15552 24676 15564
rect 24631 15524 24676 15552
rect 24397 15515 24455 15521
rect 24670 15512 24676 15524
rect 24728 15512 24734 15564
rect 25958 15552 25964 15564
rect 25919 15524 25964 15552
rect 25958 15512 25964 15524
rect 26016 15512 26022 15564
rect 21376 15456 21680 15484
rect 21269 15447 21327 15453
rect 21818 15444 21824 15496
rect 21876 15484 21882 15496
rect 22002 15484 22008 15496
rect 21876 15456 22008 15484
rect 21876 15444 21882 15456
rect 22002 15444 22008 15456
rect 22060 15444 22066 15496
rect 22186 15484 22192 15496
rect 22147 15456 22192 15484
rect 22186 15444 22192 15456
rect 22244 15444 22250 15496
rect 22281 15487 22339 15493
rect 22281 15453 22293 15487
rect 22327 15453 22339 15487
rect 22281 15447 22339 15453
rect 22557 15487 22615 15493
rect 22557 15453 22569 15487
rect 22603 15453 22615 15487
rect 22557 15447 22615 15453
rect 16071 15413 16129 15419
rect 17028 15419 17086 15425
rect 15841 15379 15899 15385
rect 17028 15385 17040 15419
rect 17074 15416 17086 15419
rect 21082 15416 21088 15428
rect 17074 15388 21088 15416
rect 17074 15385 17086 15388
rect 17028 15379 17086 15385
rect 21082 15376 21088 15388
rect 21140 15376 21146 15428
rect 22296 15416 22324 15447
rect 22204 15388 22324 15416
rect 22572 15416 22600 15447
rect 23290 15444 23296 15496
rect 23348 15484 23354 15496
rect 23385 15487 23443 15493
rect 23385 15484 23397 15487
rect 23348 15456 23397 15484
rect 23348 15444 23354 15456
rect 23385 15453 23397 15456
rect 23431 15453 23443 15487
rect 23385 15447 23443 15453
rect 23842 15444 23848 15496
rect 23900 15444 23906 15496
rect 23860 15416 23888 15444
rect 22572 15388 23888 15416
rect 26228 15419 26286 15425
rect 22204 15360 22232 15388
rect 26228 15385 26240 15419
rect 26274 15416 26286 15419
rect 26326 15416 26332 15428
rect 26274 15388 26332 15416
rect 26274 15385 26286 15388
rect 26228 15379 26286 15385
rect 26326 15376 26332 15388
rect 26384 15376 26390 15428
rect 8294 15348 8300 15360
rect 8128 15320 8300 15348
rect 7009 15311 7067 15317
rect 8294 15308 8300 15320
rect 8352 15348 8358 15360
rect 15930 15348 15936 15360
rect 8352 15320 15936 15348
rect 8352 15308 8358 15320
rect 15930 15308 15936 15320
rect 15988 15308 15994 15360
rect 16209 15351 16267 15357
rect 16209 15317 16221 15351
rect 16255 15348 16267 15351
rect 16942 15348 16948 15360
rect 16255 15320 16948 15348
rect 16255 15317 16267 15320
rect 16209 15311 16267 15317
rect 16942 15308 16948 15320
rect 17000 15308 17006 15360
rect 19334 15308 19340 15360
rect 19392 15348 19398 15360
rect 20622 15348 20628 15360
rect 19392 15320 20628 15348
rect 19392 15308 19398 15320
rect 20622 15308 20628 15320
rect 20680 15308 20686 15360
rect 20714 15308 20720 15360
rect 20772 15348 20778 15360
rect 21177 15351 21235 15357
rect 21177 15348 21189 15351
rect 20772 15320 21189 15348
rect 20772 15308 20778 15320
rect 21177 15317 21189 15320
rect 21223 15317 21235 15351
rect 21177 15311 21235 15317
rect 22186 15308 22192 15360
rect 22244 15308 22250 15360
rect 22741 15351 22799 15357
rect 22741 15317 22753 15351
rect 22787 15348 22799 15351
rect 23842 15348 23848 15360
rect 22787 15320 23848 15348
rect 22787 15317 22799 15320
rect 22741 15311 22799 15317
rect 23842 15308 23848 15320
rect 23900 15308 23906 15360
rect 25222 15308 25228 15360
rect 25280 15348 25286 15360
rect 25866 15348 25872 15360
rect 25280 15320 25872 15348
rect 25280 15308 25286 15320
rect 25866 15308 25872 15320
rect 25924 15308 25930 15360
rect 1104 15258 28060 15280
rect 1104 15206 9935 15258
rect 9987 15206 9999 15258
rect 10051 15206 10063 15258
rect 10115 15206 10127 15258
rect 10179 15206 10191 15258
rect 10243 15206 18920 15258
rect 18972 15206 18984 15258
rect 19036 15206 19048 15258
rect 19100 15206 19112 15258
rect 19164 15206 19176 15258
rect 19228 15206 28060 15258
rect 1104 15184 28060 15206
rect 1394 15104 1400 15156
rect 1452 15144 1458 15156
rect 1670 15144 1676 15156
rect 1452 15116 1676 15144
rect 1452 15104 1458 15116
rect 1670 15104 1676 15116
rect 1728 15104 1734 15156
rect 1854 15144 1860 15156
rect 1815 15116 1860 15144
rect 1854 15104 1860 15116
rect 1912 15104 1918 15156
rect 2501 15147 2559 15153
rect 2501 15113 2513 15147
rect 2547 15144 2559 15147
rect 5166 15144 5172 15156
rect 5224 15153 5230 15156
rect 5224 15147 5253 15153
rect 2547 15116 4384 15144
rect 5105 15116 5172 15144
rect 2547 15113 2559 15116
rect 2501 15107 2559 15113
rect 2866 15076 2872 15088
rect 2056 15048 2872 15076
rect 2056 15017 2084 15048
rect 2866 15036 2872 15048
rect 2924 15036 2930 15088
rect 2041 15011 2099 15017
rect 2041 14977 2053 15011
rect 2087 14977 2099 15011
rect 3412 15011 3470 15017
rect 2041 14971 2099 14977
rect 2685 14995 2743 15001
rect 2685 14961 2697 14995
rect 2731 14961 2743 14995
rect 3412 14977 3424 15011
rect 3458 15008 3470 15011
rect 3786 15008 3792 15020
rect 3458 14980 3792 15008
rect 3458 14977 3470 14980
rect 3412 14971 3470 14977
rect 3786 14968 3792 14980
rect 3844 14968 3850 15020
rect 4356 15008 4384 15116
rect 5166 15104 5172 15116
rect 5241 15144 5253 15147
rect 6454 15144 6460 15156
rect 5241 15116 6460 15144
rect 5241 15113 5253 15116
rect 5224 15107 5253 15113
rect 5224 15104 5230 15107
rect 6454 15104 6460 15116
rect 6512 15144 6518 15156
rect 6565 15147 6623 15153
rect 6565 15144 6577 15147
rect 6512 15116 6577 15144
rect 6512 15104 6518 15116
rect 6565 15113 6577 15116
rect 6611 15113 6623 15147
rect 6730 15144 6736 15156
rect 6691 15116 6736 15144
rect 6565 15107 6623 15113
rect 6730 15104 6736 15116
rect 6788 15104 6794 15156
rect 6822 15104 6828 15156
rect 6880 15144 6886 15156
rect 7469 15147 7527 15153
rect 7469 15144 7481 15147
rect 6880 15116 7481 15144
rect 6880 15104 6886 15116
rect 7469 15113 7481 15116
rect 7515 15113 7527 15147
rect 7469 15107 7527 15113
rect 8205 15147 8263 15153
rect 8205 15113 8217 15147
rect 8251 15144 8263 15147
rect 8294 15144 8300 15156
rect 8251 15116 8300 15144
rect 8251 15113 8263 15116
rect 8205 15107 8263 15113
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 9125 15147 9183 15153
rect 9125 15113 9137 15147
rect 9171 15144 9183 15147
rect 9214 15144 9220 15156
rect 9171 15116 9220 15144
rect 9171 15113 9183 15116
rect 9125 15107 9183 15113
rect 4430 15036 4436 15088
rect 4488 15076 4494 15088
rect 4985 15079 5043 15085
rect 4985 15076 4997 15079
rect 4488 15048 4997 15076
rect 4488 15036 4494 15048
rect 4985 15045 4997 15048
rect 5031 15076 5043 15079
rect 6365 15079 6423 15085
rect 6365 15076 6377 15079
rect 5031 15048 6377 15076
rect 5031 15045 5043 15048
rect 4985 15039 5043 15045
rect 6365 15045 6377 15048
rect 6411 15076 6423 15079
rect 9140 15076 9168 15107
rect 9214 15104 9220 15116
rect 9272 15104 9278 15156
rect 10873 15147 10931 15153
rect 9600 15116 10824 15144
rect 6411 15048 7144 15076
rect 6411 15045 6423 15048
rect 6365 15039 6423 15045
rect 4356 14980 6960 15008
rect 2685 14955 2743 14961
rect 2700 14884 2728 14955
rect 3145 14943 3203 14949
rect 3145 14909 3157 14943
rect 3191 14909 3203 14943
rect 3145 14903 3203 14909
rect 2682 14832 2688 14884
rect 2740 14832 2746 14884
rect 3160 14804 3188 14903
rect 4154 14832 4160 14884
rect 4212 14872 4218 14884
rect 5353 14875 5411 14881
rect 5353 14872 5365 14875
rect 4212 14844 5365 14872
rect 4212 14832 4218 14844
rect 5353 14841 5365 14844
rect 5399 14841 5411 14875
rect 5353 14835 5411 14841
rect 4338 14804 4344 14816
rect 3160 14776 4344 14804
rect 4338 14764 4344 14776
rect 4396 14764 4402 14816
rect 4525 14807 4583 14813
rect 4525 14773 4537 14807
rect 4571 14804 4583 14807
rect 5169 14807 5227 14813
rect 5169 14804 5181 14807
rect 4571 14776 5181 14804
rect 4571 14773 4583 14776
rect 4525 14767 4583 14773
rect 5169 14773 5181 14776
rect 5215 14773 5227 14807
rect 5169 14767 5227 14773
rect 6362 14764 6368 14816
rect 6420 14804 6426 14816
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 6420 14776 6561 14804
rect 6420 14764 6426 14776
rect 6549 14773 6561 14776
rect 6595 14773 6607 14807
rect 6932 14804 6960 14980
rect 7116 14872 7144 15048
rect 7392 15048 9168 15076
rect 7392 15017 7420 15048
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 14977 7435 15011
rect 7377 14971 7435 14977
rect 7561 15011 7619 15017
rect 7561 14977 7573 15011
rect 7607 14977 7619 15011
rect 7561 14971 7619 14977
rect 7576 14940 7604 14971
rect 7926 14968 7932 15020
rect 7984 15008 7990 15020
rect 8113 15011 8171 15017
rect 8113 15008 8125 15011
rect 7984 14980 8125 15008
rect 7984 14968 7990 14980
rect 8113 14977 8125 14980
rect 8159 14977 8171 15011
rect 8113 14971 8171 14977
rect 8202 14968 8208 15020
rect 8260 15008 8266 15020
rect 8260 14980 8616 15008
rect 8260 14968 8266 14980
rect 8294 14940 8300 14952
rect 7576 14912 8300 14940
rect 8294 14900 8300 14912
rect 8352 14900 8358 14952
rect 8588 14940 8616 14980
rect 8662 14968 8668 15020
rect 8720 15008 8726 15020
rect 8757 15011 8815 15017
rect 8757 15008 8769 15011
rect 8720 14980 8769 15008
rect 8720 14968 8726 14980
rect 8757 14977 8769 14980
rect 8803 14977 8815 15011
rect 9600 15008 9628 15116
rect 9766 15036 9772 15088
rect 9824 15076 9830 15088
rect 9861 15079 9919 15085
rect 9861 15076 9873 15079
rect 9824 15048 9873 15076
rect 9824 15036 9830 15048
rect 9861 15045 9873 15048
rect 9907 15045 9919 15079
rect 10796 15076 10824 15116
rect 10873 15113 10885 15147
rect 10919 15144 10931 15147
rect 13107 15147 13165 15153
rect 13107 15144 13119 15147
rect 10919 15116 13119 15144
rect 10919 15113 10931 15116
rect 10873 15107 10931 15113
rect 13107 15113 13119 15116
rect 13153 15144 13165 15147
rect 13722 15144 13728 15156
rect 13153 15116 13728 15144
rect 13153 15113 13165 15116
rect 13107 15107 13165 15113
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 14385 15147 14443 15153
rect 14385 15144 14397 15147
rect 14108 15116 14397 15144
rect 11517 15079 11575 15085
rect 10796 15048 10907 15076
rect 9861 15039 9919 15045
rect 8757 14971 8815 14977
rect 8864 14980 9628 15008
rect 8864 14949 8892 14980
rect 9674 14968 9680 15020
rect 9732 15008 9738 15020
rect 10594 15008 10600 15020
rect 9732 14980 10600 15008
rect 9732 14968 9738 14980
rect 10594 14968 10600 14980
rect 10652 15008 10658 15020
rect 10781 15011 10839 15017
rect 10781 15008 10793 15011
rect 10652 14980 10793 15008
rect 10652 14968 10658 14980
rect 10781 14977 10793 14980
rect 10827 14977 10839 15011
rect 10879 15008 10907 15048
rect 11517 15045 11529 15079
rect 11563 15045 11575 15079
rect 11517 15039 11575 15045
rect 11733 15079 11791 15085
rect 11733 15045 11745 15079
rect 11779 15076 11791 15079
rect 11779 15048 12296 15076
rect 11779 15045 11791 15048
rect 11733 15039 11791 15045
rect 10965 15011 11023 15017
rect 10965 15008 10977 15011
rect 10879 14980 10977 15008
rect 10781 14971 10839 14977
rect 10965 14977 10977 14980
rect 11011 15008 11023 15011
rect 11330 15008 11336 15020
rect 11011 14980 11336 15008
rect 11011 14977 11023 14980
rect 10965 14971 11023 14977
rect 11330 14968 11336 14980
rect 11388 14968 11394 15020
rect 8849 14943 8907 14949
rect 8849 14940 8861 14943
rect 8588 14912 8861 14940
rect 8849 14909 8861 14912
rect 8895 14909 8907 14943
rect 10870 14940 10876 14952
rect 8849 14903 8907 14909
rect 8956 14912 10876 14940
rect 8956 14872 8984 14912
rect 10870 14900 10876 14912
rect 10928 14900 10934 14952
rect 11422 14900 11428 14952
rect 11480 14940 11486 14952
rect 11532 14940 11560 15039
rect 12268 15008 12296 15048
rect 12342 15036 12348 15088
rect 12400 15076 12406 15088
rect 12897 15079 12955 15085
rect 12897 15076 12909 15079
rect 12400 15048 12909 15076
rect 12400 15036 12406 15048
rect 12897 15045 12909 15048
rect 12943 15045 12955 15079
rect 12897 15039 12955 15045
rect 13354 15036 13360 15088
rect 13412 15076 13418 15088
rect 14108 15076 14136 15116
rect 14385 15113 14397 15116
rect 14431 15144 14443 15147
rect 15838 15144 15844 15156
rect 15896 15153 15902 15156
rect 15896 15147 15915 15153
rect 14431 15116 15844 15144
rect 14431 15113 14443 15116
rect 14385 15107 14443 15113
rect 15838 15104 15844 15116
rect 15903 15113 15915 15147
rect 15896 15107 15915 15113
rect 16025 15147 16083 15153
rect 16025 15113 16037 15147
rect 16071 15113 16083 15147
rect 16025 15107 16083 15113
rect 17129 15147 17187 15153
rect 17129 15113 17141 15147
rect 17175 15144 17187 15147
rect 19334 15144 19340 15156
rect 17175 15116 19340 15144
rect 17175 15113 17187 15116
rect 17129 15107 17187 15113
rect 15896 15104 15902 15107
rect 13412 15048 14136 15076
rect 14185 15079 14243 15085
rect 13412 15036 13418 15048
rect 14185 15045 14197 15079
rect 14231 15045 14243 15079
rect 14185 15039 14243 15045
rect 15657 15079 15715 15085
rect 15657 15045 15669 15079
rect 15703 15076 15715 15079
rect 16040 15076 16068 15107
rect 19334 15104 19340 15116
rect 19392 15104 19398 15156
rect 19521 15147 19579 15153
rect 19521 15113 19533 15147
rect 19567 15144 19579 15147
rect 26237 15147 26295 15153
rect 26237 15144 26249 15147
rect 19567 15116 20096 15144
rect 19567 15113 19579 15116
rect 19521 15107 19579 15113
rect 20068 15076 20096 15116
rect 20364 15116 20760 15144
rect 20257 15079 20315 15085
rect 15703 15048 16008 15076
rect 16040 15048 20024 15076
rect 20068 15048 20208 15076
rect 15703 15045 15715 15048
rect 15657 15039 15715 15045
rect 12618 15008 12624 15020
rect 12268 14980 12624 15008
rect 12618 14968 12624 14980
rect 12676 14968 12682 15020
rect 13078 14968 13084 15020
rect 13136 15008 13142 15020
rect 13722 15008 13728 15020
rect 13136 14980 13728 15008
rect 13136 14968 13142 14980
rect 13722 14968 13728 14980
rect 13780 14968 13786 15020
rect 11698 14940 11704 14952
rect 11480 14912 11704 14940
rect 11480 14900 11486 14912
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 13262 14940 13268 14952
rect 11900 14912 13268 14940
rect 7116 14844 8984 14872
rect 9858 14832 9864 14884
rect 9916 14872 9922 14884
rect 10778 14872 10784 14884
rect 9916 14844 10784 14872
rect 9916 14832 9922 14844
rect 10778 14832 10784 14844
rect 10836 14832 10842 14884
rect 11900 14881 11928 14912
rect 13262 14900 13268 14912
rect 13320 14900 13326 14952
rect 11885 14875 11943 14881
rect 11885 14841 11897 14875
rect 11931 14841 11943 14875
rect 11885 14835 11943 14841
rect 12158 14832 12164 14884
rect 12216 14872 12222 14884
rect 14200 14872 14228 15039
rect 14826 15008 14832 15020
rect 12216 14844 14228 14872
rect 14292 14980 14832 15008
rect 12216 14832 12222 14844
rect 7834 14804 7840 14816
rect 6932 14776 7840 14804
rect 6549 14767 6607 14773
rect 7834 14764 7840 14776
rect 7892 14764 7898 14816
rect 8941 14807 8999 14813
rect 8941 14773 8953 14807
rect 8987 14804 8999 14807
rect 9674 14804 9680 14816
rect 8987 14776 9680 14804
rect 8987 14773 8999 14776
rect 8941 14767 8999 14773
rect 9674 14764 9680 14776
rect 9732 14764 9738 14816
rect 9953 14807 10011 14813
rect 9953 14773 9965 14807
rect 9999 14804 10011 14807
rect 11330 14804 11336 14816
rect 9999 14776 11336 14804
rect 9999 14773 10011 14776
rect 9953 14767 10011 14773
rect 11330 14764 11336 14776
rect 11388 14764 11394 14816
rect 11698 14804 11704 14816
rect 11659 14776 11704 14804
rect 11698 14764 11704 14776
rect 11756 14764 11762 14816
rect 13078 14804 13084 14816
rect 13039 14776 13084 14804
rect 13078 14764 13084 14776
rect 13136 14764 13142 14816
rect 13265 14807 13323 14813
rect 13265 14773 13277 14807
rect 13311 14804 13323 14807
rect 14292 14804 14320 14980
rect 14826 14968 14832 14980
rect 14884 14968 14890 15020
rect 15197 15011 15255 15017
rect 15197 14977 15209 15011
rect 15243 15008 15255 15011
rect 15980 15008 16008 15048
rect 16574 15008 16580 15020
rect 15243 14980 15900 15008
rect 15980 14980 16580 15008
rect 15243 14977 15255 14980
rect 15197 14971 15255 14977
rect 14384 14912 15516 14940
rect 14384 14813 14412 14912
rect 14553 14875 14611 14881
rect 14553 14841 14565 14875
rect 14599 14872 14611 14875
rect 15378 14872 15384 14884
rect 14599 14844 15384 14872
rect 14599 14841 14611 14844
rect 14553 14835 14611 14841
rect 15378 14832 15384 14844
rect 15436 14832 15442 14884
rect 13311 14776 14320 14804
rect 14369 14807 14427 14813
rect 13311 14773 13323 14776
rect 13265 14767 13323 14773
rect 14369 14773 14381 14807
rect 14415 14773 14427 14807
rect 15010 14804 15016 14816
rect 14971 14776 15016 14804
rect 14369 14767 14427 14773
rect 15010 14764 15016 14776
rect 15068 14764 15074 14816
rect 15488 14804 15516 14912
rect 15872 14872 15900 14980
rect 16574 14968 16580 14980
rect 16632 14968 16638 15020
rect 16761 15011 16819 15017
rect 16761 14977 16773 15011
rect 16807 14977 16819 15011
rect 16761 14971 16819 14977
rect 16776 14940 16804 14971
rect 16850 14968 16856 15020
rect 16908 15008 16914 15020
rect 16945 15011 17003 15017
rect 16945 15008 16957 15011
rect 16908 14980 16957 15008
rect 16908 14968 16914 14980
rect 16945 14977 16957 14980
rect 16991 15008 17003 15011
rect 17402 15008 17408 15020
rect 16991 14980 17408 15008
rect 16991 14977 17003 14980
rect 16945 14971 17003 14977
rect 17402 14968 17408 14980
rect 17460 14968 17466 15020
rect 17954 14968 17960 15020
rect 18012 15008 18018 15020
rect 18141 15011 18199 15017
rect 18141 15008 18153 15011
rect 18012 14980 18153 15008
rect 18012 14968 18018 14980
rect 18141 14977 18153 14980
rect 18187 14977 18199 15011
rect 18141 14971 18199 14977
rect 18408 15011 18466 15017
rect 18408 14977 18420 15011
rect 18454 15008 18466 15011
rect 18690 15008 18696 15020
rect 18454 14980 18696 15008
rect 18454 14977 18466 14980
rect 18408 14971 18466 14977
rect 18690 14968 18696 14980
rect 18748 14968 18754 15020
rect 19996 15017 20024 15048
rect 19981 15011 20039 15017
rect 19981 14977 19993 15011
rect 20027 14977 20039 15011
rect 19981 14971 20039 14977
rect 20074 15011 20132 15017
rect 20074 14977 20086 15011
rect 20120 14977 20132 15011
rect 20074 14971 20132 14977
rect 17862 14940 17868 14952
rect 16776 14912 17868 14940
rect 17862 14900 17868 14912
rect 17920 14900 17926 14952
rect 19886 14900 19892 14952
rect 19944 14940 19950 14952
rect 20088 14940 20116 14971
rect 19944 14912 20116 14940
rect 20180 14940 20208 15048
rect 20257 15045 20269 15079
rect 20303 15076 20315 15079
rect 20364 15076 20392 15116
rect 20732 15088 20760 15116
rect 22020 15116 26249 15144
rect 20303 15048 20392 15076
rect 20303 15045 20315 15048
rect 20257 15039 20315 15045
rect 20714 15036 20720 15088
rect 20772 15036 20778 15088
rect 20349 15011 20407 15017
rect 20349 14977 20361 15011
rect 20395 14977 20407 15011
rect 20349 14971 20407 14977
rect 20487 15011 20545 15017
rect 20487 14977 20499 15011
rect 20533 15008 20545 15011
rect 20533 15006 20668 15008
rect 20533 14980 20760 15006
rect 20533 14977 20545 14980
rect 20640 14978 20760 14980
rect 20487 14971 20545 14977
rect 20364 14940 20392 14971
rect 20180 14912 20392 14940
rect 20732 14940 20760 14978
rect 20806 14968 20812 15020
rect 20864 15008 20870 15020
rect 22020 15017 22048 15116
rect 26237 15113 26249 15116
rect 26283 15113 26295 15147
rect 26237 15107 26295 15113
rect 22112 15048 27200 15076
rect 21269 15011 21327 15017
rect 21269 15008 21281 15011
rect 20864 14980 21281 15008
rect 20864 14968 20870 14980
rect 21269 14977 21281 14980
rect 21315 14977 21327 15011
rect 21269 14971 21327 14977
rect 22005 15011 22063 15017
rect 22005 14977 22017 15011
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 21174 14940 21180 14952
rect 20732 14912 21180 14940
rect 19944 14900 19950 14912
rect 21174 14900 21180 14912
rect 21232 14900 21238 14952
rect 16206 14872 16212 14884
rect 15872 14844 16212 14872
rect 16206 14832 16212 14844
rect 16264 14832 16270 14884
rect 16666 14832 16672 14884
rect 16724 14872 16730 14884
rect 16850 14872 16856 14884
rect 16724 14844 16856 14872
rect 16724 14832 16730 14844
rect 16850 14832 16856 14844
rect 16908 14832 16914 14884
rect 22112 14872 22140 15048
rect 22186 14968 22192 15020
rect 22244 15010 22250 15020
rect 22281 15011 22339 15017
rect 22281 15010 22293 15011
rect 22244 14982 22293 15010
rect 22244 14968 22250 14982
rect 22281 14977 22293 14982
rect 22327 15010 22339 15011
rect 22327 15008 22407 15010
rect 23106 15008 23112 15020
rect 22327 14982 23112 15008
rect 22327 14977 22339 14982
rect 22379 14980 23112 14982
rect 22281 14971 22339 14977
rect 23106 14968 23112 14980
rect 23164 14968 23170 15020
rect 23201 15011 23259 15017
rect 23201 14977 23213 15011
rect 23247 15008 23259 15011
rect 24394 15008 24400 15020
rect 23247 14980 24400 15008
rect 23247 14977 23259 14980
rect 23201 14971 23259 14977
rect 24394 14968 24400 14980
rect 24452 14968 24458 15020
rect 24670 14968 24676 15020
rect 24728 15008 24734 15020
rect 25501 15011 25559 15017
rect 25501 15008 25513 15011
rect 24728 14980 25513 15008
rect 24728 14968 24734 14980
rect 25501 14977 25513 14980
rect 25547 14977 25559 15011
rect 25682 15008 25688 15020
rect 25643 14980 25688 15008
rect 25501 14971 25559 14977
rect 25682 14968 25688 14980
rect 25740 14968 25746 15020
rect 26053 15011 26111 15017
rect 26053 14977 26065 15011
rect 26099 15008 26111 15011
rect 26142 15008 26148 15020
rect 26099 14980 26148 15008
rect 26099 14977 26111 14980
rect 26053 14971 26111 14977
rect 26142 14968 26148 14980
rect 26200 14968 26206 15020
rect 27172 15017 27200 15048
rect 27157 15011 27215 15017
rect 27157 14977 27169 15011
rect 27203 14977 27215 15011
rect 27157 14971 27215 14977
rect 22554 14900 22560 14952
rect 22612 14940 22618 14952
rect 23290 14940 23296 14952
rect 22612 14912 22784 14940
rect 23251 14912 23296 14940
rect 22612 14900 22618 14912
rect 22756 14881 22784 14912
rect 23290 14900 23296 14912
rect 23348 14900 23354 14952
rect 24213 14943 24271 14949
rect 24213 14940 24225 14943
rect 23400 14912 24225 14940
rect 16960 14844 17264 14872
rect 15841 14807 15899 14813
rect 15841 14804 15853 14807
rect 15488 14776 15853 14804
rect 15841 14773 15853 14776
rect 15887 14804 15899 14807
rect 16022 14804 16028 14816
rect 15887 14776 16028 14804
rect 15887 14773 15899 14776
rect 15841 14767 15899 14773
rect 16022 14764 16028 14776
rect 16080 14764 16086 14816
rect 16390 14764 16396 14816
rect 16448 14804 16454 14816
rect 16960 14804 16988 14844
rect 16448 14776 16988 14804
rect 17236 14804 17264 14844
rect 19076 14844 22140 14872
rect 22741 14875 22799 14881
rect 19076 14804 19104 14844
rect 22741 14841 22753 14875
rect 22787 14841 22799 14875
rect 22741 14835 22799 14841
rect 23198 14832 23204 14884
rect 23256 14872 23262 14884
rect 23400 14872 23428 14912
rect 24213 14909 24225 14912
rect 24259 14909 24271 14943
rect 24213 14903 24271 14909
rect 24489 14943 24547 14949
rect 24489 14909 24501 14943
rect 24535 14940 24547 14943
rect 25130 14940 25136 14952
rect 24535 14912 25136 14940
rect 24535 14909 24547 14912
rect 24489 14903 24547 14909
rect 25130 14900 25136 14912
rect 25188 14940 25194 14952
rect 25700 14940 25728 14968
rect 25188 14912 25728 14940
rect 25777 14943 25835 14949
rect 25188 14900 25194 14912
rect 25777 14909 25789 14943
rect 25823 14909 25835 14943
rect 25777 14903 25835 14909
rect 23256 14844 23428 14872
rect 23256 14832 23262 14844
rect 23474 14832 23480 14884
rect 23532 14872 23538 14884
rect 25792 14872 25820 14903
rect 25866 14900 25872 14952
rect 25924 14940 25930 14952
rect 25924 14912 25969 14940
rect 25924 14900 25930 14912
rect 23532 14844 25820 14872
rect 26973 14875 27031 14881
rect 23532 14832 23538 14844
rect 26973 14841 26985 14875
rect 27019 14841 27031 14875
rect 26973 14835 27031 14841
rect 17236 14776 19104 14804
rect 16448 14764 16454 14776
rect 19150 14764 19156 14816
rect 19208 14804 19214 14816
rect 20625 14807 20683 14813
rect 20625 14804 20637 14807
rect 19208 14776 20637 14804
rect 19208 14764 19214 14776
rect 20625 14773 20637 14776
rect 20671 14773 20683 14807
rect 21082 14804 21088 14816
rect 21043 14776 21088 14804
rect 20625 14767 20683 14773
rect 21082 14764 21088 14776
rect 21140 14764 21146 14816
rect 21818 14804 21824 14816
rect 21779 14776 21824 14804
rect 21818 14764 21824 14776
rect 21876 14764 21882 14816
rect 22189 14807 22247 14813
rect 22189 14773 22201 14807
rect 22235 14804 22247 14807
rect 22922 14804 22928 14816
rect 22235 14776 22928 14804
rect 22235 14773 22247 14776
rect 22189 14767 22247 14773
rect 22922 14764 22928 14776
rect 22980 14764 22986 14816
rect 24210 14764 24216 14816
rect 24268 14804 24274 14816
rect 26988 14804 27016 14835
rect 24268 14776 27016 14804
rect 24268 14764 24274 14776
rect 1104 14714 28060 14736
rect 1104 14662 5442 14714
rect 5494 14662 5506 14714
rect 5558 14662 5570 14714
rect 5622 14662 5634 14714
rect 5686 14662 5698 14714
rect 5750 14662 14428 14714
rect 14480 14662 14492 14714
rect 14544 14662 14556 14714
rect 14608 14662 14620 14714
rect 14672 14662 14684 14714
rect 14736 14662 23413 14714
rect 23465 14662 23477 14714
rect 23529 14662 23541 14714
rect 23593 14662 23605 14714
rect 23657 14662 23669 14714
rect 23721 14662 28060 14714
rect 1104 14640 28060 14662
rect 3786 14600 3792 14612
rect 3747 14572 3792 14600
rect 3786 14560 3792 14572
rect 3844 14560 3850 14612
rect 8846 14560 8852 14612
rect 8904 14600 8910 14612
rect 8941 14603 8999 14609
rect 8941 14600 8953 14603
rect 8904 14572 8953 14600
rect 8904 14560 8910 14572
rect 8941 14569 8953 14572
rect 8987 14569 8999 14603
rect 8941 14563 8999 14569
rect 9030 14560 9036 14612
rect 9088 14600 9094 14612
rect 9088 14572 9674 14600
rect 9088 14560 9094 14572
rect 9646 14532 9674 14572
rect 9766 14560 9772 14612
rect 9824 14600 9830 14612
rect 9953 14603 10011 14609
rect 9953 14600 9965 14603
rect 9824 14572 9965 14600
rect 9824 14560 9830 14572
rect 9953 14569 9965 14572
rect 9999 14569 10011 14603
rect 11698 14600 11704 14612
rect 9953 14563 10011 14569
rect 10152 14572 11704 14600
rect 9858 14532 9864 14544
rect 9646 14504 9864 14532
rect 9858 14492 9864 14504
rect 9916 14492 9922 14544
rect 4338 14424 4344 14476
rect 4396 14464 4402 14476
rect 6457 14467 6515 14473
rect 6457 14464 6469 14467
rect 4396 14436 6469 14464
rect 4396 14424 4402 14436
rect 6457 14433 6469 14436
rect 6503 14433 6515 14467
rect 6457 14427 6515 14433
rect 8386 14424 8392 14476
rect 8444 14464 8450 14476
rect 9033 14467 9091 14473
rect 9033 14464 9045 14467
rect 8444 14436 9045 14464
rect 8444 14424 8450 14436
rect 9033 14433 9045 14436
rect 9079 14433 9091 14467
rect 9033 14427 9091 14433
rect 1397 14399 1455 14405
rect 1397 14365 1409 14399
rect 1443 14396 1455 14399
rect 2038 14396 2044 14408
rect 1443 14368 2044 14396
rect 1443 14365 1455 14368
rect 1397 14359 1455 14365
rect 2038 14356 2044 14368
rect 2096 14356 2102 14408
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14396 4031 14399
rect 4154 14396 4160 14408
rect 4019 14368 4160 14396
rect 4019 14365 4031 14368
rect 3973 14359 4031 14365
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 4246 14356 4252 14408
rect 4304 14396 4310 14408
rect 4617 14399 4675 14405
rect 4617 14396 4629 14399
rect 4304 14368 4629 14396
rect 4304 14356 4310 14368
rect 4617 14365 4629 14368
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 5261 14399 5319 14405
rect 5261 14365 5273 14399
rect 5307 14365 5319 14399
rect 5261 14359 5319 14365
rect 5997 14399 6055 14405
rect 5997 14365 6009 14399
rect 6043 14396 6055 14399
rect 6270 14396 6276 14408
rect 6043 14368 6276 14396
rect 6043 14365 6055 14368
rect 5997 14359 6055 14365
rect 1670 14337 1676 14340
rect 1664 14291 1676 14337
rect 1728 14328 1734 14340
rect 3142 14328 3148 14340
rect 1728 14300 1764 14328
rect 2792 14300 3148 14328
rect 1670 14288 1676 14291
rect 1728 14288 1734 14300
rect 2792 14269 2820 14300
rect 3142 14288 3148 14300
rect 3200 14288 3206 14340
rect 5276 14328 5304 14359
rect 6270 14356 6276 14368
rect 6328 14356 6334 14408
rect 7190 14356 7196 14408
rect 7248 14396 7254 14408
rect 7742 14396 7748 14408
rect 7248 14368 7748 14396
rect 7248 14356 7254 14368
rect 7742 14356 7748 14368
rect 7800 14356 7806 14408
rect 8662 14356 8668 14408
rect 8720 14396 8726 14408
rect 9217 14399 9275 14405
rect 9217 14396 9229 14399
rect 8720 14368 9229 14396
rect 8720 14356 8726 14368
rect 9217 14365 9229 14368
rect 9263 14365 9275 14399
rect 9217 14359 9275 14365
rect 9766 14356 9772 14408
rect 9824 14396 9830 14408
rect 10152 14405 10180 14572
rect 11698 14560 11704 14572
rect 11756 14560 11762 14612
rect 12342 14560 12348 14612
rect 12400 14600 12406 14612
rect 12621 14603 12679 14609
rect 12621 14600 12633 14603
rect 12400 14572 12633 14600
rect 12400 14560 12406 14572
rect 12621 14569 12633 14572
rect 12667 14569 12679 14603
rect 12621 14563 12679 14569
rect 13078 14560 13084 14612
rect 13136 14600 13142 14612
rect 13265 14603 13323 14609
rect 13265 14600 13277 14603
rect 13136 14572 13277 14600
rect 13136 14560 13142 14572
rect 13265 14569 13277 14572
rect 13311 14600 13323 14603
rect 15289 14603 15347 14609
rect 15289 14600 15301 14603
rect 13311 14572 15301 14600
rect 13311 14569 13323 14572
rect 13265 14563 13323 14569
rect 15289 14569 15301 14572
rect 15335 14600 15347 14603
rect 16022 14600 16028 14612
rect 15335 14572 16028 14600
rect 15335 14569 15347 14572
rect 15289 14563 15347 14569
rect 16022 14560 16028 14572
rect 16080 14560 16086 14612
rect 16117 14603 16175 14609
rect 16117 14569 16129 14603
rect 16163 14600 16175 14603
rect 16574 14600 16580 14612
rect 16163 14572 16580 14600
rect 16163 14569 16175 14572
rect 16117 14563 16175 14569
rect 16574 14560 16580 14572
rect 16632 14560 16638 14612
rect 18782 14600 18788 14612
rect 17696 14572 18788 14600
rect 11146 14532 11152 14544
rect 10428 14504 11152 14532
rect 10428 14473 10456 14504
rect 11146 14492 11152 14504
rect 11204 14492 11210 14544
rect 11793 14535 11851 14541
rect 11793 14501 11805 14535
rect 11839 14532 11851 14535
rect 14553 14535 14611 14541
rect 11839 14504 14520 14532
rect 11839 14501 11851 14504
rect 11793 14495 11851 14501
rect 10413 14467 10471 14473
rect 10413 14433 10425 14467
rect 10459 14433 10471 14467
rect 10413 14427 10471 14433
rect 10686 14424 10692 14476
rect 10744 14464 10750 14476
rect 10962 14464 10968 14476
rect 10744 14436 10968 14464
rect 10744 14424 10750 14436
rect 10962 14424 10968 14436
rect 11020 14424 11026 14476
rect 11057 14467 11115 14473
rect 11057 14433 11069 14467
rect 11103 14464 11115 14467
rect 12158 14464 12164 14476
rect 11103 14436 12164 14464
rect 11103 14433 11115 14436
rect 11057 14427 11115 14433
rect 12158 14424 12164 14436
rect 12216 14424 12222 14476
rect 13906 14424 13912 14476
rect 13964 14464 13970 14476
rect 14492 14464 14520 14504
rect 14553 14501 14565 14535
rect 14599 14532 14611 14535
rect 14599 14504 14872 14532
rect 14599 14501 14611 14504
rect 14553 14495 14611 14501
rect 14844 14476 14872 14504
rect 15010 14492 15016 14544
rect 15068 14532 15074 14544
rect 17586 14532 17592 14544
rect 15068 14504 17592 14532
rect 15068 14492 15074 14504
rect 17586 14492 17592 14504
rect 17644 14492 17650 14544
rect 13964 14436 14428 14464
rect 14492 14436 14780 14464
rect 13964 14424 13970 14436
rect 10137 14399 10195 14405
rect 10137 14396 10149 14399
rect 9824 14368 10149 14396
rect 9824 14356 9830 14368
rect 10137 14365 10149 14368
rect 10183 14365 10195 14399
rect 10318 14396 10324 14408
rect 10279 14368 10324 14396
rect 10137 14359 10195 14365
rect 10318 14356 10324 14368
rect 10376 14356 10382 14408
rect 10594 14356 10600 14408
rect 10652 14396 10658 14408
rect 11241 14399 11299 14405
rect 11241 14396 11253 14399
rect 10652 14368 11253 14396
rect 10652 14356 10658 14368
rect 11241 14365 11253 14368
rect 11287 14365 11299 14399
rect 11241 14359 11299 14365
rect 11514 14356 11520 14408
rect 11572 14396 11578 14408
rect 14400 14405 14428 14436
rect 11701 14399 11759 14405
rect 11701 14396 11713 14399
rect 11572 14368 11713 14396
rect 11572 14356 11578 14368
rect 11701 14365 11713 14368
rect 11747 14365 11759 14399
rect 13449 14399 13507 14405
rect 13449 14396 13461 14399
rect 11701 14359 11759 14365
rect 11808 14368 13461 14396
rect 6454 14328 6460 14340
rect 5276 14300 6460 14328
rect 6454 14288 6460 14300
rect 6512 14288 6518 14340
rect 6730 14337 6736 14340
rect 6724 14291 6736 14337
rect 6788 14328 6794 14340
rect 8941 14331 8999 14337
rect 6788 14300 6824 14328
rect 6730 14288 6736 14291
rect 6788 14288 6794 14300
rect 8941 14297 8953 14331
rect 8987 14328 8999 14331
rect 9490 14328 9496 14340
rect 8987 14300 9496 14328
rect 8987 14297 8999 14300
rect 8941 14291 8999 14297
rect 9490 14288 9496 14300
rect 9548 14288 9554 14340
rect 11330 14288 11336 14340
rect 11388 14328 11394 14340
rect 11808 14328 11836 14368
rect 13449 14365 13461 14368
rect 13495 14365 13507 14399
rect 13449 14359 13507 14365
rect 14278 14399 14336 14405
rect 14278 14365 14290 14399
rect 14324 14365 14336 14399
rect 14278 14359 14336 14365
rect 14370 14399 14428 14405
rect 14370 14365 14382 14399
rect 14416 14365 14428 14399
rect 14370 14359 14428 14365
rect 11388 14300 11836 14328
rect 11388 14288 11394 14300
rect 11882 14288 11888 14340
rect 11940 14328 11946 14340
rect 12437 14331 12495 14337
rect 12437 14328 12449 14331
rect 11940 14300 12449 14328
rect 11940 14288 11946 14300
rect 12437 14297 12449 14300
rect 12483 14297 12495 14331
rect 12437 14291 12495 14297
rect 12618 14288 12624 14340
rect 12676 14337 12682 14340
rect 12676 14331 12695 14337
rect 12683 14297 12695 14331
rect 12676 14291 12695 14297
rect 12676 14288 12682 14291
rect 13170 14288 13176 14340
rect 13228 14328 13234 14340
rect 14093 14331 14151 14337
rect 14093 14328 14105 14331
rect 13228 14300 14105 14328
rect 13228 14288 13234 14300
rect 14093 14297 14105 14300
rect 14139 14297 14151 14331
rect 14292 14328 14320 14359
rect 14458 14356 14464 14408
rect 14516 14396 14522 14408
rect 14599 14399 14657 14405
rect 14599 14396 14611 14399
rect 14516 14368 14611 14396
rect 14516 14356 14522 14368
rect 14599 14365 14611 14368
rect 14645 14365 14657 14399
rect 14752 14396 14780 14436
rect 14826 14424 14832 14476
rect 14884 14424 14890 14476
rect 17696 14464 17724 14572
rect 18782 14560 18788 14572
rect 18840 14600 18846 14612
rect 19886 14600 19892 14612
rect 18840 14572 19892 14600
rect 18840 14560 18846 14572
rect 19886 14560 19892 14572
rect 19944 14560 19950 14612
rect 21542 14600 21548 14612
rect 20088 14572 21548 14600
rect 17862 14492 17868 14544
rect 17920 14532 17926 14544
rect 18046 14532 18052 14544
rect 17920 14504 18052 14532
rect 17920 14492 17926 14504
rect 18046 14492 18052 14504
rect 18104 14532 18110 14544
rect 19610 14532 19616 14544
rect 18104 14504 19616 14532
rect 18104 14492 18110 14504
rect 19610 14492 19616 14504
rect 19668 14492 19674 14544
rect 19334 14464 19340 14476
rect 15796 14436 17724 14464
rect 17972 14436 19340 14464
rect 15796 14396 15824 14436
rect 15930 14396 15936 14408
rect 14752 14368 15824 14396
rect 15891 14368 15936 14396
rect 14599 14359 14657 14365
rect 15930 14356 15936 14368
rect 15988 14356 15994 14408
rect 16022 14356 16028 14408
rect 16080 14396 16086 14408
rect 17218 14396 17224 14408
rect 16080 14368 17224 14396
rect 16080 14356 16086 14368
rect 17218 14356 17224 14368
rect 17276 14356 17282 14408
rect 17862 14396 17868 14408
rect 17823 14368 17868 14396
rect 17862 14356 17868 14368
rect 17920 14356 17926 14408
rect 15010 14328 15016 14340
rect 14292 14300 15016 14328
rect 14093 14291 14151 14297
rect 15010 14288 15016 14300
rect 15068 14288 15074 14340
rect 15105 14331 15163 14337
rect 15105 14297 15117 14331
rect 15151 14328 15163 14331
rect 15194 14328 15200 14340
rect 15151 14300 15200 14328
rect 15151 14297 15163 14300
rect 15105 14291 15163 14297
rect 15194 14288 15200 14300
rect 15252 14288 15258 14340
rect 15305 14331 15363 14337
rect 15305 14297 15317 14331
rect 15351 14328 15363 14331
rect 15838 14328 15844 14340
rect 15351 14300 15844 14328
rect 15351 14297 15363 14300
rect 15305 14291 15363 14297
rect 15838 14288 15844 14300
rect 15896 14288 15902 14340
rect 16666 14288 16672 14340
rect 16724 14328 16730 14340
rect 16761 14331 16819 14337
rect 16761 14328 16773 14331
rect 16724 14300 16773 14328
rect 16724 14288 16730 14300
rect 16761 14297 16773 14300
rect 16807 14328 16819 14331
rect 17972 14328 18000 14436
rect 19334 14424 19340 14436
rect 19392 14464 19398 14476
rect 19518 14464 19524 14476
rect 19392 14436 19524 14464
rect 19392 14424 19398 14436
rect 19518 14424 19524 14436
rect 19576 14424 19582 14476
rect 18049 14399 18107 14405
rect 18049 14365 18061 14399
rect 18095 14396 18107 14399
rect 18690 14396 18696 14408
rect 18095 14368 18696 14396
rect 18095 14365 18107 14368
rect 18049 14359 18107 14365
rect 18690 14356 18696 14368
rect 18748 14356 18754 14408
rect 18782 14356 18788 14408
rect 18840 14396 18846 14408
rect 18840 14368 19564 14396
rect 18840 14356 18846 14368
rect 16807 14300 18000 14328
rect 18708 14328 18736 14356
rect 19150 14328 19156 14340
rect 18708 14300 19156 14328
rect 16807 14297 16819 14300
rect 16761 14291 16819 14297
rect 19150 14288 19156 14300
rect 19208 14288 19214 14340
rect 19334 14328 19340 14340
rect 19295 14300 19340 14328
rect 19334 14288 19340 14300
rect 19392 14288 19398 14340
rect 2777 14263 2835 14269
rect 2777 14229 2789 14263
rect 2823 14229 2835 14263
rect 2777 14223 2835 14229
rect 2866 14220 2872 14272
rect 2924 14260 2930 14272
rect 4433 14263 4491 14269
rect 4433 14260 4445 14263
rect 2924 14232 4445 14260
rect 2924 14220 2930 14232
rect 4433 14229 4445 14232
rect 4479 14229 4491 14263
rect 5074 14260 5080 14272
rect 5035 14232 5080 14260
rect 4433 14223 4491 14229
rect 5074 14220 5080 14232
rect 5132 14220 5138 14272
rect 5810 14260 5816 14272
rect 5771 14232 5816 14260
rect 5810 14220 5816 14232
rect 5868 14220 5874 14272
rect 7006 14220 7012 14272
rect 7064 14260 7070 14272
rect 7837 14263 7895 14269
rect 7837 14260 7849 14263
rect 7064 14232 7849 14260
rect 7064 14220 7070 14232
rect 7837 14229 7849 14232
rect 7883 14260 7895 14263
rect 8202 14260 8208 14272
rect 7883 14232 8208 14260
rect 7883 14229 7895 14232
rect 7837 14223 7895 14229
rect 8202 14220 8208 14232
rect 8260 14220 8266 14272
rect 9401 14263 9459 14269
rect 9401 14229 9413 14263
rect 9447 14260 9459 14263
rect 10594 14260 10600 14272
rect 9447 14232 10600 14260
rect 9447 14229 9459 14232
rect 9401 14223 9459 14229
rect 10594 14220 10600 14232
rect 10652 14220 10658 14272
rect 12805 14263 12863 14269
rect 12805 14229 12817 14263
rect 12851 14260 12863 14263
rect 13262 14260 13268 14272
rect 12851 14232 13268 14260
rect 12851 14229 12863 14232
rect 12805 14223 12863 14229
rect 13262 14220 13268 14232
rect 13320 14220 13326 14272
rect 15470 14260 15476 14272
rect 15431 14232 15476 14260
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 16853 14263 16911 14269
rect 16853 14229 16865 14263
rect 16899 14260 16911 14263
rect 17770 14260 17776 14272
rect 16899 14232 17776 14260
rect 16899 14229 16911 14232
rect 16853 14223 16911 14229
rect 17770 14220 17776 14232
rect 17828 14220 17834 14272
rect 18233 14263 18291 14269
rect 18233 14229 18245 14263
rect 18279 14260 18291 14263
rect 18414 14260 18420 14272
rect 18279 14232 18420 14260
rect 18279 14229 18291 14232
rect 18233 14223 18291 14229
rect 18414 14220 18420 14232
rect 18472 14220 18478 14272
rect 18506 14220 18512 14272
rect 18564 14260 18570 14272
rect 19429 14263 19487 14269
rect 19429 14260 19441 14263
rect 18564 14232 19441 14260
rect 18564 14220 18570 14232
rect 19429 14229 19441 14232
rect 19475 14229 19487 14263
rect 19536 14260 19564 14368
rect 20088 14328 20116 14572
rect 21542 14560 21548 14572
rect 21600 14560 21606 14612
rect 22278 14600 22284 14612
rect 22239 14572 22284 14600
rect 22278 14560 22284 14572
rect 22336 14560 22342 14612
rect 23106 14560 23112 14612
rect 23164 14600 23170 14612
rect 27341 14603 27399 14609
rect 27341 14600 27353 14603
rect 23164 14572 27353 14600
rect 23164 14560 23170 14572
rect 27341 14569 27353 14572
rect 27387 14569 27399 14603
rect 27341 14563 27399 14569
rect 21818 14492 21824 14544
rect 21876 14532 21882 14544
rect 21876 14504 24808 14532
rect 21876 14492 21882 14504
rect 21542 14424 21548 14476
rect 21600 14464 21606 14476
rect 22925 14467 22983 14473
rect 22925 14464 22937 14467
rect 21600 14436 22937 14464
rect 21600 14424 21606 14436
rect 22925 14433 22937 14436
rect 22971 14464 22983 14467
rect 23290 14464 23296 14476
rect 22971 14436 23296 14464
rect 22971 14433 22983 14436
rect 22925 14427 22983 14433
rect 23290 14424 23296 14436
rect 23348 14424 23354 14476
rect 23750 14424 23756 14476
rect 23808 14464 23814 14476
rect 24397 14467 24455 14473
rect 24397 14464 24409 14467
rect 23808 14436 24409 14464
rect 23808 14424 23814 14436
rect 24397 14433 24409 14436
rect 24443 14433 24455 14467
rect 24397 14427 24455 14433
rect 20165 14399 20223 14405
rect 20165 14365 20177 14399
rect 20211 14396 20223 14399
rect 21910 14396 21916 14408
rect 20211 14368 21916 14396
rect 20211 14365 20223 14368
rect 20165 14359 20223 14365
rect 21910 14356 21916 14368
rect 21968 14356 21974 14408
rect 24210 14396 24216 14408
rect 22066 14368 24216 14396
rect 20410 14331 20468 14337
rect 20410 14328 20422 14331
rect 20088 14300 20422 14328
rect 20410 14297 20422 14300
rect 20456 14297 20468 14331
rect 22066 14328 22094 14368
rect 24210 14356 24216 14368
rect 24268 14356 24274 14408
rect 24673 14399 24731 14405
rect 24673 14365 24685 14399
rect 24719 14365 24731 14399
rect 24780 14396 24808 14504
rect 25958 14464 25964 14476
rect 25919 14436 25964 14464
rect 25958 14424 25964 14436
rect 26016 14424 26022 14476
rect 26217 14399 26275 14405
rect 26217 14396 26229 14399
rect 24780 14368 26229 14396
rect 24673 14359 24731 14365
rect 26217 14365 26229 14368
rect 26263 14365 26275 14399
rect 26217 14359 26275 14365
rect 20410 14291 20468 14297
rect 20548 14300 22094 14328
rect 20548 14260 20576 14300
rect 22278 14288 22284 14340
rect 22336 14328 22342 14340
rect 22649 14331 22707 14337
rect 22649 14328 22661 14331
rect 22336 14300 22661 14328
rect 22336 14288 22342 14300
rect 22649 14297 22661 14300
rect 22695 14297 22707 14331
rect 23658 14328 23664 14340
rect 23619 14300 23664 14328
rect 22649 14291 22707 14297
rect 23658 14288 23664 14300
rect 23716 14288 23722 14340
rect 23845 14331 23903 14337
rect 23845 14297 23857 14331
rect 23891 14328 23903 14331
rect 24302 14328 24308 14340
rect 23891 14300 24308 14328
rect 23891 14297 23903 14300
rect 23845 14291 23903 14297
rect 21542 14260 21548 14272
rect 19536 14232 20576 14260
rect 21503 14232 21548 14260
rect 19429 14223 19487 14229
rect 21542 14220 21548 14232
rect 21600 14220 21606 14272
rect 22094 14220 22100 14272
rect 22152 14260 22158 14272
rect 22741 14263 22799 14269
rect 22741 14260 22753 14263
rect 22152 14232 22753 14260
rect 22152 14220 22158 14232
rect 22741 14229 22753 14232
rect 22787 14229 22799 14263
rect 22741 14223 22799 14229
rect 22922 14220 22928 14272
rect 22980 14260 22986 14272
rect 23860 14260 23888 14291
rect 24302 14288 24308 14300
rect 24360 14288 24366 14340
rect 24688 14328 24716 14359
rect 25866 14328 25872 14340
rect 24688 14300 25872 14328
rect 22980 14232 23888 14260
rect 22980 14220 22986 14232
rect 24210 14220 24216 14272
rect 24268 14260 24274 14272
rect 24688 14260 24716 14300
rect 25866 14288 25872 14300
rect 25924 14288 25930 14340
rect 24268 14232 24716 14260
rect 24268 14220 24274 14232
rect 1104 14170 28060 14192
rect 1104 14118 9935 14170
rect 9987 14118 9999 14170
rect 10051 14118 10063 14170
rect 10115 14118 10127 14170
rect 10179 14118 10191 14170
rect 10243 14118 18920 14170
rect 18972 14118 18984 14170
rect 19036 14118 19048 14170
rect 19100 14118 19112 14170
rect 19164 14118 19176 14170
rect 19228 14118 28060 14170
rect 1104 14096 28060 14118
rect 1670 14056 1676 14068
rect 1631 14028 1676 14056
rect 1670 14016 1676 14028
rect 1728 14016 1734 14068
rect 3142 14016 3148 14068
rect 3200 14056 3206 14068
rect 3970 14056 3976 14068
rect 3200 14028 3976 14056
rect 3200 14016 3206 14028
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 6730 14056 6736 14068
rect 6691 14028 6736 14056
rect 6730 14016 6736 14028
rect 6788 14016 6794 14068
rect 8662 14016 8668 14068
rect 8720 14056 8726 14068
rect 9217 14059 9275 14065
rect 8720 14028 8892 14056
rect 8720 14016 8726 14028
rect 4338 13988 4344 14000
rect 2608 13960 4344 13988
rect 1854 13920 1860 13932
rect 1815 13892 1860 13920
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 2608 13929 2636 13960
rect 4338 13948 4344 13960
rect 4396 13948 4402 14000
rect 4700 13991 4758 13997
rect 4700 13957 4712 13991
rect 4746 13988 4758 13991
rect 5810 13988 5816 14000
rect 4746 13960 5816 13988
rect 4746 13957 4758 13960
rect 4700 13951 4758 13957
rect 5810 13948 5816 13960
rect 5868 13948 5874 14000
rect 7929 13991 7987 13997
rect 7929 13957 7941 13991
rect 7975 13988 7987 13991
rect 8294 13988 8300 14000
rect 7975 13960 8300 13988
rect 7975 13957 7987 13960
rect 7929 13951 7987 13957
rect 8294 13948 8300 13960
rect 8352 13948 8358 14000
rect 8478 13948 8484 14000
rect 8536 13988 8542 14000
rect 8573 13991 8631 13997
rect 8573 13988 8585 13991
rect 8536 13960 8585 13988
rect 8536 13948 8542 13960
rect 8573 13957 8585 13960
rect 8619 13957 8631 13991
rect 8573 13951 8631 13957
rect 2866 13929 2872 13932
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13889 2651 13923
rect 2593 13883 2651 13889
rect 2860 13883 2872 13929
rect 2924 13920 2930 13932
rect 6917 13923 6975 13929
rect 2924 13892 2960 13920
rect 1670 13812 1676 13864
rect 1728 13852 1734 13864
rect 2038 13852 2044 13864
rect 1728 13824 2044 13852
rect 1728 13812 1734 13824
rect 2038 13812 2044 13824
rect 2096 13852 2102 13864
rect 2608 13852 2636 13883
rect 2866 13880 2872 13883
rect 2924 13880 2930 13892
rect 6917 13889 6929 13923
rect 6963 13920 6975 13923
rect 7742 13920 7748 13932
rect 6963 13892 7748 13920
rect 6963 13889 6975 13892
rect 6917 13883 6975 13889
rect 7742 13880 7748 13892
rect 7800 13880 7806 13932
rect 8386 13880 8392 13932
rect 8444 13920 8450 13932
rect 8720 13923 8778 13929
rect 8720 13920 8732 13923
rect 8444 13892 8732 13920
rect 8444 13880 8450 13892
rect 8720 13889 8732 13892
rect 8766 13889 8778 13923
rect 8720 13883 8778 13889
rect 2096 13824 2636 13852
rect 2096 13812 2102 13824
rect 4338 13812 4344 13864
rect 4396 13852 4402 13864
rect 4433 13855 4491 13861
rect 4433 13852 4445 13855
rect 4396 13824 4445 13852
rect 4396 13812 4402 13824
rect 4433 13821 4445 13824
rect 4479 13821 4491 13855
rect 8864 13852 8892 14028
rect 9217 14025 9229 14059
rect 9263 14056 9275 14059
rect 10686 14056 10692 14068
rect 9263 14028 10692 14056
rect 9263 14025 9275 14028
rect 9217 14019 9275 14025
rect 10686 14016 10692 14028
rect 10744 14016 10750 14068
rect 10778 14016 10784 14068
rect 10836 14056 10842 14068
rect 10836 14028 10881 14056
rect 10836 14016 10842 14028
rect 11514 14016 11520 14068
rect 11572 14056 11578 14068
rect 12371 14059 12429 14065
rect 11572 14028 12204 14056
rect 11572 14016 11578 14028
rect 12176 13997 12204 14028
rect 12371 14025 12383 14059
rect 12417 14056 12429 14059
rect 12618 14056 12624 14068
rect 12417 14028 12624 14056
rect 12417 14025 12429 14028
rect 12371 14019 12429 14025
rect 12618 14016 12624 14028
rect 12676 14016 12682 14068
rect 12710 14016 12716 14068
rect 12768 14056 12774 14068
rect 12894 14056 12900 14068
rect 12768 14028 12900 14056
rect 12768 14016 12774 14028
rect 12894 14016 12900 14028
rect 12952 14016 12958 14068
rect 14458 14056 14464 14068
rect 14419 14028 14464 14056
rect 14458 14016 14464 14028
rect 14516 14016 14522 14068
rect 15010 14016 15016 14068
rect 15068 14056 15074 14068
rect 15121 14059 15179 14065
rect 15121 14056 15133 14059
rect 15068 14028 15133 14056
rect 15068 14016 15074 14028
rect 15121 14025 15133 14028
rect 15167 14025 15179 14059
rect 15286 14056 15292 14068
rect 15247 14028 15292 14056
rect 15121 14019 15179 14025
rect 15286 14016 15292 14028
rect 15344 14016 15350 14068
rect 15470 14016 15476 14068
rect 15528 14056 15534 14068
rect 18506 14056 18512 14068
rect 15528 14028 18512 14056
rect 15528 14016 15534 14028
rect 18506 14016 18512 14028
rect 18564 14016 18570 14068
rect 18782 14056 18788 14068
rect 18607 14028 18788 14056
rect 12161 13991 12219 13997
rect 12161 13957 12173 13991
rect 12207 13957 12219 13991
rect 12161 13951 12219 13957
rect 13538 13948 13544 14000
rect 13596 13948 13602 14000
rect 14642 13948 14648 14000
rect 14700 13988 14706 14000
rect 14921 13991 14979 13997
rect 14921 13988 14933 13991
rect 14700 13960 14933 13988
rect 14700 13948 14706 13960
rect 14921 13957 14933 13960
rect 14967 13988 14979 13991
rect 15654 13988 15660 14000
rect 14967 13960 15660 13988
rect 14967 13957 14979 13960
rect 14921 13951 14979 13957
rect 15654 13948 15660 13960
rect 15712 13988 15718 14000
rect 15749 13991 15807 13997
rect 15749 13988 15761 13991
rect 15712 13960 15761 13988
rect 15712 13948 15718 13960
rect 15749 13957 15761 13960
rect 15795 13957 15807 13991
rect 15749 13951 15807 13957
rect 15965 13991 16023 13997
rect 15965 13957 15977 13991
rect 16011 13988 16023 13991
rect 16574 13988 16580 14000
rect 16011 13960 16580 13988
rect 16011 13957 16023 13960
rect 15965 13951 16023 13957
rect 16574 13948 16580 13960
rect 16632 13948 16638 14000
rect 16936 13991 16994 13997
rect 16936 13957 16948 13991
rect 16982 13988 16994 13991
rect 18607 13988 18635 14028
rect 18782 14016 18788 14028
rect 18840 14016 18846 14068
rect 19153 14059 19211 14065
rect 19153 14025 19165 14059
rect 19199 14056 19211 14059
rect 19242 14056 19248 14068
rect 19199 14028 19248 14056
rect 19199 14025 19211 14028
rect 19153 14019 19211 14025
rect 19242 14016 19248 14028
rect 19300 14016 19306 14068
rect 20714 14016 20720 14068
rect 20772 14056 20778 14068
rect 22005 14059 22063 14065
rect 22005 14056 22017 14059
rect 20772 14028 20944 14056
rect 20772 14016 20778 14028
rect 19518 13988 19524 14000
rect 16982 13960 18635 13988
rect 18708 13960 19524 13988
rect 16982 13957 16994 13960
rect 16936 13951 16994 13957
rect 9769 13923 9827 13929
rect 9769 13889 9781 13923
rect 9815 13920 9827 13923
rect 10505 13923 10563 13929
rect 9815 13892 10468 13920
rect 9815 13889 9827 13892
rect 9769 13883 9827 13889
rect 8941 13855 8999 13861
rect 8941 13852 8953 13855
rect 8864 13824 8953 13852
rect 4433 13815 4491 13821
rect 8941 13821 8953 13824
rect 8987 13821 8999 13855
rect 10045 13855 10103 13861
rect 10045 13852 10057 13855
rect 8941 13815 8999 13821
rect 9784 13824 10057 13852
rect 9784 13796 9812 13824
rect 10045 13821 10057 13824
rect 10091 13821 10103 13855
rect 10440 13852 10468 13892
rect 10505 13889 10517 13923
rect 10551 13920 10563 13923
rect 10686 13920 10692 13932
rect 10551 13892 10692 13920
rect 10551 13889 10563 13892
rect 10505 13883 10563 13889
rect 10686 13880 10692 13892
rect 10744 13920 10750 13932
rect 11422 13920 11428 13932
rect 10744 13892 11428 13920
rect 10744 13880 10750 13892
rect 11422 13880 11428 13892
rect 11480 13880 11486 13932
rect 11514 13880 11520 13932
rect 11572 13920 11578 13932
rect 13348 13923 13406 13929
rect 11572 13892 11617 13920
rect 11572 13880 11578 13892
rect 13348 13889 13360 13923
rect 13394 13920 13406 13923
rect 13556 13920 13584 13948
rect 18414 13920 18420 13932
rect 13394 13892 13584 13920
rect 14573 13892 18420 13920
rect 13394 13889 13406 13892
rect 13348 13883 13406 13889
rect 10781 13855 10839 13861
rect 10781 13852 10793 13855
rect 10440 13824 10793 13852
rect 10045 13815 10103 13821
rect 10781 13821 10793 13824
rect 10827 13852 10839 13855
rect 11146 13852 11152 13864
rect 10827 13824 11152 13852
rect 10827 13821 10839 13824
rect 10781 13815 10839 13821
rect 11146 13812 11152 13824
rect 11204 13812 11210 13864
rect 11606 13852 11612 13864
rect 11567 13824 11612 13852
rect 11606 13812 11612 13824
rect 11664 13812 11670 13864
rect 11698 13812 11704 13864
rect 11756 13852 11762 13864
rect 13081 13855 13139 13861
rect 13081 13852 13093 13855
rect 11756 13824 13093 13852
rect 11756 13812 11762 13824
rect 13081 13821 13093 13824
rect 13127 13821 13139 13855
rect 13081 13815 13139 13821
rect 8113 13787 8171 13793
rect 8113 13753 8125 13787
rect 8159 13784 8171 13787
rect 8202 13784 8208 13796
rect 8159 13756 8208 13784
rect 8159 13753 8171 13756
rect 8113 13747 8171 13753
rect 8202 13744 8208 13756
rect 8260 13744 8266 13796
rect 9766 13744 9772 13796
rect 9824 13744 9830 13796
rect 9861 13787 9919 13793
rect 9861 13753 9873 13787
rect 9907 13784 9919 13787
rect 10318 13784 10324 13796
rect 9907 13756 10324 13784
rect 9907 13753 9919 13756
rect 9861 13747 9919 13753
rect 10318 13744 10324 13756
rect 10376 13744 10382 13796
rect 10594 13784 10600 13796
rect 10555 13756 10600 13784
rect 10594 13744 10600 13756
rect 10652 13744 10658 13796
rect 2866 13676 2872 13728
rect 2924 13716 2930 13728
rect 3234 13716 3240 13728
rect 2924 13688 3240 13716
rect 2924 13676 2930 13688
rect 3234 13676 3240 13688
rect 3292 13676 3298 13728
rect 3973 13719 4031 13725
rect 3973 13685 3985 13719
rect 4019 13716 4031 13719
rect 4154 13716 4160 13728
rect 4019 13688 4160 13716
rect 4019 13685 4031 13688
rect 3973 13679 4031 13685
rect 4154 13676 4160 13688
rect 4212 13716 4218 13728
rect 5166 13716 5172 13728
rect 4212 13688 5172 13716
rect 4212 13676 4218 13688
rect 5166 13676 5172 13688
rect 5224 13676 5230 13728
rect 5350 13676 5356 13728
rect 5408 13716 5414 13728
rect 5813 13719 5871 13725
rect 5813 13716 5825 13719
rect 5408 13688 5825 13716
rect 5408 13676 5414 13688
rect 5813 13685 5825 13688
rect 5859 13685 5871 13719
rect 8846 13716 8852 13728
rect 8807 13688 8852 13716
rect 5813 13679 5871 13685
rect 8846 13676 8852 13688
rect 8904 13676 8910 13728
rect 9950 13716 9956 13728
rect 9911 13688 9956 13716
rect 9950 13676 9956 13688
rect 10008 13676 10014 13728
rect 10410 13676 10416 13728
rect 10468 13716 10474 13728
rect 11146 13716 11152 13728
rect 10468 13688 11152 13716
rect 10468 13676 10474 13688
rect 11146 13676 11152 13688
rect 11204 13676 11210 13728
rect 12342 13716 12348 13728
rect 12303 13688 12348 13716
rect 12342 13676 12348 13688
rect 12400 13676 12406 13728
rect 12529 13719 12587 13725
rect 12529 13685 12541 13719
rect 12575 13716 12587 13719
rect 14573 13716 14601 13892
rect 18414 13880 18420 13892
rect 18472 13880 18478 13932
rect 18506 13880 18512 13932
rect 18564 13920 18570 13932
rect 18708 13929 18736 13960
rect 19518 13948 19524 13960
rect 19576 13948 19582 14000
rect 19886 13988 19892 14000
rect 19847 13960 19892 13988
rect 19886 13948 19892 13960
rect 19944 13948 19950 14000
rect 20916 13997 20944 14028
rect 21744 14028 22017 14056
rect 20901 13991 20959 13997
rect 20901 13957 20913 13991
rect 20947 13957 20959 13991
rect 20901 13951 20959 13957
rect 20993 13991 21051 13997
rect 20993 13957 21005 13991
rect 21039 13988 21051 13991
rect 21542 13988 21548 14000
rect 21039 13960 21548 13988
rect 21039 13957 21051 13960
rect 20993 13951 21051 13957
rect 21542 13948 21548 13960
rect 21600 13948 21606 14000
rect 18657 13923 18736 13929
rect 18564 13892 18609 13920
rect 18564 13880 18570 13892
rect 18657 13889 18669 13923
rect 18703 13892 18736 13923
rect 18785 13923 18843 13929
rect 18703 13889 18715 13892
rect 18657 13883 18715 13889
rect 18785 13889 18797 13923
rect 18831 13889 18843 13923
rect 18785 13883 18843 13889
rect 16390 13852 16396 13864
rect 16132 13824 16396 13852
rect 14734 13744 14740 13796
rect 14792 13784 14798 13796
rect 16132 13793 16160 13824
rect 16390 13812 16396 13824
rect 16448 13812 16454 13864
rect 16666 13852 16672 13864
rect 16627 13824 16672 13852
rect 16666 13812 16672 13824
rect 16724 13812 16730 13864
rect 16117 13787 16175 13793
rect 14792 13756 16084 13784
rect 14792 13744 14798 13756
rect 12575 13688 14601 13716
rect 15105 13719 15163 13725
rect 12575 13685 12587 13688
rect 12529 13679 12587 13685
rect 15105 13685 15117 13719
rect 15151 13716 15163 13719
rect 15286 13716 15292 13728
rect 15151 13688 15292 13716
rect 15151 13685 15163 13688
rect 15105 13679 15163 13685
rect 15286 13676 15292 13688
rect 15344 13716 15350 13728
rect 15838 13716 15844 13728
rect 15344 13688 15844 13716
rect 15344 13676 15350 13688
rect 15838 13676 15844 13688
rect 15896 13716 15902 13728
rect 15933 13719 15991 13725
rect 15933 13716 15945 13719
rect 15896 13688 15945 13716
rect 15896 13676 15902 13688
rect 15933 13685 15945 13688
rect 15979 13685 15991 13719
rect 16056 13716 16084 13756
rect 16117 13753 16129 13787
rect 16163 13753 16175 13787
rect 16117 13747 16175 13753
rect 17862 13744 17868 13796
rect 17920 13784 17926 13796
rect 17920 13756 18635 13784
rect 17920 13744 17926 13756
rect 17770 13716 17776 13728
rect 16056 13688 17776 13716
rect 15933 13679 15991 13685
rect 17770 13676 17776 13688
rect 17828 13676 17834 13728
rect 17954 13676 17960 13728
rect 18012 13716 18018 13728
rect 18049 13719 18107 13725
rect 18049 13716 18061 13719
rect 18012 13688 18061 13716
rect 18012 13676 18018 13688
rect 18049 13685 18061 13688
rect 18095 13685 18107 13719
rect 18607 13716 18635 13756
rect 18800 13716 18828 13883
rect 18874 13880 18880 13932
rect 18932 13920 18938 13932
rect 19058 13929 19064 13932
rect 19015 13923 19064 13929
rect 18932 13892 18977 13920
rect 18932 13880 18938 13892
rect 19015 13889 19027 13923
rect 19061 13889 19064 13923
rect 19015 13883 19064 13889
rect 19058 13880 19064 13883
rect 19116 13880 19122 13932
rect 19610 13880 19616 13932
rect 19668 13920 19674 13932
rect 21174 13929 21180 13932
rect 19705 13923 19763 13929
rect 19705 13920 19717 13923
rect 19668 13892 19717 13920
rect 19668 13880 19674 13892
rect 19705 13889 19717 13892
rect 19751 13889 19763 13923
rect 20614 13923 20672 13929
rect 20614 13920 20626 13923
rect 19705 13883 19763 13889
rect 20548 13892 20626 13920
rect 19150 13812 19156 13864
rect 19208 13852 19214 13864
rect 20548 13852 20576 13892
rect 20614 13889 20626 13892
rect 20660 13889 20672 13923
rect 20614 13883 20672 13889
rect 20718 13923 20776 13929
rect 20718 13889 20730 13923
rect 20764 13889 20776 13923
rect 20718 13883 20776 13889
rect 21131 13923 21180 13929
rect 21131 13889 21143 13923
rect 21177 13889 21180 13923
rect 21131 13883 21180 13889
rect 19208 13824 20576 13852
rect 19208 13812 19214 13824
rect 20073 13787 20131 13793
rect 20073 13753 20085 13787
rect 20119 13784 20131 13787
rect 20346 13784 20352 13796
rect 20119 13756 20352 13784
rect 20119 13753 20131 13756
rect 20073 13747 20131 13753
rect 20346 13744 20352 13756
rect 20404 13744 20410 13796
rect 20622 13744 20628 13796
rect 20680 13784 20686 13796
rect 20733 13784 20761 13883
rect 21174 13880 21180 13883
rect 21232 13880 21238 13932
rect 21744 13796 21772 14028
rect 22005 14025 22017 14028
rect 22051 14025 22063 14059
rect 25130 14056 25136 14068
rect 22005 14019 22063 14025
rect 24044 14028 25136 14056
rect 22572 13960 23796 13988
rect 21818 13880 21824 13932
rect 21876 13920 21882 13932
rect 22572 13929 22600 13960
rect 22557 13923 22615 13929
rect 22557 13920 22569 13923
rect 21876 13892 21921 13920
rect 22020 13892 22569 13920
rect 21876 13880 21882 13892
rect 21910 13812 21916 13864
rect 21968 13852 21974 13864
rect 22020 13852 22048 13892
rect 22557 13889 22569 13892
rect 22603 13889 22615 13923
rect 22557 13883 22615 13889
rect 22646 13880 22652 13932
rect 22704 13920 22710 13932
rect 22741 13923 22799 13929
rect 22741 13920 22753 13923
rect 22704 13892 22753 13920
rect 22704 13880 22710 13892
rect 22741 13889 22753 13892
rect 22787 13889 22799 13923
rect 23106 13920 23112 13932
rect 23067 13892 23112 13920
rect 22741 13883 22799 13889
rect 23106 13880 23112 13892
rect 23164 13880 23170 13932
rect 23198 13880 23204 13932
rect 23256 13920 23262 13932
rect 23768 13929 23796 13960
rect 24044 13944 24072 14028
rect 25130 14016 25136 14028
rect 25188 14016 25194 14068
rect 26237 14059 26295 14065
rect 26237 14025 26249 14059
rect 26283 14056 26295 14059
rect 26786 14056 26792 14068
rect 26283 14028 26792 14056
rect 26283 14025 26295 14028
rect 26237 14019 26295 14025
rect 26786 14016 26792 14028
rect 26844 14016 26850 14068
rect 26973 14059 27031 14065
rect 26973 14025 26985 14059
rect 27019 14025 27031 14059
rect 26973 14019 27031 14025
rect 24210 13988 24216 14000
rect 23952 13942 24072 13944
rect 23943 13935 24072 13942
rect 23925 13929 24072 13935
rect 24136 13960 24216 13988
rect 24136 13929 24164 13960
rect 24210 13948 24216 13960
rect 24268 13948 24274 14000
rect 24854 13988 24860 14000
rect 24320 13960 24860 13988
rect 24320 13929 24348 13960
rect 24854 13948 24860 13960
rect 24912 13948 24918 14000
rect 25682 13948 25688 14000
rect 25740 13988 25746 14000
rect 26988 13988 27016 14019
rect 25740 13960 27016 13988
rect 25740 13948 25746 13960
rect 23293 13923 23351 13929
rect 23293 13920 23305 13923
rect 23256 13892 23305 13920
rect 23256 13880 23262 13892
rect 23293 13889 23305 13892
rect 23339 13889 23351 13923
rect 23293 13883 23351 13889
rect 23753 13923 23811 13929
rect 23753 13889 23765 13923
rect 23799 13889 23811 13923
rect 23925 13895 23937 13929
rect 23971 13916 24072 13929
rect 24121 13923 24179 13929
rect 23971 13895 23983 13916
rect 23925 13889 23983 13895
rect 24121 13889 24133 13923
rect 24167 13889 24179 13923
rect 23753 13883 23811 13889
rect 24121 13883 24179 13889
rect 24305 13923 24363 13929
rect 24305 13889 24317 13923
rect 24351 13889 24363 13923
rect 24305 13883 24363 13889
rect 24670 13880 24676 13932
rect 24728 13920 24734 13932
rect 24949 13923 25007 13929
rect 24949 13920 24961 13923
rect 24728 13892 24961 13920
rect 24728 13880 24734 13892
rect 24949 13889 24961 13892
rect 24995 13889 25007 13923
rect 25130 13920 25136 13932
rect 25091 13892 25136 13920
rect 24949 13883 25007 13889
rect 25130 13880 25136 13892
rect 25188 13880 25194 13932
rect 25498 13920 25504 13932
rect 25459 13892 25504 13920
rect 25498 13880 25504 13892
rect 25556 13880 25562 13932
rect 26421 13923 26479 13929
rect 26421 13889 26433 13923
rect 26467 13920 26479 13923
rect 26510 13920 26516 13932
rect 26467 13892 26516 13920
rect 26467 13889 26479 13892
rect 26421 13883 26479 13889
rect 26510 13880 26516 13892
rect 26568 13880 26574 13932
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13889 27215 13923
rect 27157 13883 27215 13889
rect 21968 13824 22048 13852
rect 21968 13812 21974 13824
rect 22186 13812 22192 13864
rect 22244 13852 22250 13864
rect 22833 13855 22891 13861
rect 22833 13852 22845 13855
rect 22244 13824 22845 13852
rect 22244 13812 22250 13824
rect 22833 13821 22845 13824
rect 22879 13821 22891 13855
rect 22833 13815 22891 13821
rect 22925 13855 22983 13861
rect 22925 13821 22937 13855
rect 22971 13852 22983 13855
rect 23474 13852 23480 13864
rect 22971 13824 23480 13852
rect 22971 13821 22983 13824
rect 22925 13815 22983 13821
rect 23474 13812 23480 13824
rect 23532 13812 23538 13864
rect 24029 13855 24087 13861
rect 24029 13821 24041 13855
rect 24075 13821 24087 13855
rect 24029 13815 24087 13821
rect 20680 13756 20761 13784
rect 21269 13787 21327 13793
rect 20680 13744 20686 13756
rect 21269 13753 21281 13787
rect 21315 13784 21327 13787
rect 21542 13784 21548 13796
rect 21315 13756 21548 13784
rect 21315 13753 21327 13756
rect 21269 13747 21327 13753
rect 21542 13744 21548 13756
rect 21600 13744 21606 13796
rect 21726 13744 21732 13796
rect 21784 13744 21790 13796
rect 23106 13744 23112 13796
rect 23164 13784 23170 13796
rect 24044 13784 24072 13815
rect 24210 13812 24216 13864
rect 24268 13852 24274 13864
rect 24489 13855 24547 13861
rect 24489 13852 24501 13855
rect 24268 13824 24501 13852
rect 24268 13812 24274 13824
rect 24489 13821 24501 13824
rect 24535 13821 24547 13855
rect 24489 13815 24547 13821
rect 25225 13855 25283 13861
rect 25225 13821 25237 13855
rect 25271 13821 25283 13855
rect 25225 13815 25283 13821
rect 25317 13855 25375 13861
rect 25317 13821 25329 13855
rect 25363 13852 25375 13855
rect 25406 13852 25412 13864
rect 25363 13824 25412 13852
rect 25363 13821 25375 13824
rect 25317 13815 25375 13821
rect 23164 13756 24072 13784
rect 23164 13744 23170 13756
rect 25130 13744 25136 13796
rect 25188 13784 25194 13796
rect 25240 13784 25268 13815
rect 25406 13812 25412 13824
rect 25464 13852 25470 13864
rect 25866 13852 25872 13864
rect 25464 13824 25872 13852
rect 25464 13812 25470 13824
rect 25866 13812 25872 13824
rect 25924 13812 25930 13864
rect 26050 13812 26056 13864
rect 26108 13852 26114 13864
rect 27172 13852 27200 13883
rect 26108 13824 27200 13852
rect 26108 13812 26114 13824
rect 26878 13784 26884 13796
rect 25188 13756 25268 13784
rect 25608 13756 26884 13784
rect 25188 13744 25194 13756
rect 19518 13716 19524 13728
rect 18607 13688 19524 13716
rect 18049 13679 18107 13685
rect 19518 13676 19524 13688
rect 19576 13716 19582 13728
rect 20714 13716 20720 13728
rect 19576 13688 20720 13716
rect 19576 13676 19582 13688
rect 20714 13676 20720 13688
rect 20772 13676 20778 13728
rect 22094 13676 22100 13728
rect 22152 13716 22158 13728
rect 25608 13716 25636 13756
rect 26878 13744 26884 13756
rect 26936 13744 26942 13796
rect 22152 13688 25636 13716
rect 25685 13719 25743 13725
rect 22152 13676 22158 13688
rect 25685 13685 25697 13719
rect 25731 13716 25743 13719
rect 26142 13716 26148 13728
rect 25731 13688 26148 13716
rect 25731 13685 25743 13688
rect 25685 13679 25743 13685
rect 26142 13676 26148 13688
rect 26200 13676 26206 13728
rect 1104 13626 28060 13648
rect 1104 13574 5442 13626
rect 5494 13574 5506 13626
rect 5558 13574 5570 13626
rect 5622 13574 5634 13626
rect 5686 13574 5698 13626
rect 5750 13574 14428 13626
rect 14480 13574 14492 13626
rect 14544 13574 14556 13626
rect 14608 13574 14620 13626
rect 14672 13574 14684 13626
rect 14736 13574 23413 13626
rect 23465 13574 23477 13626
rect 23529 13574 23541 13626
rect 23593 13574 23605 13626
rect 23657 13574 23669 13626
rect 23721 13574 28060 13626
rect 1104 13552 28060 13574
rect 5261 13515 5319 13521
rect 5261 13481 5273 13515
rect 5307 13512 5319 13515
rect 5350 13512 5356 13524
rect 5307 13484 5356 13512
rect 5307 13481 5319 13484
rect 5261 13475 5319 13481
rect 5350 13472 5356 13484
rect 5408 13472 5414 13524
rect 7285 13515 7343 13521
rect 7285 13512 7297 13515
rect 6656 13484 7297 13512
rect 3878 13404 3884 13456
rect 3936 13444 3942 13456
rect 6656 13444 6684 13484
rect 7285 13481 7297 13484
rect 7331 13481 7343 13515
rect 7285 13475 7343 13481
rect 8297 13515 8355 13521
rect 8297 13481 8309 13515
rect 8343 13512 8355 13515
rect 8478 13512 8484 13524
rect 8343 13484 8484 13512
rect 8343 13481 8355 13484
rect 8297 13475 8355 13481
rect 8478 13472 8484 13484
rect 8536 13472 8542 13524
rect 10686 13512 10692 13524
rect 8864 13484 10692 13512
rect 3936 13416 6684 13444
rect 3936 13404 3942 13416
rect 4338 13336 4344 13388
rect 4396 13376 4402 13388
rect 4617 13379 4675 13385
rect 4617 13376 4629 13379
rect 4396 13348 4629 13376
rect 4396 13336 4402 13348
rect 4617 13345 4629 13348
rect 4663 13345 4675 13379
rect 4617 13339 4675 13345
rect 5166 13336 5172 13388
rect 5224 13376 5230 13388
rect 5353 13379 5411 13385
rect 5353 13376 5365 13379
rect 5224 13348 5365 13376
rect 5224 13336 5230 13348
rect 5353 13345 5365 13348
rect 5399 13345 5411 13379
rect 5353 13339 5411 13345
rect 1581 13311 1639 13317
rect 1581 13277 1593 13311
rect 1627 13308 1639 13311
rect 1670 13308 1676 13320
rect 1627 13280 1676 13308
rect 1627 13277 1639 13280
rect 1581 13271 1639 13277
rect 1670 13268 1676 13280
rect 1728 13268 1734 13320
rect 6656 13317 6684 13416
rect 6733 13447 6791 13453
rect 6733 13413 6745 13447
rect 6779 13444 6791 13447
rect 8662 13444 8668 13456
rect 6779 13416 8668 13444
rect 6779 13413 6791 13416
rect 6733 13407 6791 13413
rect 8662 13404 8668 13416
rect 8720 13404 8726 13456
rect 8864 13376 8892 13484
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 14090 13472 14096 13524
rect 14148 13512 14154 13524
rect 15010 13512 15016 13524
rect 14148 13484 15016 13512
rect 14148 13472 14154 13484
rect 15010 13472 15016 13484
rect 15068 13472 15074 13524
rect 16574 13472 16580 13524
rect 16632 13512 16638 13524
rect 17586 13512 17592 13524
rect 16632 13484 17592 13512
rect 16632 13472 16638 13484
rect 17586 13472 17592 13484
rect 17644 13472 17650 13524
rect 18782 13512 18788 13524
rect 18248 13484 18788 13512
rect 11054 13404 11060 13456
rect 11112 13444 11118 13456
rect 11514 13444 11520 13456
rect 11112 13416 11520 13444
rect 11112 13404 11118 13416
rect 11514 13404 11520 13416
rect 11572 13404 11578 13456
rect 18248 13444 18276 13484
rect 18782 13472 18788 13484
rect 18840 13512 18846 13524
rect 19058 13512 19064 13524
rect 18840 13484 19064 13512
rect 18840 13472 18846 13484
rect 19058 13472 19064 13484
rect 19116 13472 19122 13524
rect 19889 13515 19947 13521
rect 19889 13481 19901 13515
rect 19935 13512 19947 13515
rect 20346 13512 20352 13524
rect 19935 13484 20352 13512
rect 19935 13481 19947 13484
rect 19889 13475 19947 13481
rect 20346 13472 20352 13484
rect 20404 13472 20410 13524
rect 20898 13472 20904 13524
rect 20956 13512 20962 13524
rect 21726 13512 21732 13524
rect 20956 13484 21732 13512
rect 20956 13472 20962 13484
rect 21726 13472 21732 13484
rect 21784 13472 21790 13524
rect 22186 13472 22192 13524
rect 22244 13512 22250 13524
rect 23014 13512 23020 13524
rect 22244 13484 23020 13512
rect 22244 13472 22250 13484
rect 23014 13472 23020 13484
rect 23072 13472 23078 13524
rect 26234 13512 26240 13524
rect 23492 13484 26240 13512
rect 23492 13456 23520 13484
rect 26234 13472 26240 13484
rect 26292 13472 26298 13524
rect 26878 13472 26884 13524
rect 26936 13512 26942 13524
rect 27341 13515 27399 13521
rect 27341 13512 27353 13515
rect 26936 13484 27353 13512
rect 26936 13472 26942 13484
rect 27341 13481 27353 13484
rect 27387 13481 27399 13515
rect 27341 13475 27399 13481
rect 22094 13444 22100 13456
rect 17425 13416 18276 13444
rect 19306 13416 22100 13444
rect 10502 13376 10508 13388
rect 8404 13348 8892 13376
rect 8956 13348 10508 13376
rect 6641 13311 6699 13317
rect 6641 13277 6653 13311
rect 6687 13277 6699 13311
rect 6641 13271 6699 13277
rect 6733 13311 6791 13317
rect 6733 13277 6745 13311
rect 6779 13308 6791 13311
rect 7006 13308 7012 13320
rect 6779 13280 7012 13308
rect 6779 13277 6791 13280
rect 6733 13271 6791 13277
rect 7006 13268 7012 13280
rect 7064 13268 7070 13320
rect 8404 13317 8432 13348
rect 7193 13311 7251 13317
rect 7193 13277 7205 13311
rect 7239 13277 7251 13311
rect 7193 13271 7251 13277
rect 8205 13311 8263 13317
rect 8205 13277 8217 13311
rect 8251 13308 8263 13311
rect 8389 13311 8447 13317
rect 8251 13280 8340 13308
rect 8251 13277 8263 13280
rect 8205 13271 8263 13277
rect 1848 13243 1906 13249
rect 1848 13209 1860 13243
rect 1894 13240 1906 13243
rect 2498 13240 2504 13252
rect 1894 13212 2504 13240
rect 1894 13209 1906 13212
rect 1848 13203 1906 13209
rect 2498 13200 2504 13212
rect 2556 13200 2562 13252
rect 4433 13243 4491 13249
rect 4433 13209 4445 13243
rect 4479 13240 4491 13243
rect 4614 13240 4620 13252
rect 4479 13212 4620 13240
rect 4479 13209 4491 13212
rect 4433 13203 4491 13209
rect 4614 13200 4620 13212
rect 4672 13200 4678 13252
rect 5077 13243 5135 13249
rect 5077 13209 5089 13243
rect 5123 13209 5135 13243
rect 5442 13240 5448 13252
rect 5403 13212 5448 13240
rect 5077 13203 5135 13209
rect 2961 13175 3019 13181
rect 2961 13141 2973 13175
rect 3007 13172 3019 13175
rect 4062 13172 4068 13184
rect 3007 13144 4068 13172
rect 3007 13141 3019 13144
rect 2961 13135 3019 13141
rect 4062 13132 4068 13144
rect 4120 13172 4126 13184
rect 5092 13172 5120 13203
rect 5442 13200 5448 13212
rect 5500 13200 5506 13252
rect 6457 13243 6515 13249
rect 6457 13209 6469 13243
rect 6503 13240 6515 13243
rect 7208 13240 7236 13271
rect 6503 13212 7236 13240
rect 6503 13209 6515 13212
rect 6457 13203 6515 13209
rect 4120 13144 5120 13172
rect 5169 13175 5227 13181
rect 4120 13132 4126 13144
rect 5169 13141 5181 13175
rect 5215 13172 5227 13175
rect 6472 13172 6500 13203
rect 5215 13144 6500 13172
rect 7653 13175 7711 13181
rect 5215 13141 5227 13144
rect 5169 13135 5227 13141
rect 7653 13141 7665 13175
rect 7699 13172 7711 13175
rect 7926 13172 7932 13184
rect 7699 13144 7932 13172
rect 7699 13141 7711 13144
rect 7653 13135 7711 13141
rect 7926 13132 7932 13144
rect 7984 13132 7990 13184
rect 8312 13172 8340 13280
rect 8389 13277 8401 13311
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 8478 13268 8484 13320
rect 8536 13308 8542 13320
rect 8956 13317 8984 13348
rect 10502 13336 10508 13348
rect 10560 13336 10566 13388
rect 11330 13376 11336 13388
rect 11291 13348 11336 13376
rect 11330 13336 11336 13348
rect 11388 13376 11394 13388
rect 12161 13379 12219 13385
rect 12161 13376 12173 13379
rect 11388 13348 12173 13376
rect 11388 13336 11394 13348
rect 12161 13345 12173 13348
rect 12207 13345 12219 13379
rect 12161 13339 12219 13345
rect 14553 13379 14611 13385
rect 14553 13345 14565 13379
rect 14599 13376 14611 13379
rect 15930 13376 15936 13388
rect 14599 13348 15936 13376
rect 14599 13345 14611 13348
rect 14553 13339 14611 13345
rect 15930 13336 15936 13348
rect 15988 13376 15994 13388
rect 17425 13376 17453 13416
rect 19306 13376 19334 13416
rect 22094 13404 22100 13416
rect 22152 13404 22158 13456
rect 23474 13404 23480 13456
rect 23532 13404 23538 13456
rect 15988 13348 17453 13376
rect 15988 13336 15994 13348
rect 8941 13311 8999 13317
rect 8941 13308 8953 13311
rect 8536 13280 8953 13308
rect 8536 13268 8542 13280
rect 8941 13277 8953 13280
rect 8987 13277 8999 13311
rect 8941 13271 8999 13277
rect 9217 13311 9275 13317
rect 9217 13277 9229 13311
rect 9263 13308 9275 13311
rect 9674 13308 9680 13320
rect 9263 13280 9680 13308
rect 9263 13277 9275 13280
rect 9217 13271 9275 13277
rect 9674 13268 9680 13280
rect 9732 13308 9738 13320
rect 11517 13311 11575 13317
rect 11517 13308 11529 13311
rect 9732 13280 11529 13308
rect 9732 13268 9738 13280
rect 11517 13277 11529 13280
rect 11563 13277 11575 13311
rect 11517 13271 11575 13277
rect 12342 13268 12348 13320
rect 12400 13308 12406 13320
rect 12437 13311 12495 13317
rect 12437 13308 12449 13311
rect 12400 13280 12449 13308
rect 12400 13268 12406 13280
rect 12437 13277 12449 13280
rect 12483 13308 12495 13311
rect 13538 13308 13544 13320
rect 12483 13280 13544 13308
rect 12483 13277 12495 13280
rect 12437 13271 12495 13277
rect 13538 13268 13544 13280
rect 13596 13268 13602 13320
rect 14274 13308 14280 13320
rect 14235 13280 14280 13308
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 15378 13268 15384 13320
rect 15436 13308 15442 13320
rect 15565 13311 15623 13317
rect 15565 13308 15577 13311
rect 15436 13280 15577 13308
rect 15436 13268 15442 13280
rect 15565 13277 15577 13280
rect 15611 13277 15623 13311
rect 15565 13271 15623 13277
rect 15654 13268 15660 13320
rect 15712 13308 15718 13320
rect 16045 13317 16073 13348
rect 16030 13311 16088 13317
rect 15712 13280 15757 13308
rect 15712 13268 15718 13280
rect 16030 13277 16042 13311
rect 16076 13277 16088 13311
rect 16942 13308 16948 13320
rect 16903 13280 16948 13308
rect 16030 13271 16088 13277
rect 16942 13268 16948 13280
rect 17000 13268 17006 13320
rect 17126 13317 17132 13320
rect 17093 13311 17132 13317
rect 17093 13277 17105 13311
rect 17093 13271 17132 13277
rect 17126 13268 17132 13271
rect 17184 13268 17190 13320
rect 17425 13317 17453 13348
rect 18156 13348 19334 13376
rect 17410 13311 17468 13317
rect 17410 13277 17422 13311
rect 17456 13277 17468 13311
rect 17410 13271 17468 13277
rect 17770 13268 17776 13320
rect 17828 13308 17834 13320
rect 18156 13317 18184 13348
rect 19886 13336 19892 13388
rect 19944 13376 19950 13388
rect 19944 13348 20116 13376
rect 19944 13336 19950 13348
rect 20088 13320 20116 13348
rect 20714 13336 20720 13388
rect 20772 13376 20778 13388
rect 20901 13379 20959 13385
rect 20901 13376 20913 13379
rect 20772 13348 20913 13376
rect 20772 13336 20778 13348
rect 20901 13345 20913 13348
rect 20947 13345 20959 13379
rect 20901 13339 20959 13345
rect 23566 13336 23572 13388
rect 23624 13376 23630 13388
rect 25041 13379 25099 13385
rect 25041 13376 25053 13379
rect 23624 13348 25053 13376
rect 23624 13336 23630 13348
rect 25041 13345 25053 13348
rect 25087 13345 25099 13379
rect 25041 13339 25099 13345
rect 25133 13379 25191 13385
rect 25133 13345 25145 13379
rect 25179 13376 25191 13379
rect 25406 13376 25412 13388
rect 25179 13348 25412 13376
rect 25179 13345 25191 13348
rect 25133 13339 25191 13345
rect 25406 13336 25412 13348
rect 25464 13336 25470 13388
rect 18049 13311 18107 13317
rect 18049 13308 18061 13311
rect 17828 13280 18061 13308
rect 17828 13268 17834 13280
rect 18049 13277 18061 13280
rect 18095 13277 18107 13311
rect 18049 13271 18107 13277
rect 18142 13311 18200 13317
rect 18142 13277 18154 13311
rect 18188 13277 18200 13311
rect 18417 13311 18475 13317
rect 18417 13310 18429 13311
rect 18340 13308 18429 13310
rect 18142 13271 18200 13277
rect 18248 13282 18429 13308
rect 18248 13280 18368 13282
rect 9030 13200 9036 13252
rect 9088 13240 9094 13252
rect 10597 13243 10655 13249
rect 10597 13240 10609 13243
rect 9088 13212 10609 13240
rect 9088 13200 9094 13212
rect 10597 13209 10609 13212
rect 10643 13209 10655 13243
rect 10597 13203 10655 13209
rect 11701 13243 11759 13249
rect 11701 13209 11713 13243
rect 11747 13240 11759 13243
rect 15838 13240 15844 13252
rect 11747 13212 15844 13240
rect 11747 13209 11759 13212
rect 11701 13203 11759 13209
rect 15838 13200 15844 13212
rect 15896 13200 15902 13252
rect 15930 13200 15936 13252
rect 15988 13240 15994 13252
rect 17221 13243 17279 13249
rect 15988 13212 16033 13240
rect 15988 13200 15994 13212
rect 17221 13209 17233 13243
rect 17267 13209 17279 13243
rect 17221 13203 17279 13209
rect 17313 13243 17371 13249
rect 17313 13209 17325 13243
rect 17359 13240 17371 13243
rect 17954 13240 17960 13252
rect 17359 13212 17960 13240
rect 17359 13209 17371 13212
rect 17313 13203 17371 13209
rect 9766 13172 9772 13184
rect 8312 13144 9772 13172
rect 9766 13132 9772 13144
rect 9824 13172 9830 13184
rect 10778 13172 10784 13184
rect 9824 13144 10784 13172
rect 9824 13132 9830 13144
rect 10778 13132 10784 13144
rect 10836 13132 10842 13184
rect 14090 13132 14096 13184
rect 14148 13172 14154 13184
rect 16209 13175 16267 13181
rect 16209 13172 16221 13175
rect 14148 13144 16221 13172
rect 14148 13132 14154 13144
rect 16209 13141 16221 13144
rect 16255 13141 16267 13175
rect 17236 13172 17264 13203
rect 17954 13200 17960 13212
rect 18012 13200 18018 13252
rect 17862 13172 17868 13184
rect 17236 13144 17868 13172
rect 16209 13135 16267 13141
rect 17862 13132 17868 13144
rect 17920 13132 17926 13184
rect 18046 13132 18052 13184
rect 18104 13172 18110 13184
rect 18248 13172 18276 13280
rect 18417 13277 18429 13282
rect 18463 13277 18475 13311
rect 18417 13271 18475 13277
rect 18555 13311 18613 13317
rect 18555 13277 18567 13311
rect 18601 13308 18613 13311
rect 18782 13308 18788 13320
rect 18601 13280 18788 13308
rect 18601 13277 18613 13280
rect 18555 13271 18613 13277
rect 18782 13268 18788 13280
rect 18840 13268 18846 13320
rect 19245 13311 19303 13317
rect 19245 13277 19257 13311
rect 19291 13277 19303 13311
rect 19245 13271 19303 13277
rect 19393 13311 19451 13317
rect 19393 13277 19405 13311
rect 19439 13277 19451 13311
rect 19621 13311 19679 13317
rect 19621 13298 19633 13311
rect 19667 13298 19679 13311
rect 19393 13271 19451 13277
rect 18325 13243 18383 13249
rect 18325 13209 18337 13243
rect 18371 13240 18383 13243
rect 18371 13212 18460 13240
rect 18371 13209 18383 13212
rect 18325 13203 18383 13209
rect 18432 13184 18460 13212
rect 19150 13200 19156 13252
rect 19208 13240 19214 13252
rect 19260 13240 19288 13271
rect 19208 13212 19288 13240
rect 19208 13200 19214 13212
rect 18104 13144 18276 13172
rect 18104 13132 18110 13144
rect 18414 13132 18420 13184
rect 18472 13132 18478 13184
rect 18506 13132 18512 13184
rect 18564 13172 18570 13184
rect 18693 13175 18751 13181
rect 18693 13172 18705 13175
rect 18564 13144 18705 13172
rect 18564 13132 18570 13144
rect 18693 13141 18705 13144
rect 18739 13141 18751 13175
rect 19408 13172 19436 13271
rect 19518 13240 19524 13252
rect 19479 13212 19524 13240
rect 19518 13200 19524 13212
rect 19576 13200 19582 13252
rect 19610 13246 19616 13298
rect 19668 13271 19679 13298
rect 19710 13311 19768 13317
rect 19710 13277 19722 13311
rect 19756 13298 19768 13311
rect 19756 13277 20015 13298
rect 19710 13271 20015 13277
rect 19668 13246 19674 13271
rect 19720 13270 20015 13271
rect 19987 13240 20015 13270
rect 20070 13268 20076 13320
rect 20128 13268 20134 13320
rect 20622 13308 20628 13320
rect 20583 13280 20628 13308
rect 20622 13268 20628 13280
rect 20680 13308 20686 13320
rect 21818 13308 21824 13320
rect 20680 13280 21824 13308
rect 20680 13268 20686 13280
rect 21818 13268 21824 13280
rect 21876 13268 21882 13320
rect 21910 13268 21916 13320
rect 21968 13308 21974 13320
rect 22373 13311 22431 13317
rect 22373 13308 22385 13311
rect 21968 13280 22385 13308
rect 21968 13268 21974 13280
rect 22373 13277 22385 13280
rect 22419 13308 22431 13311
rect 23750 13308 23756 13320
rect 22419 13280 23756 13308
rect 22419 13277 22431 13280
rect 22373 13271 22431 13277
rect 23750 13268 23756 13280
rect 23808 13268 23814 13320
rect 24670 13268 24676 13320
rect 24728 13308 24734 13320
rect 24765 13311 24823 13317
rect 24765 13308 24777 13311
rect 24728 13280 24777 13308
rect 24728 13268 24734 13280
rect 24765 13277 24777 13280
rect 24811 13277 24823 13311
rect 24946 13308 24952 13320
rect 24907 13280 24952 13308
rect 24765 13271 24823 13277
rect 24946 13268 24952 13280
rect 25004 13268 25010 13320
rect 25317 13311 25375 13317
rect 25317 13277 25329 13311
rect 25363 13308 25375 13311
rect 25590 13308 25596 13320
rect 25363 13280 25596 13308
rect 25363 13277 25375 13280
rect 25317 13271 25375 13277
rect 25590 13268 25596 13280
rect 25648 13268 25654 13320
rect 25958 13308 25964 13320
rect 25919 13280 25964 13308
rect 25958 13268 25964 13280
rect 26016 13268 26022 13320
rect 21174 13240 21180 13252
rect 19987 13212 21180 13240
rect 21174 13200 21180 13212
rect 21232 13200 21238 13252
rect 22640 13243 22698 13249
rect 22640 13209 22652 13243
rect 22686 13240 22698 13243
rect 23290 13240 23296 13252
rect 22686 13212 23296 13240
rect 22686 13209 22698 13212
rect 22640 13203 22698 13209
rect 23290 13200 23296 13212
rect 23348 13200 23354 13252
rect 26228 13243 26286 13249
rect 26228 13209 26240 13243
rect 26274 13240 26286 13243
rect 26418 13240 26424 13252
rect 26274 13212 26424 13240
rect 26274 13209 26286 13212
rect 26228 13203 26286 13209
rect 26418 13200 26424 13212
rect 26476 13200 26482 13252
rect 20070 13172 20076 13184
rect 19408 13144 20076 13172
rect 18693 13135 18751 13141
rect 20070 13132 20076 13144
rect 20128 13132 20134 13184
rect 20714 13132 20720 13184
rect 20772 13172 20778 13184
rect 22094 13172 22100 13184
rect 20772 13144 22100 13172
rect 20772 13132 20778 13144
rect 22094 13132 22100 13144
rect 22152 13132 22158 13184
rect 22278 13132 22284 13184
rect 22336 13172 22342 13184
rect 23753 13175 23811 13181
rect 23753 13172 23765 13175
rect 22336 13144 23765 13172
rect 22336 13132 22342 13144
rect 23753 13141 23765 13144
rect 23799 13172 23811 13175
rect 24026 13172 24032 13184
rect 23799 13144 24032 13172
rect 23799 13141 23811 13144
rect 23753 13135 23811 13141
rect 24026 13132 24032 13144
rect 24084 13132 24090 13184
rect 25406 13132 25412 13184
rect 25464 13172 25470 13184
rect 25501 13175 25559 13181
rect 25501 13172 25513 13175
rect 25464 13144 25513 13172
rect 25464 13132 25470 13144
rect 25501 13141 25513 13144
rect 25547 13141 25559 13175
rect 25501 13135 25559 13141
rect 1104 13082 28060 13104
rect 1104 13030 9935 13082
rect 9987 13030 9999 13082
rect 10051 13030 10063 13082
rect 10115 13030 10127 13082
rect 10179 13030 10191 13082
rect 10243 13030 18920 13082
rect 18972 13030 18984 13082
rect 19036 13030 19048 13082
rect 19100 13030 19112 13082
rect 19164 13030 19176 13082
rect 19228 13030 28060 13082
rect 1104 13008 28060 13030
rect 3053 12971 3111 12977
rect 3053 12937 3065 12971
rect 3099 12968 3111 12971
rect 4246 12968 4252 12980
rect 3099 12940 4252 12968
rect 3099 12937 3111 12940
rect 3053 12931 3111 12937
rect 4246 12928 4252 12940
rect 4304 12928 4310 12980
rect 4614 12928 4620 12980
rect 4672 12968 4678 12980
rect 6733 12971 6791 12977
rect 6733 12968 6745 12971
rect 4672 12940 6745 12968
rect 4672 12928 4678 12940
rect 6733 12937 6745 12940
rect 6779 12937 6791 12971
rect 7466 12968 7472 12980
rect 6733 12931 6791 12937
rect 7392 12940 7472 12968
rect 2685 12903 2743 12909
rect 2685 12869 2697 12903
rect 2731 12900 2743 12903
rect 3602 12900 3608 12912
rect 2731 12872 3608 12900
rect 2731 12869 2743 12872
rect 2685 12863 2743 12869
rect 3602 12860 3608 12872
rect 3660 12860 3666 12912
rect 4338 12900 4344 12912
rect 3988 12872 4344 12900
rect 1765 12835 1823 12841
rect 1765 12801 1777 12835
rect 1811 12801 1823 12835
rect 1765 12795 1823 12801
rect 1949 12835 2007 12841
rect 1949 12801 1961 12835
rect 1995 12832 2007 12835
rect 2038 12832 2044 12844
rect 1995 12804 2044 12832
rect 1995 12801 2007 12804
rect 1949 12795 2007 12801
rect 1780 12764 1808 12795
rect 2038 12792 2044 12804
rect 2096 12832 2102 12844
rect 3988 12841 4016 12872
rect 4338 12860 4344 12872
rect 4396 12860 4402 12912
rect 4706 12860 4712 12912
rect 4764 12900 4770 12912
rect 4890 12900 4896 12912
rect 4764 12872 4896 12900
rect 4764 12860 4770 12872
rect 4890 12860 4896 12872
rect 4948 12860 4954 12912
rect 5534 12860 5540 12912
rect 5592 12900 5598 12912
rect 6362 12900 6368 12912
rect 5592 12872 6368 12900
rect 5592 12860 5598 12872
rect 6362 12860 6368 12872
rect 6420 12860 6426 12912
rect 6641 12903 6699 12909
rect 6641 12869 6653 12903
rect 6687 12900 6699 12903
rect 6914 12900 6920 12912
rect 6687 12872 6920 12900
rect 6687 12869 6699 12872
rect 6641 12863 6699 12869
rect 6914 12860 6920 12872
rect 6972 12860 6978 12912
rect 2869 12835 2927 12841
rect 2869 12832 2881 12835
rect 2096 12804 2881 12832
rect 2096 12792 2102 12804
rect 2869 12801 2881 12804
rect 2915 12801 2927 12835
rect 2869 12795 2927 12801
rect 3973 12835 4031 12841
rect 3973 12801 3985 12835
rect 4019 12801 4031 12835
rect 3973 12795 4031 12801
rect 4240 12835 4298 12841
rect 4240 12801 4252 12835
rect 4286 12832 4298 12835
rect 5074 12832 5080 12844
rect 4286 12804 5080 12832
rect 4286 12801 4298 12804
rect 4240 12795 4298 12801
rect 5074 12792 5080 12804
rect 5132 12792 5138 12844
rect 7006 12792 7012 12844
rect 7064 12792 7070 12844
rect 3418 12764 3424 12776
rect 1780 12736 3424 12764
rect 3418 12724 3424 12736
rect 3476 12724 3482 12776
rect 6362 12724 6368 12776
rect 6420 12764 6426 12776
rect 7024 12764 7052 12792
rect 6420 12736 7052 12764
rect 6420 12724 6426 12736
rect 5074 12656 5080 12708
rect 5132 12696 5138 12708
rect 5353 12699 5411 12705
rect 5353 12696 5365 12699
rect 5132 12668 5365 12696
rect 5132 12656 5138 12668
rect 5353 12665 5365 12668
rect 5399 12696 5411 12699
rect 5442 12696 5448 12708
rect 5399 12668 5448 12696
rect 5399 12665 5411 12668
rect 5353 12659 5411 12665
rect 5442 12656 5448 12668
rect 5500 12656 5506 12708
rect 7392 12696 7420 12940
rect 7466 12928 7472 12940
rect 7524 12928 7530 12980
rect 8297 12971 8355 12977
rect 8297 12937 8309 12971
rect 8343 12968 8355 12971
rect 8478 12968 8484 12980
rect 8343 12940 8484 12968
rect 8343 12937 8355 12940
rect 8297 12931 8355 12937
rect 8478 12928 8484 12940
rect 8536 12928 8542 12980
rect 9217 12971 9275 12977
rect 9217 12937 9229 12971
rect 9263 12968 9275 12971
rect 10318 12968 10324 12980
rect 9263 12940 10324 12968
rect 9263 12937 9275 12940
rect 9217 12931 9275 12937
rect 9306 12900 9312 12912
rect 7484 12872 9312 12900
rect 7484 12841 7512 12872
rect 9306 12860 9312 12872
rect 9364 12860 9370 12912
rect 10152 12909 10180 12940
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 11146 12928 11152 12980
rect 11204 12968 11210 12980
rect 11701 12971 11759 12977
rect 11701 12968 11713 12971
rect 11204 12940 11713 12968
rect 11204 12928 11210 12940
rect 11701 12937 11713 12940
rect 11747 12937 11759 12971
rect 11701 12931 11759 12937
rect 13357 12971 13415 12977
rect 13357 12937 13369 12971
rect 13403 12968 13415 12971
rect 13998 12968 14004 12980
rect 13403 12940 14004 12968
rect 13403 12937 13415 12940
rect 13357 12931 13415 12937
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 16666 12928 16672 12980
rect 16724 12968 16730 12980
rect 17773 12971 17831 12977
rect 17773 12968 17785 12971
rect 16724 12940 17785 12968
rect 16724 12928 16730 12940
rect 10137 12903 10195 12909
rect 10137 12869 10149 12903
rect 10183 12869 10195 12903
rect 10137 12863 10195 12869
rect 10229 12903 10287 12909
rect 10229 12869 10241 12903
rect 10275 12900 10287 12903
rect 10778 12900 10784 12912
rect 10275 12872 10784 12900
rect 10275 12869 10287 12872
rect 10229 12863 10287 12869
rect 10778 12860 10784 12872
rect 10836 12900 10842 12912
rect 10962 12900 10968 12912
rect 10836 12872 10968 12900
rect 10836 12860 10842 12872
rect 10962 12860 10968 12872
rect 11020 12860 11026 12912
rect 14185 12903 14243 12909
rect 14185 12900 14197 12903
rect 11348 12872 14197 12900
rect 7469 12835 7527 12841
rect 7469 12801 7481 12835
rect 7515 12801 7527 12835
rect 7926 12832 7932 12844
rect 7887 12804 7932 12832
rect 7469 12795 7527 12801
rect 7926 12792 7932 12804
rect 7984 12792 7990 12844
rect 8386 12792 8392 12844
rect 8444 12832 8450 12844
rect 9122 12841 9128 12844
rect 8757 12835 8815 12841
rect 8757 12832 8769 12835
rect 8444 12804 8769 12832
rect 8444 12792 8450 12804
rect 8757 12801 8769 12804
rect 8803 12801 8815 12835
rect 8757 12795 8815 12801
rect 9073 12835 9128 12841
rect 9073 12801 9085 12835
rect 9119 12801 9128 12835
rect 9073 12795 9128 12801
rect 9122 12792 9128 12795
rect 9180 12792 9186 12844
rect 9214 12792 9220 12844
rect 9272 12832 9278 12844
rect 9766 12832 9772 12844
rect 9272 12804 9772 12832
rect 9272 12792 9278 12804
rect 8021 12767 8079 12773
rect 8021 12733 8033 12767
rect 8067 12764 8079 12767
rect 8846 12764 8852 12776
rect 8067 12736 8852 12764
rect 8067 12733 8079 12736
rect 8021 12727 8079 12733
rect 7392 12668 7880 12696
rect 7852 12640 7880 12668
rect 8036 12640 8064 12727
rect 8846 12724 8852 12736
rect 8904 12724 8910 12776
rect 2133 12631 2191 12637
rect 2133 12597 2145 12631
rect 2179 12628 2191 12631
rect 2682 12628 2688 12640
rect 2179 12600 2688 12628
rect 2179 12597 2191 12600
rect 2133 12591 2191 12597
rect 2682 12588 2688 12600
rect 2740 12588 2746 12640
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 4338 12628 4344 12640
rect 4212 12600 4344 12628
rect 4212 12588 4218 12600
rect 4338 12588 4344 12600
rect 4396 12588 4402 12640
rect 6638 12588 6644 12640
rect 6696 12628 6702 12640
rect 6822 12628 6828 12640
rect 6696 12600 6828 12628
rect 6696 12588 6702 12600
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 7285 12631 7343 12637
rect 7285 12597 7297 12631
rect 7331 12628 7343 12631
rect 7374 12628 7380 12640
rect 7331 12600 7380 12628
rect 7331 12597 7343 12600
rect 7285 12591 7343 12597
rect 7374 12588 7380 12600
rect 7432 12588 7438 12640
rect 7834 12588 7840 12640
rect 7892 12588 7898 12640
rect 8018 12588 8024 12640
rect 8076 12588 8082 12640
rect 8113 12631 8171 12637
rect 8113 12597 8125 12631
rect 8159 12628 8171 12631
rect 8386 12628 8392 12640
rect 8159 12600 8392 12628
rect 8159 12597 8171 12600
rect 8113 12591 8171 12597
rect 8386 12588 8392 12600
rect 8444 12588 8450 12640
rect 8662 12588 8668 12640
rect 8720 12628 8726 12640
rect 8757 12631 8815 12637
rect 8757 12628 8769 12631
rect 8720 12600 8769 12628
rect 8720 12588 8726 12600
rect 8757 12597 8769 12600
rect 8803 12597 8815 12631
rect 9416 12628 9444 12804
rect 9766 12792 9772 12804
rect 9824 12792 9830 12844
rect 10042 12792 10048 12844
rect 10100 12832 10106 12844
rect 10367 12835 10425 12841
rect 10100 12804 10145 12832
rect 10100 12792 10106 12804
rect 10367 12801 10379 12835
rect 10413 12832 10425 12835
rect 11348 12832 11376 12872
rect 14185 12869 14197 12872
rect 14231 12900 14243 12903
rect 14274 12900 14280 12912
rect 14231 12872 14280 12900
rect 14231 12869 14243 12872
rect 14185 12863 14243 12869
rect 14274 12860 14280 12872
rect 14332 12860 14338 12912
rect 15105 12903 15163 12909
rect 15105 12869 15117 12903
rect 15151 12900 15163 12903
rect 16022 12900 16028 12912
rect 15151 12872 16028 12900
rect 15151 12869 15163 12872
rect 15105 12863 15163 12869
rect 16022 12860 16028 12872
rect 16080 12900 16086 12912
rect 16390 12900 16396 12912
rect 16080 12872 16396 12900
rect 16080 12860 16086 12872
rect 16390 12860 16396 12872
rect 16448 12860 16454 12912
rect 17512 12856 17540 12940
rect 17773 12937 17785 12940
rect 17819 12937 17831 12971
rect 17773 12931 17831 12937
rect 17862 12928 17868 12980
rect 17920 12968 17926 12980
rect 18414 12968 18420 12980
rect 17920 12940 18420 12968
rect 17920 12928 17926 12940
rect 18414 12928 18420 12940
rect 18472 12968 18478 12980
rect 19518 12968 19524 12980
rect 18472 12940 19524 12968
rect 18472 12928 18478 12940
rect 19518 12928 19524 12940
rect 19576 12928 19582 12980
rect 19610 12928 19616 12980
rect 19668 12968 19674 12980
rect 19705 12971 19763 12977
rect 19705 12968 19717 12971
rect 19668 12940 19717 12968
rect 19668 12928 19674 12940
rect 19705 12937 19717 12940
rect 19751 12937 19763 12971
rect 19705 12931 19763 12937
rect 20070 12928 20076 12980
rect 20128 12968 20134 12980
rect 21358 12968 21364 12980
rect 20128 12940 21364 12968
rect 20128 12928 20134 12940
rect 21358 12928 21364 12940
rect 21416 12928 21422 12980
rect 21818 12928 21824 12980
rect 21876 12968 21882 12980
rect 22002 12968 22008 12980
rect 21876 12940 22008 12968
rect 21876 12928 21882 12940
rect 22002 12928 22008 12940
rect 22060 12928 22066 12980
rect 22370 12928 22376 12980
rect 22428 12968 22434 12980
rect 22465 12971 22523 12977
rect 22465 12968 22477 12971
rect 22428 12940 22477 12968
rect 22428 12928 22434 12940
rect 22465 12937 22477 12940
rect 22511 12937 22523 12971
rect 22465 12931 22523 12937
rect 22833 12971 22891 12977
rect 22833 12937 22845 12971
rect 22879 12968 22891 12971
rect 24670 12968 24676 12980
rect 22879 12940 24676 12968
rect 22879 12937 22891 12940
rect 22833 12931 22891 12937
rect 24670 12928 24676 12940
rect 24728 12968 24734 12980
rect 25041 12971 25099 12977
rect 25041 12968 25053 12971
rect 24728 12940 25053 12968
rect 24728 12928 24734 12940
rect 25041 12937 25053 12940
rect 25087 12937 25099 12971
rect 25041 12931 25099 12937
rect 18138 12860 18144 12912
rect 18196 12900 18202 12912
rect 18322 12900 18328 12912
rect 18196 12872 18328 12900
rect 18196 12860 18202 12872
rect 18322 12860 18328 12872
rect 18380 12860 18386 12912
rect 18592 12903 18650 12909
rect 18592 12869 18604 12903
rect 18638 12900 18650 12903
rect 23474 12900 23480 12912
rect 18638 12872 23480 12900
rect 18638 12869 18650 12872
rect 18592 12863 18650 12869
rect 23474 12860 23480 12872
rect 23532 12860 23538 12912
rect 23750 12900 23756 12912
rect 23676 12872 23756 12900
rect 11514 12832 11520 12844
rect 10413 12804 11376 12832
rect 11475 12804 11520 12832
rect 10413 12802 10468 12804
rect 10413 12801 10425 12802
rect 10367 12795 10425 12801
rect 10382 12764 10410 12795
rect 11514 12792 11520 12804
rect 11572 12792 11578 12844
rect 12250 12832 12256 12844
rect 12211 12804 12256 12832
rect 12250 12792 12256 12804
rect 12308 12792 12314 12844
rect 12437 12835 12495 12841
rect 12437 12801 12449 12835
rect 12483 12801 12495 12835
rect 13262 12832 13268 12844
rect 13223 12804 13268 12832
rect 12437 12795 12495 12801
rect 9646 12736 10410 12764
rect 10505 12767 10563 12773
rect 9490 12656 9496 12708
rect 9548 12696 9554 12708
rect 9646 12696 9674 12736
rect 10505 12733 10517 12767
rect 10551 12764 10563 12767
rect 10594 12764 10600 12776
rect 10551 12736 10600 12764
rect 10551 12733 10563 12736
rect 10505 12727 10563 12733
rect 10594 12724 10600 12736
rect 10652 12724 10658 12776
rect 12158 12724 12164 12776
rect 12216 12764 12222 12776
rect 12452 12764 12480 12795
rect 13262 12792 13268 12804
rect 13320 12792 13326 12844
rect 14826 12792 14832 12844
rect 14884 12832 14890 12844
rect 14921 12835 14979 12841
rect 14921 12832 14933 12835
rect 14884 12804 14933 12832
rect 14884 12792 14890 12804
rect 14921 12801 14933 12804
rect 14967 12801 14979 12835
rect 14921 12795 14979 12801
rect 16117 12835 16175 12841
rect 16117 12801 16129 12835
rect 16163 12832 16175 12835
rect 16574 12832 16580 12844
rect 16163 12804 16580 12832
rect 16163 12801 16175 12804
rect 16117 12795 16175 12801
rect 13538 12764 13544 12776
rect 12216 12736 12480 12764
rect 13451 12736 13544 12764
rect 12216 12724 12222 12736
rect 13538 12724 13544 12736
rect 13596 12764 13602 12776
rect 14936 12764 14964 12795
rect 16574 12792 16580 12804
rect 16632 12792 16638 12844
rect 17126 12832 17132 12844
rect 17087 12804 17132 12832
rect 17126 12792 17132 12804
rect 17184 12792 17190 12844
rect 17512 12828 17623 12856
rect 13596 12736 14964 12764
rect 13596 12724 13602 12736
rect 15654 12724 15660 12776
rect 15712 12764 15718 12776
rect 17595 12764 17623 12828
rect 17681 12835 17739 12841
rect 17681 12801 17693 12835
rect 17727 12830 17739 12835
rect 18414 12832 18420 12844
rect 17788 12830 18420 12832
rect 17727 12804 18420 12830
rect 17727 12802 17816 12804
rect 17727 12801 17739 12802
rect 17681 12795 17739 12801
rect 18414 12792 18420 12804
rect 18472 12792 18478 12844
rect 19058 12792 19064 12844
rect 19116 12832 19122 12844
rect 20346 12832 20352 12844
rect 19116 12804 20352 12832
rect 19116 12792 19122 12804
rect 20346 12792 20352 12804
rect 20404 12792 20410 12844
rect 20714 12832 20720 12844
rect 20675 12804 20720 12832
rect 20714 12792 20720 12804
rect 20772 12792 20778 12844
rect 20898 12832 20904 12844
rect 20859 12804 20904 12832
rect 20898 12792 20904 12804
rect 20956 12792 20962 12844
rect 20993 12835 21051 12841
rect 20993 12801 21005 12835
rect 21039 12801 21051 12835
rect 20993 12795 21051 12801
rect 21085 12835 21143 12841
rect 21085 12801 21097 12835
rect 21131 12832 21143 12835
rect 21174 12832 21180 12844
rect 21131 12804 21180 12832
rect 21131 12801 21143 12804
rect 21085 12795 21143 12801
rect 18325 12767 18383 12773
rect 18325 12764 18337 12767
rect 15712 12736 17448 12764
rect 17595 12736 18337 12764
rect 15712 12724 15718 12736
rect 14366 12696 14372 12708
rect 9548 12668 9674 12696
rect 14279 12668 14372 12696
rect 9548 12656 9554 12668
rect 14366 12656 14372 12668
rect 14424 12696 14430 12708
rect 15194 12696 15200 12708
rect 14424 12668 15200 12696
rect 14424 12656 14430 12668
rect 15194 12656 15200 12668
rect 15252 12656 15258 12708
rect 15933 12699 15991 12705
rect 15933 12665 15945 12699
rect 15979 12696 15991 12699
rect 17310 12696 17316 12708
rect 15979 12668 17316 12696
rect 15979 12665 15991 12668
rect 15933 12659 15991 12665
rect 17310 12656 17316 12668
rect 17368 12656 17374 12708
rect 9861 12631 9919 12637
rect 9861 12628 9873 12631
rect 9416 12600 9873 12628
rect 8757 12591 8815 12597
rect 9861 12597 9873 12600
rect 9907 12597 9919 12631
rect 12342 12628 12348 12640
rect 12303 12600 12348 12628
rect 9861 12591 9919 12597
rect 12342 12588 12348 12600
rect 12400 12588 12406 12640
rect 12802 12588 12808 12640
rect 12860 12628 12866 12640
rect 12897 12631 12955 12637
rect 12897 12628 12909 12631
rect 12860 12600 12909 12628
rect 12860 12588 12866 12600
rect 12897 12597 12909 12600
rect 12943 12597 12955 12631
rect 12897 12591 12955 12597
rect 16022 12588 16028 12640
rect 16080 12628 16086 12640
rect 16206 12628 16212 12640
rect 16080 12600 16212 12628
rect 16080 12588 16086 12600
rect 16206 12588 16212 12600
rect 16264 12588 16270 12640
rect 16850 12588 16856 12640
rect 16908 12628 16914 12640
rect 16945 12631 17003 12637
rect 16945 12628 16957 12631
rect 16908 12600 16957 12628
rect 16908 12588 16914 12600
rect 16945 12597 16957 12600
rect 16991 12597 17003 12631
rect 17420 12628 17448 12736
rect 18325 12733 18337 12736
rect 18371 12733 18383 12767
rect 21008 12764 21036 12795
rect 21174 12792 21180 12804
rect 21232 12792 21238 12844
rect 22005 12835 22063 12841
rect 22005 12832 22017 12835
rect 21652 12804 22017 12832
rect 21542 12764 21548 12776
rect 21008 12736 21548 12764
rect 18325 12727 18383 12733
rect 21542 12724 21548 12736
rect 21600 12724 21606 12776
rect 21652 12696 21680 12804
rect 22005 12801 22017 12804
rect 22051 12801 22063 12835
rect 22005 12795 22063 12801
rect 22278 12792 22284 12844
rect 22336 12832 22342 12844
rect 22646 12832 22652 12844
rect 22336 12804 22652 12832
rect 22336 12792 22342 12804
rect 22646 12792 22652 12804
rect 22704 12792 22710 12844
rect 23676 12841 23704 12872
rect 23750 12860 23756 12872
rect 23808 12900 23814 12912
rect 25958 12900 25964 12912
rect 23808 12872 25964 12900
rect 23808 12860 23814 12872
rect 25958 12860 25964 12872
rect 26016 12860 26022 12912
rect 23934 12841 23940 12844
rect 23661 12835 23719 12841
rect 23661 12801 23673 12835
rect 23707 12801 23719 12835
rect 23661 12795 23719 12801
rect 23928 12795 23940 12841
rect 23992 12832 23998 12844
rect 23992 12804 24028 12832
rect 23934 12792 23940 12795
rect 23992 12792 23998 12804
rect 24854 12792 24860 12844
rect 24912 12832 24918 12844
rect 25774 12832 25780 12844
rect 24912 12804 25780 12832
rect 24912 12792 24918 12804
rect 25774 12792 25780 12804
rect 25832 12792 25838 12844
rect 26142 12832 26148 12844
rect 26103 12804 26148 12832
rect 26142 12792 26148 12804
rect 26200 12792 26206 12844
rect 27341 12835 27399 12841
rect 27341 12832 27353 12835
rect 26243 12804 27353 12832
rect 22922 12764 22928 12776
rect 22883 12736 22928 12764
rect 22922 12724 22928 12736
rect 22980 12724 22986 12776
rect 23109 12767 23167 12773
rect 23109 12733 23121 12767
rect 23155 12764 23167 12767
rect 23382 12764 23388 12776
rect 23155 12736 23388 12764
rect 23155 12733 23167 12736
rect 23109 12727 23167 12733
rect 23382 12724 23388 12736
rect 23440 12724 23446 12776
rect 24762 12724 24768 12776
rect 24820 12764 24826 12776
rect 26243 12764 26271 12804
rect 27341 12801 27353 12804
rect 27387 12801 27399 12835
rect 27341 12795 27399 12801
rect 24820 12736 26271 12764
rect 26421 12767 26479 12773
rect 24820 12724 24826 12736
rect 26421 12733 26433 12767
rect 26467 12764 26479 12767
rect 26602 12764 26608 12776
rect 26467 12736 26608 12764
rect 26467 12733 26479 12736
rect 26421 12727 26479 12733
rect 26602 12724 26608 12736
rect 26660 12724 26666 12776
rect 19996 12668 21680 12696
rect 19996 12640 20024 12668
rect 21726 12656 21732 12708
rect 21784 12696 21790 12708
rect 23566 12696 23572 12708
rect 21784 12668 23572 12696
rect 21784 12656 21790 12668
rect 23566 12656 23572 12668
rect 23624 12656 23630 12708
rect 25961 12699 26019 12705
rect 25961 12665 25973 12699
rect 26007 12696 26019 12699
rect 26234 12696 26240 12708
rect 26007 12668 26240 12696
rect 26007 12665 26019 12668
rect 25961 12659 26019 12665
rect 26234 12656 26240 12668
rect 26292 12656 26298 12708
rect 19886 12628 19892 12640
rect 17420 12600 19892 12628
rect 16945 12591 17003 12597
rect 19886 12588 19892 12600
rect 19944 12588 19950 12640
rect 19978 12588 19984 12640
rect 20036 12588 20042 12640
rect 20346 12588 20352 12640
rect 20404 12628 20410 12640
rect 21269 12631 21327 12637
rect 21269 12628 21281 12631
rect 20404 12600 21281 12628
rect 20404 12588 20410 12600
rect 21269 12597 21281 12600
rect 21315 12597 21327 12631
rect 21269 12591 21327 12597
rect 21358 12588 21364 12640
rect 21416 12628 21422 12640
rect 21634 12628 21640 12640
rect 21416 12600 21640 12628
rect 21416 12588 21422 12600
rect 21634 12588 21640 12600
rect 21692 12588 21698 12640
rect 21821 12631 21879 12637
rect 21821 12597 21833 12631
rect 21867 12628 21879 12631
rect 22094 12628 22100 12640
rect 21867 12600 22100 12628
rect 21867 12597 21879 12600
rect 21821 12591 21879 12597
rect 22094 12588 22100 12600
rect 22152 12588 22158 12640
rect 26326 12588 26332 12640
rect 26384 12628 26390 12640
rect 26384 12600 26429 12628
rect 26384 12588 26390 12600
rect 27062 12588 27068 12640
rect 27120 12628 27126 12640
rect 27157 12631 27215 12637
rect 27157 12628 27169 12631
rect 27120 12600 27169 12628
rect 27120 12588 27126 12600
rect 27157 12597 27169 12600
rect 27203 12597 27215 12631
rect 27157 12591 27215 12597
rect 27522 12588 27528 12640
rect 27580 12628 27586 12640
rect 28074 12628 28080 12640
rect 27580 12600 28080 12628
rect 27580 12588 27586 12600
rect 28074 12588 28080 12600
rect 28132 12588 28138 12640
rect 1104 12538 28060 12560
rect 1104 12486 5442 12538
rect 5494 12486 5506 12538
rect 5558 12486 5570 12538
rect 5622 12486 5634 12538
rect 5686 12486 5698 12538
rect 5750 12486 14428 12538
rect 14480 12486 14492 12538
rect 14544 12486 14556 12538
rect 14608 12486 14620 12538
rect 14672 12486 14684 12538
rect 14736 12486 23413 12538
rect 23465 12486 23477 12538
rect 23529 12486 23541 12538
rect 23593 12486 23605 12538
rect 23657 12486 23669 12538
rect 23721 12486 28060 12538
rect 1104 12464 28060 12486
rect 1854 12384 1860 12436
rect 1912 12424 1918 12436
rect 2041 12427 2099 12433
rect 2041 12424 2053 12427
rect 1912 12396 2053 12424
rect 1912 12384 1918 12396
rect 2041 12393 2053 12396
rect 2087 12393 2099 12427
rect 2498 12424 2504 12436
rect 2459 12396 2504 12424
rect 2041 12387 2099 12393
rect 2498 12384 2504 12396
rect 2556 12384 2562 12436
rect 3418 12384 3424 12436
rect 3476 12424 3482 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 3476 12396 3801 12424
rect 3476 12384 3482 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 3970 12424 3976 12436
rect 3789 12387 3847 12393
rect 3896 12396 3976 12424
rect 2958 12316 2964 12368
rect 3016 12356 3022 12368
rect 3896 12356 3924 12396
rect 3970 12384 3976 12396
rect 4028 12384 4034 12436
rect 4338 12384 4344 12436
rect 4396 12424 4402 12436
rect 4522 12424 4528 12436
rect 4396 12396 4528 12424
rect 4396 12384 4402 12396
rect 4522 12384 4528 12396
rect 4580 12384 4586 12436
rect 7742 12424 7748 12436
rect 7703 12396 7748 12424
rect 7742 12384 7748 12396
rect 7800 12384 7806 12436
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 10321 12427 10379 12433
rect 10321 12424 10333 12427
rect 10100 12396 10333 12424
rect 10100 12384 10106 12396
rect 10321 12393 10333 12396
rect 10367 12393 10379 12427
rect 12986 12424 12992 12436
rect 10321 12387 10379 12393
rect 10419 12396 12992 12424
rect 3016 12328 3924 12356
rect 4249 12359 4307 12365
rect 3016 12316 3022 12328
rect 4249 12325 4261 12359
rect 4295 12325 4307 12359
rect 4249 12319 4307 12325
rect 2130 12248 2136 12300
rect 2188 12288 2194 12300
rect 2498 12288 2504 12300
rect 2188 12260 2504 12288
rect 2188 12248 2194 12260
rect 2498 12248 2504 12260
rect 2556 12248 2562 12300
rect 2682 12220 2688 12232
rect 2643 12192 2688 12220
rect 2682 12180 2688 12192
rect 2740 12180 2746 12232
rect 3418 12180 3424 12232
rect 3476 12220 3482 12232
rect 3973 12223 4031 12229
rect 3973 12220 3985 12223
rect 3476 12192 3985 12220
rect 3476 12180 3482 12192
rect 3973 12189 3985 12192
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 4120 12192 4165 12220
rect 4120 12180 4126 12192
rect 1670 12152 1676 12164
rect 1631 12124 1676 12152
rect 1670 12112 1676 12124
rect 1728 12112 1734 12164
rect 1857 12155 1915 12161
rect 1857 12121 1869 12155
rect 1903 12152 1915 12155
rect 2130 12152 2136 12164
rect 1903 12124 2136 12152
rect 1903 12121 1915 12124
rect 1857 12115 1915 12121
rect 2130 12112 2136 12124
rect 2188 12112 2194 12164
rect 3970 12044 3976 12096
rect 4028 12084 4034 12096
rect 4264 12084 4292 12319
rect 5718 12316 5724 12368
rect 5776 12356 5782 12368
rect 5994 12356 6000 12368
rect 5776 12328 6000 12356
rect 5776 12316 5782 12328
rect 5994 12316 6000 12328
rect 6052 12316 6058 12368
rect 6822 12316 6828 12368
rect 6880 12356 6886 12368
rect 8018 12356 8024 12368
rect 6880 12328 8024 12356
rect 6880 12316 6886 12328
rect 8018 12316 8024 12328
rect 8076 12316 8082 12368
rect 8938 12356 8944 12368
rect 8220 12328 8944 12356
rect 4982 12248 4988 12300
rect 5040 12288 5046 12300
rect 7377 12291 7435 12297
rect 5040 12260 5672 12288
rect 5040 12248 5046 12260
rect 4341 12223 4399 12229
rect 4341 12189 4353 12223
rect 4387 12220 4399 12223
rect 4706 12220 4712 12232
rect 4387 12192 4712 12220
rect 4387 12189 4399 12192
rect 4341 12183 4399 12189
rect 4706 12180 4712 12192
rect 4764 12180 4770 12232
rect 5350 12220 5356 12232
rect 5311 12192 5356 12220
rect 5350 12180 5356 12192
rect 5408 12180 5414 12232
rect 5644 12229 5672 12260
rect 6012 12260 6776 12288
rect 6012 12232 6040 12260
rect 5629 12223 5687 12229
rect 5629 12189 5641 12223
rect 5675 12189 5687 12223
rect 5629 12183 5687 12189
rect 5721 12223 5779 12229
rect 5721 12189 5733 12223
rect 5767 12220 5779 12223
rect 5994 12220 6000 12232
rect 5767 12192 6000 12220
rect 5767 12189 5779 12192
rect 5721 12183 5779 12189
rect 5994 12180 6000 12192
rect 6052 12180 6058 12232
rect 6362 12220 6368 12232
rect 6323 12192 6368 12220
rect 6362 12180 6368 12192
rect 6420 12180 6426 12232
rect 6638 12220 6644 12232
rect 6599 12192 6644 12220
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 6748 12229 6776 12260
rect 7377 12257 7389 12291
rect 7423 12288 7435 12291
rect 8220 12288 8248 12328
rect 8938 12316 8944 12328
rect 8996 12356 9002 12368
rect 9585 12359 9643 12365
rect 9585 12356 9597 12359
rect 8996 12328 9597 12356
rect 8996 12316 9002 12328
rect 9585 12325 9597 12328
rect 9631 12325 9643 12359
rect 9585 12319 9643 12325
rect 9766 12316 9772 12368
rect 9824 12356 9830 12368
rect 10419 12356 10447 12396
rect 12986 12384 12992 12396
rect 13044 12384 13050 12436
rect 13081 12427 13139 12433
rect 13081 12393 13093 12427
rect 13127 12424 13139 12427
rect 13262 12424 13268 12436
rect 13127 12396 13268 12424
rect 13127 12393 13139 12396
rect 13081 12387 13139 12393
rect 13262 12384 13268 12396
rect 13320 12384 13326 12436
rect 15657 12427 15715 12433
rect 14200 12396 15608 12424
rect 9824 12328 10447 12356
rect 9824 12316 9830 12328
rect 7423 12260 8248 12288
rect 8297 12291 8355 12297
rect 7423 12257 7435 12260
rect 7377 12251 7435 12257
rect 8297 12257 8309 12291
rect 8343 12288 8355 12291
rect 10594 12288 10600 12300
rect 8343 12260 10600 12288
rect 8343 12257 8355 12260
rect 8297 12251 8355 12257
rect 10594 12248 10600 12260
rect 10652 12248 10658 12300
rect 11698 12288 11704 12300
rect 11659 12260 11704 12288
rect 11698 12248 11704 12260
rect 11756 12248 11762 12300
rect 13262 12248 13268 12300
rect 13320 12288 13326 12300
rect 13446 12288 13452 12300
rect 13320 12260 13452 12288
rect 13320 12248 13326 12260
rect 13446 12248 13452 12260
rect 13504 12248 13510 12300
rect 6733 12223 6791 12229
rect 6733 12189 6745 12223
rect 6779 12189 6791 12223
rect 6733 12183 6791 12189
rect 7561 12223 7619 12229
rect 7561 12189 7573 12223
rect 7607 12189 7619 12223
rect 7561 12183 7619 12189
rect 8205 12223 8263 12229
rect 8205 12189 8217 12223
rect 8251 12220 8263 12223
rect 10318 12220 10324 12232
rect 8251 12192 10324 12220
rect 8251 12189 8263 12192
rect 8205 12183 8263 12189
rect 5534 12152 5540 12164
rect 5495 12124 5540 12152
rect 5534 12112 5540 12124
rect 5592 12152 5598 12164
rect 6549 12155 6607 12161
rect 6549 12152 6561 12155
rect 5592 12124 6561 12152
rect 5592 12112 5598 12124
rect 6549 12121 6561 12124
rect 6595 12121 6607 12155
rect 7576 12152 7604 12183
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 10502 12220 10508 12232
rect 10463 12192 10508 12220
rect 10502 12180 10508 12192
rect 10560 12180 10566 12232
rect 10781 12223 10839 12229
rect 10781 12220 10793 12223
rect 10612 12192 10793 12220
rect 6549 12115 6607 12121
rect 6932 12124 7604 12152
rect 5902 12084 5908 12096
rect 4028 12056 4292 12084
rect 5863 12056 5908 12084
rect 4028 12044 4034 12056
rect 5902 12044 5908 12056
rect 5960 12044 5966 12096
rect 6932 12093 6960 12124
rect 8294 12112 8300 12164
rect 8352 12152 8358 12164
rect 8846 12152 8852 12164
rect 8352 12124 8852 12152
rect 8352 12112 8358 12124
rect 8846 12112 8852 12124
rect 8904 12152 8910 12164
rect 9401 12155 9459 12161
rect 9401 12152 9413 12155
rect 8904 12124 9413 12152
rect 8904 12112 8910 12124
rect 9401 12121 9413 12124
rect 9447 12121 9459 12155
rect 9401 12115 9459 12121
rect 9582 12112 9588 12164
rect 9640 12152 9646 12164
rect 10612 12152 10640 12192
rect 10781 12189 10793 12192
rect 10827 12189 10839 12223
rect 11968 12223 12026 12229
rect 11968 12220 11980 12223
rect 10781 12183 10839 12189
rect 11900 12192 11980 12220
rect 9640 12124 10640 12152
rect 10689 12155 10747 12161
rect 9640 12112 9646 12124
rect 10689 12121 10701 12155
rect 10735 12152 10747 12155
rect 11606 12152 11612 12164
rect 10735 12124 11612 12152
rect 10735 12121 10747 12124
rect 10689 12115 10747 12121
rect 11606 12112 11612 12124
rect 11664 12112 11670 12164
rect 11900 12096 11928 12192
rect 11968 12189 11980 12192
rect 12014 12189 12026 12223
rect 11968 12183 12026 12189
rect 14200 12152 14228 12396
rect 15580 12356 15608 12396
rect 15657 12393 15669 12427
rect 15703 12424 15715 12427
rect 15930 12424 15936 12436
rect 15703 12396 15936 12424
rect 15703 12393 15715 12396
rect 15657 12387 15715 12393
rect 15930 12384 15936 12396
rect 15988 12384 15994 12436
rect 17589 12427 17647 12433
rect 16224 12396 17540 12424
rect 16224 12356 16252 12396
rect 15580 12328 16252 12356
rect 17512 12356 17540 12396
rect 17589 12393 17601 12427
rect 17635 12424 17647 12427
rect 18046 12424 18052 12436
rect 17635 12396 18052 12424
rect 17635 12393 17647 12396
rect 17589 12387 17647 12393
rect 18046 12384 18052 12396
rect 18104 12384 18110 12436
rect 18417 12427 18475 12433
rect 18417 12393 18429 12427
rect 18463 12424 18475 12427
rect 21542 12424 21548 12436
rect 18463 12396 21128 12424
rect 21503 12396 21548 12424
rect 18463 12393 18475 12396
rect 18417 12387 18475 12393
rect 20070 12356 20076 12368
rect 17512 12328 20076 12356
rect 20070 12316 20076 12328
rect 20128 12316 20134 12368
rect 21100 12356 21128 12396
rect 21542 12384 21548 12396
rect 21600 12384 21606 12436
rect 23290 12424 23296 12436
rect 23251 12396 23296 12424
rect 23290 12384 23296 12396
rect 23348 12384 23354 12436
rect 25409 12427 25467 12433
rect 23400 12396 25351 12424
rect 22278 12356 22284 12368
rect 21100 12328 22284 12356
rect 22278 12316 22284 12328
rect 22336 12316 22342 12368
rect 22922 12316 22928 12368
rect 22980 12356 22986 12368
rect 23400 12356 23428 12396
rect 22980 12328 23428 12356
rect 23661 12359 23719 12365
rect 22980 12316 22986 12328
rect 23661 12325 23673 12359
rect 23707 12356 23719 12359
rect 24118 12356 24124 12368
rect 23707 12328 24124 12356
rect 23707 12325 23719 12328
rect 23661 12319 23719 12325
rect 24118 12316 24124 12328
rect 24176 12316 24182 12368
rect 25323 12356 25351 12396
rect 25409 12393 25421 12427
rect 25455 12424 25467 12427
rect 26326 12424 26332 12436
rect 25455 12396 26332 12424
rect 25455 12393 25467 12396
rect 25409 12387 25467 12393
rect 26326 12384 26332 12396
rect 26384 12384 26390 12436
rect 27614 12384 27620 12436
rect 27672 12424 27678 12436
rect 27890 12424 27896 12436
rect 27672 12396 27896 12424
rect 27672 12384 27678 12396
rect 27890 12384 27896 12396
rect 27948 12384 27954 12436
rect 25323 12328 25544 12356
rect 25516 12300 25544 12328
rect 18046 12248 18052 12300
rect 18104 12288 18110 12300
rect 19058 12288 19064 12300
rect 18104 12260 19064 12288
rect 18104 12248 18110 12260
rect 18248 12229 18276 12260
rect 19058 12248 19064 12260
rect 19116 12248 19122 12300
rect 19702 12288 19708 12300
rect 19663 12260 19708 12288
rect 19702 12248 19708 12260
rect 19760 12248 19766 12300
rect 21174 12248 21180 12300
rect 21232 12288 21238 12300
rect 23753 12291 23811 12297
rect 21232 12260 22324 12288
rect 21232 12248 21238 12260
rect 22296 12232 22324 12260
rect 23753 12257 23765 12291
rect 23799 12288 23811 12291
rect 24026 12288 24032 12300
rect 23799 12260 24032 12288
rect 23799 12257 23811 12260
rect 23753 12251 23811 12257
rect 24026 12248 24032 12260
rect 24084 12248 24090 12300
rect 25498 12288 25504 12300
rect 25411 12260 25504 12288
rect 25498 12248 25504 12260
rect 25556 12248 25562 12300
rect 25958 12288 25964 12300
rect 25919 12260 25964 12288
rect 25958 12248 25964 12260
rect 26016 12248 26022 12300
rect 27430 12248 27436 12300
rect 27488 12288 27494 12300
rect 27614 12288 27620 12300
rect 27488 12260 27620 12288
rect 27488 12248 27494 12260
rect 27614 12248 27620 12260
rect 27672 12248 27678 12300
rect 14277 12223 14335 12229
rect 14277 12189 14289 12223
rect 14323 12220 14335 12223
rect 16209 12223 16267 12229
rect 16209 12220 16221 12223
rect 14323 12192 16221 12220
rect 14323 12189 14335 12192
rect 14277 12183 14335 12189
rect 16209 12189 16221 12192
rect 16255 12220 16267 12223
rect 18233 12223 18291 12229
rect 16255 12192 16712 12220
rect 16255 12189 16267 12192
rect 16209 12183 16267 12189
rect 16684 12164 16712 12192
rect 18233 12189 18245 12223
rect 18279 12189 18291 12223
rect 19337 12223 19395 12229
rect 19337 12220 19349 12223
rect 18233 12183 18291 12189
rect 18340 12192 19349 12220
rect 14522 12155 14580 12161
rect 14522 12152 14534 12155
rect 14200 12124 14534 12152
rect 14522 12121 14534 12124
rect 14568 12121 14580 12155
rect 14522 12115 14580 12121
rect 15930 12112 15936 12164
rect 15988 12152 15994 12164
rect 16454 12155 16512 12161
rect 16454 12152 16466 12155
rect 15988 12124 16466 12152
rect 15988 12112 15994 12124
rect 16454 12121 16466 12124
rect 16500 12121 16512 12155
rect 16454 12115 16512 12121
rect 16666 12112 16672 12164
rect 16724 12112 16730 12164
rect 17770 12112 17776 12164
rect 17828 12152 17834 12164
rect 18049 12155 18107 12161
rect 18049 12152 18061 12155
rect 17828 12124 18061 12152
rect 17828 12112 17834 12124
rect 18049 12121 18061 12124
rect 18095 12152 18107 12155
rect 18340 12152 18368 12192
rect 19337 12189 19349 12192
rect 19383 12189 19395 12223
rect 19337 12183 19395 12189
rect 20165 12223 20223 12229
rect 20165 12189 20177 12223
rect 20211 12220 20223 12223
rect 21910 12220 21916 12232
rect 20211 12192 21916 12220
rect 20211 12189 20223 12192
rect 20165 12183 20223 12189
rect 21910 12180 21916 12192
rect 21968 12180 21974 12232
rect 22051 12223 22109 12229
rect 22051 12189 22063 12223
rect 22097 12189 22109 12223
rect 22278 12220 22284 12232
rect 22239 12192 22284 12220
rect 22051 12183 22109 12189
rect 18095 12124 18368 12152
rect 18095 12121 18107 12124
rect 18049 12115 18107 12121
rect 18598 12112 18604 12164
rect 18656 12152 18662 12164
rect 19150 12152 19156 12164
rect 18656 12124 19156 12152
rect 18656 12112 18662 12124
rect 19150 12112 19156 12124
rect 19208 12112 19214 12164
rect 19521 12155 19579 12161
rect 19521 12121 19533 12155
rect 19567 12152 19579 12155
rect 20070 12152 20076 12164
rect 19567 12124 20076 12152
rect 19567 12121 19579 12124
rect 19521 12115 19579 12121
rect 20070 12112 20076 12124
rect 20128 12112 20134 12164
rect 20432 12155 20490 12161
rect 20432 12121 20444 12155
rect 20478 12152 20490 12155
rect 20530 12152 20536 12164
rect 20478 12124 20536 12152
rect 20478 12121 20490 12124
rect 20432 12115 20490 12121
rect 20530 12112 20536 12124
rect 20588 12112 20594 12164
rect 20622 12112 20628 12164
rect 20680 12152 20686 12164
rect 20680 12124 21956 12152
rect 20680 12112 20686 12124
rect 6917 12087 6975 12093
rect 6917 12053 6929 12087
rect 6963 12053 6975 12087
rect 6917 12047 6975 12053
rect 8018 12044 8024 12096
rect 8076 12084 8082 12096
rect 8386 12084 8392 12096
rect 8076 12056 8392 12084
rect 8076 12044 8082 12056
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 11882 12044 11888 12096
rect 11940 12044 11946 12096
rect 12526 12044 12532 12096
rect 12584 12084 12590 12096
rect 12802 12084 12808 12096
rect 12584 12056 12808 12084
rect 12584 12044 12590 12056
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 12894 12044 12900 12096
rect 12952 12084 12958 12096
rect 13722 12084 13728 12096
rect 12952 12056 13728 12084
rect 12952 12044 12958 12056
rect 13722 12044 13728 12056
rect 13780 12044 13786 12096
rect 13814 12044 13820 12096
rect 13872 12084 13878 12096
rect 15838 12084 15844 12096
rect 13872 12056 15844 12084
rect 13872 12044 13878 12056
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 16206 12044 16212 12096
rect 16264 12084 16270 12096
rect 17678 12084 17684 12096
rect 16264 12056 17684 12084
rect 16264 12044 16270 12056
rect 17678 12044 17684 12056
rect 17736 12044 17742 12096
rect 21928 12084 21956 12124
rect 22066 12084 22094 12183
rect 22278 12180 22284 12192
rect 22336 12180 22342 12232
rect 23477 12223 23535 12229
rect 23477 12189 23489 12223
rect 23523 12220 23535 12223
rect 23842 12220 23848 12232
rect 23523 12192 23848 12220
rect 23523 12189 23535 12192
rect 23477 12183 23535 12189
rect 23842 12180 23848 12192
rect 23900 12180 23906 12232
rect 24394 12180 24400 12232
rect 24452 12180 24458 12232
rect 24581 12223 24639 12229
rect 24581 12189 24593 12223
rect 24627 12220 24639 12223
rect 25038 12220 25044 12232
rect 24627 12192 25044 12220
rect 24627 12189 24639 12192
rect 24581 12183 24639 12189
rect 25038 12180 25044 12192
rect 25096 12180 25102 12232
rect 25225 12223 25283 12229
rect 25225 12189 25237 12223
rect 25271 12220 25283 12223
rect 25406 12220 25412 12232
rect 25271 12192 25412 12220
rect 25271 12189 25283 12192
rect 25225 12183 25283 12189
rect 25406 12180 25412 12192
rect 25464 12180 25470 12232
rect 26234 12229 26240 12232
rect 26228 12183 26240 12229
rect 26292 12220 26298 12232
rect 26292 12192 26328 12220
rect 26234 12180 26240 12183
rect 26292 12180 26298 12192
rect 24412 12152 24440 12180
rect 26602 12152 26608 12164
rect 24412 12124 26608 12152
rect 26602 12112 26608 12124
rect 26660 12152 26666 12164
rect 26660 12124 27384 12152
rect 26660 12112 26666 12124
rect 23106 12084 23112 12096
rect 21928 12056 23112 12084
rect 23106 12044 23112 12056
rect 23164 12044 23170 12096
rect 24026 12044 24032 12096
rect 24084 12084 24090 12096
rect 24397 12087 24455 12093
rect 24397 12084 24409 12087
rect 24084 12056 24409 12084
rect 24084 12044 24090 12056
rect 24397 12053 24409 12056
rect 24443 12053 24455 12087
rect 24397 12047 24455 12053
rect 25041 12087 25099 12093
rect 25041 12053 25053 12087
rect 25087 12084 25099 12087
rect 25130 12084 25136 12096
rect 25087 12056 25136 12084
rect 25087 12053 25099 12056
rect 25041 12047 25099 12053
rect 25130 12044 25136 12056
rect 25188 12044 25194 12096
rect 27356 12093 27384 12124
rect 27341 12087 27399 12093
rect 27341 12053 27353 12087
rect 27387 12053 27399 12087
rect 27341 12047 27399 12053
rect 27430 12044 27436 12096
rect 27488 12084 27494 12096
rect 28074 12084 28080 12096
rect 27488 12056 28080 12084
rect 27488 12044 27494 12056
rect 28074 12044 28080 12056
rect 28132 12044 28138 12096
rect 1104 11994 28060 12016
rect 1104 11942 9935 11994
rect 9987 11942 9999 11994
rect 10051 11942 10063 11994
rect 10115 11942 10127 11994
rect 10179 11942 10191 11994
rect 10243 11942 18920 11994
rect 18972 11942 18984 11994
rect 19036 11942 19048 11994
rect 19100 11942 19112 11994
rect 19164 11942 19176 11994
rect 19228 11942 28060 11994
rect 1104 11920 28060 11942
rect 1670 11840 1676 11892
rect 1728 11880 1734 11892
rect 2777 11883 2835 11889
rect 2777 11880 2789 11883
rect 1728 11852 2789 11880
rect 1728 11840 1734 11852
rect 2777 11849 2789 11852
rect 2823 11849 2835 11883
rect 2777 11843 2835 11849
rect 3602 11840 3608 11892
rect 3660 11880 3666 11892
rect 3789 11883 3847 11889
rect 3789 11880 3801 11883
rect 3660 11852 3801 11880
rect 3660 11840 3666 11852
rect 3789 11849 3801 11852
rect 3835 11849 3847 11883
rect 3789 11843 3847 11849
rect 5258 11840 5264 11892
rect 5316 11840 5322 11892
rect 6270 11840 6276 11892
rect 6328 11880 6334 11892
rect 6733 11883 6791 11889
rect 6733 11880 6745 11883
rect 6328 11852 6745 11880
rect 6328 11840 6334 11852
rect 6733 11849 6745 11852
rect 6779 11849 6791 11883
rect 6733 11843 6791 11849
rect 7006 11840 7012 11892
rect 7064 11880 7070 11892
rect 7064 11852 8984 11880
rect 7064 11840 7070 11852
rect 2406 11772 2412 11824
rect 2464 11812 2470 11824
rect 4430 11812 4436 11824
rect 2464 11784 3372 11812
rect 2464 11772 2470 11784
rect 1026 11704 1032 11756
rect 1084 11744 1090 11756
rect 1670 11744 1676 11756
rect 1084 11716 1676 11744
rect 1084 11704 1090 11716
rect 1670 11704 1676 11716
rect 1728 11704 1734 11756
rect 2038 11744 2044 11756
rect 1999 11716 2044 11744
rect 2038 11704 2044 11716
rect 2096 11704 2102 11756
rect 2774 11704 2780 11756
rect 2832 11744 2838 11756
rect 3344 11753 3372 11784
rect 4080 11784 4436 11812
rect 2961 11747 3019 11753
rect 2961 11744 2973 11747
rect 2832 11716 2973 11744
rect 2832 11704 2838 11716
rect 2961 11713 2973 11716
rect 3007 11713 3019 11747
rect 2961 11707 3019 11713
rect 3053 11747 3111 11753
rect 3053 11713 3065 11747
rect 3099 11713 3111 11747
rect 3053 11707 3111 11713
rect 3329 11747 3387 11753
rect 3329 11713 3341 11747
rect 3375 11713 3387 11747
rect 3329 11707 3387 11713
rect 3068 11676 3096 11707
rect 3418 11704 3424 11756
rect 3476 11744 3482 11756
rect 4080 11753 4108 11784
rect 4430 11772 4436 11784
rect 4488 11772 4494 11824
rect 5276 11812 5304 11840
rect 5353 11815 5411 11821
rect 5353 11812 5365 11815
rect 5276 11784 5365 11812
rect 5353 11781 5365 11784
rect 5399 11781 5411 11815
rect 5353 11775 5411 11781
rect 6362 11772 6368 11824
rect 6420 11812 6426 11824
rect 6420 11784 6684 11812
rect 6420 11772 6426 11784
rect 3973 11747 4031 11753
rect 3973 11744 3985 11747
rect 3476 11716 3985 11744
rect 3476 11704 3482 11716
rect 3973 11713 3985 11716
rect 4019 11713 4031 11747
rect 3973 11707 4031 11713
rect 4065 11747 4123 11753
rect 4065 11713 4077 11747
rect 4111 11713 4123 11747
rect 4338 11744 4344 11756
rect 4299 11716 4344 11744
rect 4065 11707 4123 11713
rect 4338 11704 4344 11716
rect 4396 11704 4402 11756
rect 5074 11744 5080 11756
rect 5035 11716 5080 11744
rect 5074 11704 5080 11716
rect 5132 11704 5138 11756
rect 5261 11747 5319 11753
rect 5261 11713 5273 11747
rect 5307 11713 5319 11747
rect 5261 11707 5319 11713
rect 5445 11747 5503 11753
rect 5445 11713 5457 11747
rect 5491 11713 5503 11747
rect 5445 11707 5503 11713
rect 3878 11676 3884 11688
rect 3068 11648 3884 11676
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 4430 11636 4436 11688
rect 4488 11676 4494 11688
rect 4798 11676 4804 11688
rect 4488 11648 4804 11676
rect 4488 11636 4494 11648
rect 4798 11636 4804 11648
rect 4856 11636 4862 11688
rect 5276 11676 5304 11707
rect 5350 11676 5356 11688
rect 5276 11648 5356 11676
rect 5350 11636 5356 11648
rect 5408 11636 5414 11688
rect 5460 11676 5488 11707
rect 5902 11704 5908 11756
rect 5960 11744 5966 11756
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 5960 11716 6561 11744
rect 5960 11704 5966 11716
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 6656 11744 6684 11784
rect 7650 11772 7656 11824
rect 7708 11812 7714 11824
rect 7990 11815 8048 11821
rect 7990 11812 8002 11815
rect 7708 11784 8002 11812
rect 7708 11772 7714 11784
rect 7990 11781 8002 11784
rect 8036 11781 8048 11815
rect 8956 11812 8984 11852
rect 9030 11840 9036 11892
rect 9088 11880 9094 11892
rect 9125 11883 9183 11889
rect 9125 11880 9137 11883
rect 9088 11852 9137 11880
rect 9088 11840 9094 11852
rect 9125 11849 9137 11852
rect 9171 11880 9183 11883
rect 9582 11880 9588 11892
rect 9171 11852 9588 11880
rect 9171 11849 9183 11852
rect 9125 11843 9183 11849
rect 9582 11840 9588 11852
rect 9640 11840 9646 11892
rect 10318 11840 10324 11892
rect 10376 11880 10382 11892
rect 10965 11883 11023 11889
rect 10965 11880 10977 11883
rect 10376 11852 10977 11880
rect 10376 11840 10382 11852
rect 10965 11849 10977 11852
rect 11011 11849 11023 11883
rect 10965 11843 11023 11849
rect 11974 11840 11980 11892
rect 12032 11880 12038 11892
rect 12253 11883 12311 11889
rect 12253 11880 12265 11883
rect 12032 11852 12265 11880
rect 12032 11840 12038 11852
rect 12253 11849 12265 11852
rect 12299 11849 12311 11883
rect 12253 11843 12311 11849
rect 13648 11852 14412 11880
rect 11885 11815 11943 11821
rect 11885 11812 11897 11815
rect 8956 11784 11897 11812
rect 7990 11775 8048 11781
rect 11885 11781 11897 11784
rect 11931 11812 11943 11815
rect 13648 11812 13676 11852
rect 11931 11784 13676 11812
rect 14277 11815 14335 11821
rect 11931 11781 11943 11784
rect 11885 11775 11943 11781
rect 14277 11781 14289 11815
rect 14323 11781 14335 11815
rect 14384 11812 14412 11852
rect 14458 11840 14464 11892
rect 14516 11889 14522 11892
rect 14516 11883 14535 11889
rect 14523 11849 14535 11883
rect 14642 11880 14648 11892
rect 14603 11852 14648 11880
rect 14516 11843 14535 11849
rect 14516 11840 14522 11843
rect 14642 11840 14648 11852
rect 14700 11840 14706 11892
rect 14752 11852 16160 11880
rect 14752 11812 14780 11852
rect 14384 11784 14780 11812
rect 15565 11815 15623 11821
rect 14277 11775 14335 11781
rect 15565 11781 15577 11815
rect 15611 11781 15623 11815
rect 15565 11775 15623 11781
rect 15781 11815 15839 11821
rect 15781 11781 15793 11815
rect 15827 11812 15839 11815
rect 15930 11812 15936 11824
rect 15827 11784 15936 11812
rect 15827 11781 15839 11784
rect 15781 11775 15839 11781
rect 6656 11716 8800 11744
rect 6549 11707 6607 11713
rect 5994 11676 6000 11688
rect 5460 11648 6000 11676
rect 5994 11636 6000 11648
rect 6052 11636 6058 11688
rect 6365 11679 6423 11685
rect 6365 11645 6377 11679
rect 6411 11645 6423 11679
rect 6365 11639 6423 11645
rect 3237 11611 3295 11617
rect 3237 11577 3249 11611
rect 3283 11608 3295 11611
rect 3970 11608 3976 11620
rect 3283 11580 3976 11608
rect 3283 11577 3295 11580
rect 3237 11571 3295 11577
rect 3970 11568 3976 11580
rect 4028 11608 4034 11620
rect 4249 11611 4307 11617
rect 4249 11608 4261 11611
rect 4028 11580 4261 11608
rect 4028 11568 4034 11580
rect 4249 11577 4261 11580
rect 4295 11577 4307 11611
rect 4249 11571 4307 11577
rect 5718 11568 5724 11620
rect 5776 11608 5782 11620
rect 5776 11580 6316 11608
rect 5776 11568 5782 11580
rect 6288 11552 6316 11580
rect 1854 11540 1860 11552
rect 1815 11512 1860 11540
rect 1854 11500 1860 11512
rect 1912 11500 1918 11552
rect 5629 11543 5687 11549
rect 5629 11509 5641 11543
rect 5675 11540 5687 11543
rect 5902 11540 5908 11552
rect 5675 11512 5908 11540
rect 5675 11509 5687 11512
rect 5629 11503 5687 11509
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 6270 11500 6276 11552
rect 6328 11500 6334 11552
rect 6380 11540 6408 11639
rect 6638 11636 6644 11688
rect 6696 11676 6702 11688
rect 7745 11679 7803 11685
rect 7745 11676 7757 11679
rect 6696 11648 7757 11676
rect 6696 11636 6702 11648
rect 7745 11645 7757 11648
rect 7791 11645 7803 11679
rect 8772 11676 8800 11716
rect 9030 11704 9036 11756
rect 9088 11744 9094 11756
rect 9398 11744 9404 11756
rect 9088 11716 9404 11744
rect 9088 11704 9094 11716
rect 9398 11704 9404 11716
rect 9456 11704 9462 11756
rect 9841 11747 9899 11753
rect 9841 11744 9853 11747
rect 9508 11716 9853 11744
rect 9508 11676 9536 11716
rect 9841 11713 9853 11716
rect 9887 11713 9899 11747
rect 9841 11707 9899 11713
rect 12069 11747 12127 11753
rect 12069 11713 12081 11747
rect 12115 11744 12127 11747
rect 12710 11744 12716 11756
rect 12115 11716 12434 11744
rect 12671 11716 12716 11744
rect 12115 11713 12127 11716
rect 12069 11707 12127 11713
rect 8772 11648 9536 11676
rect 9585 11679 9643 11685
rect 7745 11639 7803 11645
rect 9585 11645 9597 11679
rect 9631 11645 9643 11679
rect 9585 11639 9643 11645
rect 8386 11540 8392 11552
rect 6380 11512 8392 11540
rect 8386 11500 8392 11512
rect 8444 11500 8450 11552
rect 9600 11540 9628 11639
rect 11698 11540 11704 11552
rect 9600 11512 11704 11540
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 11882 11500 11888 11552
rect 11940 11540 11946 11552
rect 12158 11540 12164 11552
rect 11940 11512 12164 11540
rect 11940 11500 11946 11512
rect 12158 11500 12164 11512
rect 12216 11500 12222 11552
rect 12406 11540 12434 11716
rect 12710 11704 12716 11716
rect 12768 11704 12774 11756
rect 12986 11744 12992 11756
rect 12947 11716 12992 11744
rect 12986 11704 12992 11716
rect 13044 11704 13050 11756
rect 13078 11704 13084 11756
rect 13136 11744 13142 11756
rect 13541 11747 13599 11753
rect 13541 11744 13553 11747
rect 13136 11716 13553 11744
rect 13136 11704 13142 11716
rect 13541 11713 13553 11716
rect 13587 11744 13599 11747
rect 14292 11744 14320 11775
rect 15580 11744 15608 11775
rect 15930 11772 15936 11784
rect 15988 11772 15994 11824
rect 13587 11716 15608 11744
rect 13587 11713 13599 11716
rect 13541 11707 13599 11713
rect 13446 11636 13452 11688
rect 13504 11676 13510 11688
rect 13504 11648 14504 11676
rect 13504 11636 13510 11648
rect 12989 11611 13047 11617
rect 12989 11577 13001 11611
rect 13035 11608 13047 11611
rect 13078 11608 13084 11620
rect 13035 11580 13084 11608
rect 13035 11577 13047 11580
rect 12989 11571 13047 11577
rect 13078 11568 13084 11580
rect 13136 11568 13142 11620
rect 13722 11608 13728 11620
rect 13683 11580 13728 11608
rect 13722 11568 13728 11580
rect 13780 11568 13786 11620
rect 12526 11540 12532 11552
rect 12406 11512 12532 11540
rect 12526 11500 12532 11512
rect 12584 11500 12590 11552
rect 12802 11500 12808 11552
rect 12860 11540 12866 11552
rect 13740 11540 13768 11568
rect 12860 11512 13768 11540
rect 12860 11500 12866 11512
rect 13814 11500 13820 11552
rect 13872 11540 13878 11552
rect 14274 11540 14280 11552
rect 13872 11512 14280 11540
rect 13872 11500 13878 11512
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 14476 11549 14504 11648
rect 15194 11636 15200 11688
rect 15252 11676 15258 11688
rect 16132 11676 16160 11852
rect 17310 11840 17316 11892
rect 17368 11880 17374 11892
rect 17494 11880 17500 11892
rect 17368 11852 17500 11880
rect 17368 11840 17374 11852
rect 17494 11840 17500 11852
rect 17552 11840 17558 11892
rect 18598 11880 18604 11892
rect 18559 11852 18604 11880
rect 18598 11840 18604 11852
rect 18656 11840 18662 11892
rect 19794 11880 19800 11892
rect 19536 11852 19800 11880
rect 18233 11815 18291 11821
rect 18233 11812 18245 11815
rect 16960 11784 18245 11812
rect 16960 11753 16988 11784
rect 18233 11781 18245 11784
rect 18279 11812 18291 11815
rect 19426 11812 19432 11824
rect 18279 11784 19432 11812
rect 18279 11781 18291 11784
rect 18233 11775 18291 11781
rect 19426 11772 19432 11784
rect 19484 11812 19490 11824
rect 19536 11821 19564 11852
rect 19794 11840 19800 11852
rect 19852 11840 19858 11892
rect 20070 11840 20076 11892
rect 20128 11880 20134 11892
rect 20346 11880 20352 11892
rect 20128 11852 20352 11880
rect 20128 11840 20134 11852
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 20990 11840 20996 11892
rect 21048 11880 21054 11892
rect 22002 11880 22008 11892
rect 21048 11852 22008 11880
rect 21048 11840 21054 11852
rect 22002 11840 22008 11852
rect 22060 11880 22066 11892
rect 23290 11880 23296 11892
rect 22060 11852 23296 11880
rect 22060 11840 22066 11852
rect 23290 11840 23296 11852
rect 23348 11840 23354 11892
rect 23934 11840 23940 11892
rect 23992 11880 23998 11892
rect 24029 11883 24087 11889
rect 24029 11880 24041 11883
rect 23992 11852 24041 11880
rect 23992 11840 23998 11852
rect 24029 11849 24041 11852
rect 24075 11849 24087 11883
rect 24029 11843 24087 11849
rect 25498 11840 25504 11892
rect 25556 11880 25562 11892
rect 26421 11883 26479 11889
rect 26421 11880 26433 11883
rect 25556 11852 26433 11880
rect 25556 11840 25562 11852
rect 26421 11849 26433 11852
rect 26467 11849 26479 11883
rect 26421 11843 26479 11849
rect 26602 11840 26608 11892
rect 26660 11880 26666 11892
rect 27338 11880 27344 11892
rect 26660 11852 27344 11880
rect 26660 11840 26666 11852
rect 27338 11840 27344 11852
rect 27396 11840 27402 11892
rect 19521 11815 19579 11821
rect 19521 11812 19533 11815
rect 19484 11784 19533 11812
rect 19484 11772 19490 11784
rect 19521 11781 19533 11784
rect 19567 11781 19579 11815
rect 21174 11812 21180 11824
rect 19521 11775 19579 11781
rect 19812 11784 21180 11812
rect 16945 11747 17003 11753
rect 16945 11713 16957 11747
rect 16991 11713 17003 11747
rect 16945 11707 17003 11713
rect 17221 11747 17279 11753
rect 17221 11713 17233 11747
rect 17267 11744 17279 11747
rect 17770 11744 17776 11756
rect 17267 11716 17776 11744
rect 17267 11713 17279 11716
rect 17221 11707 17279 11713
rect 17770 11704 17776 11716
rect 17828 11704 17834 11756
rect 18417 11747 18475 11753
rect 18417 11713 18429 11747
rect 18463 11744 18475 11747
rect 18874 11744 18880 11756
rect 18463 11716 18880 11744
rect 18463 11713 18475 11716
rect 18417 11707 18475 11713
rect 18874 11704 18880 11716
rect 18932 11704 18938 11756
rect 19150 11704 19156 11756
rect 19208 11744 19214 11756
rect 19812 11744 19840 11784
rect 21174 11772 21180 11784
rect 21232 11772 21238 11824
rect 21928 11784 23704 11812
rect 21928 11753 21956 11784
rect 19208 11716 19840 11744
rect 20901 11747 20959 11753
rect 19208 11704 19214 11716
rect 20901 11713 20913 11747
rect 20947 11713 20959 11747
rect 20901 11707 20959 11713
rect 21913 11747 21971 11753
rect 21913 11713 21925 11747
rect 21959 11713 21971 11747
rect 21913 11707 21971 11713
rect 19705 11679 19763 11685
rect 19705 11676 19717 11679
rect 15252 11648 16068 11676
rect 16132 11648 19717 11676
rect 15252 11636 15258 11648
rect 15838 11568 15844 11620
rect 15896 11608 15902 11620
rect 15933 11611 15991 11617
rect 15933 11608 15945 11611
rect 15896 11580 15945 11608
rect 15896 11568 15902 11580
rect 15933 11577 15945 11580
rect 15979 11577 15991 11611
rect 15933 11571 15991 11577
rect 14461 11543 14519 11549
rect 14461 11509 14473 11543
rect 14507 11540 14519 11543
rect 15286 11540 15292 11552
rect 14507 11512 15292 11540
rect 14507 11509 14519 11512
rect 14461 11503 14519 11509
rect 15286 11500 15292 11512
rect 15344 11540 15350 11552
rect 15749 11543 15807 11549
rect 15749 11540 15761 11543
rect 15344 11512 15761 11540
rect 15344 11500 15350 11512
rect 15749 11509 15761 11512
rect 15795 11509 15807 11543
rect 16040 11540 16068 11648
rect 19705 11645 19717 11648
rect 19751 11676 19763 11679
rect 19794 11676 19800 11688
rect 19751 11648 19800 11676
rect 19751 11645 19763 11648
rect 19705 11639 19763 11645
rect 19794 11636 19800 11648
rect 19852 11636 19858 11688
rect 20916 11676 20944 11707
rect 22002 11704 22008 11756
rect 22060 11744 22066 11756
rect 22097 11747 22155 11753
rect 22097 11744 22109 11747
rect 22060 11716 22109 11744
rect 22060 11704 22066 11716
rect 22097 11713 22109 11716
rect 22143 11713 22155 11747
rect 22097 11707 22155 11713
rect 22189 11747 22247 11753
rect 22189 11713 22201 11747
rect 22235 11713 22247 11747
rect 22189 11707 22247 11713
rect 21174 11676 21180 11688
rect 19904 11648 20760 11676
rect 20916 11648 21180 11676
rect 19518 11568 19524 11620
rect 19576 11608 19582 11620
rect 19904 11608 19932 11648
rect 20272 11620 20300 11648
rect 19576 11580 19932 11608
rect 19576 11568 19582 11580
rect 20254 11568 20260 11620
rect 20312 11568 20318 11620
rect 20622 11608 20628 11620
rect 20461 11580 20628 11608
rect 20461 11540 20489 11580
rect 20622 11568 20628 11580
rect 20680 11568 20686 11620
rect 20732 11608 20760 11648
rect 21174 11636 21180 11648
rect 21232 11636 21238 11688
rect 21634 11636 21640 11688
rect 21692 11676 21698 11688
rect 22204 11676 22232 11707
rect 22278 11704 22284 11756
rect 22336 11744 22342 11756
rect 22336 11716 22381 11744
rect 22336 11704 22342 11716
rect 23106 11704 23112 11756
rect 23164 11744 23170 11756
rect 23293 11747 23351 11753
rect 23293 11744 23305 11747
rect 23164 11716 23305 11744
rect 23164 11704 23170 11716
rect 23293 11713 23305 11716
rect 23339 11713 23351 11747
rect 23293 11707 23351 11713
rect 21692 11648 22232 11676
rect 23676 11676 23704 11784
rect 23750 11772 23756 11824
rect 23808 11812 23814 11824
rect 24762 11812 24768 11824
rect 23808 11784 24768 11812
rect 23808 11772 23814 11784
rect 24762 11772 24768 11784
rect 24820 11812 24826 11824
rect 24820 11784 25084 11812
rect 24820 11772 24826 11784
rect 24210 11744 24216 11756
rect 24171 11716 24216 11744
rect 24210 11704 24216 11716
rect 24268 11704 24274 11756
rect 25056 11753 25084 11784
rect 25041 11747 25099 11753
rect 25041 11713 25053 11747
rect 25087 11713 25099 11747
rect 25041 11707 25099 11713
rect 25130 11704 25136 11756
rect 25188 11744 25194 11756
rect 25297 11747 25355 11753
rect 25297 11744 25309 11747
rect 25188 11716 25309 11744
rect 25188 11704 25194 11716
rect 25297 11713 25309 11716
rect 25343 11713 25355 11747
rect 25297 11707 25355 11713
rect 25590 11704 25596 11756
rect 25648 11744 25654 11756
rect 26694 11744 26700 11756
rect 25648 11716 26700 11744
rect 25648 11704 25654 11716
rect 26694 11704 26700 11716
rect 26752 11704 26758 11756
rect 27062 11744 27068 11756
rect 27023 11716 27068 11744
rect 27062 11704 27068 11716
rect 27120 11704 27126 11756
rect 24489 11679 24547 11685
rect 24489 11676 24501 11679
rect 23676 11648 24501 11676
rect 21692 11636 21698 11648
rect 24489 11645 24501 11648
rect 24535 11676 24547 11679
rect 24670 11676 24676 11688
rect 24535 11648 24676 11676
rect 24535 11645 24547 11648
rect 24489 11639 24547 11645
rect 24670 11636 24676 11648
rect 24728 11636 24734 11688
rect 22465 11611 22523 11617
rect 22465 11608 22477 11611
rect 20732 11580 22477 11608
rect 22465 11577 22477 11580
rect 22511 11577 22523 11611
rect 27246 11608 27252 11620
rect 27207 11580 27252 11608
rect 22465 11571 22523 11577
rect 27246 11568 27252 11580
rect 27304 11568 27310 11620
rect 16040 11512 20489 11540
rect 15749 11503 15807 11509
rect 20530 11500 20536 11552
rect 20588 11540 20594 11552
rect 20717 11543 20775 11549
rect 20717 11540 20729 11543
rect 20588 11512 20729 11540
rect 20588 11500 20594 11512
rect 20717 11509 20729 11512
rect 20763 11509 20775 11543
rect 20717 11503 20775 11509
rect 22278 11500 22284 11552
rect 22336 11540 22342 11552
rect 22830 11540 22836 11552
rect 22336 11512 22836 11540
rect 22336 11500 22342 11512
rect 22830 11500 22836 11512
rect 22888 11500 22894 11552
rect 23477 11543 23535 11549
rect 23477 11509 23489 11543
rect 23523 11540 23535 11543
rect 24210 11540 24216 11552
rect 23523 11512 24216 11540
rect 23523 11509 23535 11512
rect 23477 11503 23535 11509
rect 24210 11500 24216 11512
rect 24268 11500 24274 11552
rect 24302 11500 24308 11552
rect 24360 11540 24366 11552
rect 24397 11543 24455 11549
rect 24397 11540 24409 11543
rect 24360 11512 24409 11540
rect 24360 11500 24366 11512
rect 24397 11509 24409 11512
rect 24443 11540 24455 11543
rect 26326 11540 26332 11552
rect 24443 11512 26332 11540
rect 24443 11509 24455 11512
rect 24397 11503 24455 11509
rect 26326 11500 26332 11512
rect 26384 11500 26390 11552
rect 1104 11450 28060 11472
rect 1104 11398 5442 11450
rect 5494 11398 5506 11450
rect 5558 11398 5570 11450
rect 5622 11398 5634 11450
rect 5686 11398 5698 11450
rect 5750 11398 14428 11450
rect 14480 11398 14492 11450
rect 14544 11398 14556 11450
rect 14608 11398 14620 11450
rect 14672 11398 14684 11450
rect 14736 11398 23413 11450
rect 23465 11398 23477 11450
rect 23529 11398 23541 11450
rect 23593 11398 23605 11450
rect 23657 11398 23669 11450
rect 23721 11398 28060 11450
rect 1104 11376 28060 11398
rect 6089 11339 6147 11345
rect 6089 11305 6101 11339
rect 6135 11336 6147 11339
rect 6454 11336 6460 11348
rect 6135 11308 6460 11336
rect 6135 11305 6147 11308
rect 6089 11299 6147 11305
rect 6454 11296 6460 11308
rect 6512 11296 6518 11348
rect 9306 11336 9312 11348
rect 9267 11308 9312 11336
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 9398 11296 9404 11348
rect 9456 11336 9462 11348
rect 9953 11339 10011 11345
rect 9953 11336 9965 11339
rect 9456 11308 9965 11336
rect 9456 11296 9462 11308
rect 9953 11305 9965 11308
rect 9999 11305 10011 11339
rect 10686 11336 10692 11348
rect 9953 11299 10011 11305
rect 10060 11308 10692 11336
rect 2682 11228 2688 11280
rect 2740 11268 2746 11280
rect 3878 11268 3884 11280
rect 2740 11240 3884 11268
rect 2740 11228 2746 11240
rect 3878 11228 3884 11240
rect 3936 11228 3942 11280
rect 6270 11228 6276 11280
rect 6328 11268 6334 11280
rect 7423 11271 7481 11277
rect 7423 11268 7435 11271
rect 6328 11240 7435 11268
rect 6328 11228 6334 11240
rect 7423 11237 7435 11240
rect 7469 11237 7481 11271
rect 7423 11231 7481 11237
rect 9858 11228 9864 11280
rect 9916 11268 9922 11280
rect 10060 11268 10088 11308
rect 10686 11296 10692 11308
rect 10744 11296 10750 11348
rect 11422 11296 11428 11348
rect 11480 11336 11486 11348
rect 12158 11336 12164 11348
rect 11480 11308 12164 11336
rect 11480 11296 11486 11308
rect 12158 11296 12164 11308
rect 12216 11336 12222 11348
rect 13722 11336 13728 11348
rect 12216 11308 13728 11336
rect 12216 11296 12222 11308
rect 13722 11296 13728 11308
rect 13780 11296 13786 11348
rect 13814 11296 13820 11348
rect 13872 11336 13878 11348
rect 14090 11336 14096 11348
rect 13872 11308 14096 11336
rect 13872 11296 13878 11308
rect 14090 11296 14096 11308
rect 14148 11296 14154 11348
rect 14461 11339 14519 11345
rect 14461 11305 14473 11339
rect 14507 11336 14519 11339
rect 15838 11336 15844 11348
rect 14507 11308 15844 11336
rect 14507 11305 14519 11308
rect 14461 11299 14519 11305
rect 15838 11296 15844 11308
rect 15896 11296 15902 11348
rect 17218 11336 17224 11348
rect 16592 11308 17224 11336
rect 16114 11268 16120 11280
rect 9916 11240 10088 11268
rect 10612 11240 16120 11268
rect 9916 11228 9922 11240
rect 6638 11200 6644 11212
rect 4908 11172 6644 11200
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11101 1731 11135
rect 1673 11095 1731 11101
rect 1940 11135 1998 11141
rect 1940 11101 1952 11135
rect 1986 11101 1998 11135
rect 1940 11095 1998 11101
rect 1688 10996 1716 11095
rect 1854 11024 1860 11076
rect 1912 11064 1918 11076
rect 1964 11064 1992 11095
rect 3326 11092 3332 11144
rect 3384 11132 3390 11144
rect 3510 11132 3516 11144
rect 3384 11104 3516 11132
rect 3384 11092 3390 11104
rect 3510 11092 3516 11104
rect 3568 11092 3574 11144
rect 3881 11135 3939 11141
rect 3881 11101 3893 11135
rect 3927 11132 3939 11135
rect 4908 11132 4936 11172
rect 6638 11160 6644 11172
rect 6696 11160 6702 11212
rect 6914 11160 6920 11212
rect 6972 11200 6978 11212
rect 10612 11200 10640 11240
rect 16114 11228 16120 11240
rect 16172 11228 16178 11280
rect 6972 11172 10640 11200
rect 6972 11160 6978 11172
rect 3927 11104 4936 11132
rect 5721 11135 5779 11141
rect 3927 11101 3939 11104
rect 3881 11095 3939 11101
rect 3896 11064 3924 11095
rect 4264 11076 4292 11104
rect 5721 11101 5733 11135
rect 5767 11101 5779 11135
rect 5902 11132 5908 11144
rect 5863 11104 5908 11132
rect 5721 11095 5779 11101
rect 1912 11036 1992 11064
rect 2047 11036 3924 11064
rect 4148 11067 4206 11073
rect 1912 11024 1918 11036
rect 2047 10996 2075 11036
rect 4148 11033 4160 11067
rect 4194 11033 4206 11067
rect 4148 11027 4206 11033
rect 1688 10968 2075 10996
rect 3053 10999 3111 11005
rect 3053 10965 3065 10999
rect 3099 10996 3111 10999
rect 3326 10996 3332 11008
rect 3099 10968 3332 10996
rect 3099 10965 3111 10968
rect 3053 10959 3111 10965
rect 3326 10956 3332 10968
rect 3384 10956 3390 11008
rect 4172 10996 4200 11027
rect 4246 11024 4252 11076
rect 4304 11024 4310 11076
rect 5736 11064 5764 11095
rect 5902 11092 5908 11104
rect 5960 11092 5966 11144
rect 6270 11092 6276 11144
rect 6328 11092 6334 11144
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11132 6791 11135
rect 7006 11132 7012 11144
rect 6779 11104 7012 11132
rect 6779 11101 6791 11104
rect 6733 11095 6791 11101
rect 7006 11092 7012 11104
rect 7064 11092 7070 11144
rect 7193 11135 7251 11141
rect 7193 11101 7205 11135
rect 7239 11132 7251 11135
rect 7650 11132 7656 11144
rect 7239 11104 7656 11132
rect 7239 11101 7251 11104
rect 7193 11095 7251 11101
rect 7650 11092 7656 11104
rect 7708 11132 7714 11144
rect 8846 11132 8852 11144
rect 7708 11104 8852 11132
rect 7708 11092 7714 11104
rect 8846 11092 8852 11104
rect 8904 11092 8910 11144
rect 8938 11092 8944 11144
rect 8996 11132 9002 11144
rect 9033 11135 9091 11141
rect 9033 11132 9045 11135
rect 8996 11104 9045 11132
rect 8996 11092 9002 11104
rect 9033 11101 9045 11104
rect 9079 11101 9091 11135
rect 9033 11095 9091 11101
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11132 9183 11135
rect 10502 11132 10508 11144
rect 9171 11104 10508 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 6288 11064 6316 11092
rect 6454 11064 6460 11076
rect 5092 11036 6460 11064
rect 4338 10996 4344 11008
rect 4172 10968 4344 10996
rect 4338 10956 4344 10968
rect 4396 10956 4402 11008
rect 4982 10956 4988 11008
rect 5040 10996 5046 11008
rect 5092 10996 5120 11036
rect 6454 11024 6460 11036
rect 6512 11024 6518 11076
rect 5258 10996 5264 11008
rect 5040 10968 5120 10996
rect 5219 10968 5264 10996
rect 5040 10956 5046 10968
rect 5258 10956 5264 10968
rect 5316 10956 5322 11008
rect 6549 10999 6607 11005
rect 6549 10965 6561 10999
rect 6595 10996 6607 10999
rect 6822 10996 6828 11008
rect 6595 10968 6828 10996
rect 6595 10965 6607 10968
rect 6549 10959 6607 10965
rect 6822 10956 6828 10968
rect 6880 10956 6886 11008
rect 7650 10956 7656 11008
rect 7708 10996 7714 11008
rect 8110 10996 8116 11008
rect 7708 10968 8116 10996
rect 7708 10956 7714 10968
rect 8110 10956 8116 10968
rect 8168 10956 8174 11008
rect 8386 10956 8392 11008
rect 8444 10996 8450 11008
rect 9048 10996 9076 11095
rect 10502 11092 10508 11104
rect 10560 11092 10566 11144
rect 10612 11141 10640 11172
rect 10962 11160 10968 11212
rect 11020 11200 11026 11212
rect 11020 11172 11652 11200
rect 11020 11160 11026 11172
rect 10597 11135 10655 11141
rect 10597 11101 10609 11135
rect 10643 11101 10655 11135
rect 11422 11132 11428 11144
rect 11383 11104 11428 11132
rect 10597 11095 10655 11101
rect 11422 11092 11428 11104
rect 11480 11092 11486 11144
rect 11624 11141 11652 11172
rect 13538 11160 13544 11212
rect 13596 11200 13602 11212
rect 15381 11203 15439 11209
rect 15381 11200 15393 11203
rect 13596 11172 15393 11200
rect 13596 11160 13602 11172
rect 15381 11169 15393 11172
rect 15427 11169 15439 11203
rect 15381 11163 15439 11169
rect 11609 11135 11667 11141
rect 11609 11101 11621 11135
rect 11655 11101 11667 11135
rect 11882 11132 11888 11144
rect 11843 11104 11888 11132
rect 11609 11095 11667 11101
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 12710 11132 12716 11144
rect 12671 11104 12716 11132
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 12989 11135 13047 11141
rect 12989 11101 13001 11135
rect 13035 11132 13047 11135
rect 13446 11132 13452 11144
rect 13035 11104 13452 11132
rect 13035 11101 13047 11104
rect 12989 11095 13047 11101
rect 13446 11092 13452 11104
rect 13504 11092 13510 11144
rect 13906 11092 13912 11144
rect 13964 11132 13970 11144
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13964 11104 14105 11132
rect 13964 11092 13970 11104
rect 14093 11101 14105 11104
rect 14139 11101 14151 11135
rect 14093 11095 14151 11101
rect 14274 11092 14280 11144
rect 14332 11132 14338 11144
rect 14369 11135 14427 11141
rect 14369 11132 14381 11135
rect 14332 11104 14381 11132
rect 14332 11092 14338 11104
rect 14369 11101 14381 11104
rect 14415 11101 14427 11135
rect 16482 11132 16488 11144
rect 16443 11104 16488 11132
rect 14369 11095 14427 11101
rect 16482 11092 16488 11104
rect 16540 11092 16546 11144
rect 16592 11141 16620 11308
rect 17218 11296 17224 11308
rect 17276 11296 17282 11348
rect 18693 11339 18751 11345
rect 18693 11305 18705 11339
rect 18739 11336 18751 11339
rect 18782 11336 18788 11348
rect 18739 11308 18788 11336
rect 18739 11305 18751 11308
rect 18693 11299 18751 11305
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 19797 11339 19855 11345
rect 19797 11305 19809 11339
rect 19843 11336 19855 11339
rect 20438 11336 20444 11348
rect 19843 11308 20444 11336
rect 19843 11305 19855 11308
rect 19797 11299 19855 11305
rect 20438 11296 20444 11308
rect 20496 11296 20502 11348
rect 21634 11336 21640 11348
rect 21595 11308 21640 11336
rect 21634 11296 21640 11308
rect 21692 11296 21698 11348
rect 23198 11296 23204 11348
rect 23256 11336 23262 11348
rect 26329 11339 26387 11345
rect 23256 11308 25728 11336
rect 23256 11296 23262 11308
rect 16666 11228 16672 11280
rect 16724 11268 16730 11280
rect 16724 11240 17356 11268
rect 16724 11228 16730 11240
rect 17328 11209 17356 11240
rect 24210 11228 24216 11280
rect 24268 11268 24274 11280
rect 24268 11240 25636 11268
rect 24268 11228 24274 11240
rect 16761 11203 16819 11209
rect 16761 11169 16773 11203
rect 16807 11169 16819 11203
rect 16761 11163 16819 11169
rect 17313 11203 17371 11209
rect 17313 11169 17325 11203
rect 17359 11169 17371 11203
rect 17313 11163 17371 11169
rect 16577 11135 16635 11141
rect 16577 11101 16589 11135
rect 16623 11101 16635 11135
rect 16577 11095 16635 11101
rect 9674 11024 9680 11076
rect 9732 11064 9738 11076
rect 9861 11067 9919 11073
rect 9861 11064 9873 11067
rect 9732 11036 9873 11064
rect 9732 11024 9738 11036
rect 9861 11033 9873 11036
rect 9907 11064 9919 11067
rect 10686 11064 10692 11076
rect 9907 11036 10692 11064
rect 9907 11033 9919 11036
rect 9861 11027 9919 11033
rect 10686 11024 10692 11036
rect 10744 11024 10750 11076
rect 10781 11067 10839 11073
rect 10781 11033 10793 11067
rect 10827 11064 10839 11067
rect 12618 11064 12624 11076
rect 10827 11036 12624 11064
rect 10827 11033 10839 11036
rect 10781 11027 10839 11033
rect 12618 11024 12624 11036
rect 12676 11064 12682 11076
rect 15197 11067 15255 11073
rect 15197 11064 15209 11067
rect 12676 11036 15209 11064
rect 12676 11024 12682 11036
rect 15197 11033 15209 11036
rect 15243 11033 15255 11067
rect 15197 11027 15255 11033
rect 16301 11067 16359 11073
rect 16301 11033 16313 11067
rect 16347 11033 16359 11067
rect 16301 11027 16359 11033
rect 10962 10996 10968 11008
rect 8444 10968 10968 10996
rect 8444 10956 8450 10968
rect 10962 10956 10968 10968
rect 11020 10956 11026 11008
rect 12250 10956 12256 11008
rect 12308 10996 12314 11008
rect 14182 10996 14188 11008
rect 12308 10968 14188 10996
rect 12308 10956 12314 10968
rect 14182 10956 14188 10968
rect 14240 10956 14246 11008
rect 14274 10956 14280 11008
rect 14332 10996 14338 11008
rect 14645 10999 14703 11005
rect 14645 10996 14657 10999
rect 14332 10968 14657 10996
rect 14332 10956 14338 10968
rect 14645 10965 14657 10968
rect 14691 10965 14703 10999
rect 16316 10996 16344 11027
rect 16390 11024 16396 11076
rect 16448 11064 16454 11076
rect 16776 11064 16804 11163
rect 16853 11135 16911 11141
rect 16853 11101 16865 11135
rect 16899 11101 16911 11135
rect 17328 11132 17356 11163
rect 21910 11160 21916 11212
rect 21968 11200 21974 11212
rect 22097 11203 22155 11209
rect 22097 11200 22109 11203
rect 21968 11172 22109 11200
rect 21968 11160 21974 11172
rect 22097 11169 22109 11172
rect 22143 11169 22155 11203
rect 22097 11163 22155 11169
rect 24302 11160 24308 11212
rect 24360 11200 24366 11212
rect 24489 11203 24547 11209
rect 24489 11200 24501 11203
rect 24360 11172 24501 11200
rect 24360 11160 24366 11172
rect 24489 11169 24501 11172
rect 24535 11200 24547 11203
rect 25498 11200 25504 11212
rect 24535 11172 25504 11200
rect 24535 11169 24547 11172
rect 24489 11163 24547 11169
rect 25498 11160 25504 11172
rect 25556 11160 25562 11212
rect 19702 11132 19708 11144
rect 17328 11104 19708 11132
rect 16853 11095 16911 11101
rect 16448 11036 16804 11064
rect 16868 11064 16896 11095
rect 19702 11092 19708 11104
rect 19760 11132 19766 11144
rect 20257 11135 20315 11141
rect 20257 11132 20269 11135
rect 19760 11104 20269 11132
rect 19760 11092 19766 11104
rect 20257 11101 20269 11104
rect 20303 11101 20315 11135
rect 20257 11095 20315 11101
rect 20346 11092 20352 11144
rect 20404 11132 20410 11144
rect 20513 11135 20571 11141
rect 20513 11132 20525 11135
rect 20404 11104 20525 11132
rect 20404 11092 20410 11104
rect 20513 11101 20525 11104
rect 20559 11101 20571 11135
rect 22738 11132 22744 11144
rect 20513 11095 20571 11101
rect 22296 11104 22744 11132
rect 17580 11067 17638 11073
rect 16868 11036 17540 11064
rect 16448 11024 16454 11036
rect 16482 10996 16488 11008
rect 16316 10968 16488 10996
rect 14645 10959 14703 10965
rect 16482 10956 16488 10968
rect 16540 10956 16546 11008
rect 17512 10996 17540 11036
rect 17580 11033 17592 11067
rect 17626 11064 17638 11067
rect 19150 11064 19156 11076
rect 17626 11036 19156 11064
rect 17626 11033 17638 11036
rect 17580 11027 17638 11033
rect 19150 11024 19156 11036
rect 19208 11024 19214 11076
rect 19426 11064 19432 11076
rect 19387 11036 19432 11064
rect 19426 11024 19432 11036
rect 19484 11024 19490 11076
rect 19518 11024 19524 11076
rect 19576 11064 19582 11076
rect 19613 11067 19671 11073
rect 19613 11064 19625 11067
rect 19576 11036 19625 11064
rect 19576 11024 19582 11036
rect 19613 11033 19625 11036
rect 19659 11033 19671 11067
rect 19613 11027 19671 11033
rect 19794 11024 19800 11076
rect 19852 11064 19858 11076
rect 22296 11064 22324 11104
rect 22738 11092 22744 11104
rect 22796 11092 22802 11144
rect 24394 11132 24400 11144
rect 24355 11104 24400 11132
rect 24394 11092 24400 11104
rect 24452 11092 24458 11144
rect 25608 11141 25636 11240
rect 24949 11135 25007 11141
rect 24949 11101 24961 11135
rect 24995 11101 25007 11135
rect 24949 11095 25007 11101
rect 25409 11135 25467 11141
rect 25409 11101 25421 11135
rect 25455 11101 25467 11135
rect 25409 11095 25467 11101
rect 25593 11135 25651 11141
rect 25593 11101 25605 11135
rect 25639 11101 25651 11135
rect 25700 11132 25728 11308
rect 26329 11305 26341 11339
rect 26375 11336 26387 11339
rect 26418 11336 26424 11348
rect 26375 11308 26424 11336
rect 26375 11305 26387 11308
rect 26329 11299 26387 11305
rect 26418 11296 26424 11308
rect 26476 11296 26482 11348
rect 27246 11296 27252 11348
rect 27304 11336 27310 11348
rect 27614 11336 27620 11348
rect 27304 11308 27620 11336
rect 27304 11296 27310 11308
rect 27614 11296 27620 11308
rect 27672 11296 27678 11348
rect 26326 11160 26332 11212
rect 26384 11200 26390 11212
rect 26697 11203 26755 11209
rect 26697 11200 26709 11203
rect 26384 11172 26709 11200
rect 26384 11160 26390 11172
rect 26697 11169 26709 11172
rect 26743 11169 26755 11203
rect 26697 11163 26755 11169
rect 26789 11203 26847 11209
rect 26789 11169 26801 11203
rect 26835 11200 26847 11203
rect 26878 11200 26884 11212
rect 26835 11172 26884 11200
rect 26835 11169 26847 11172
rect 26789 11163 26847 11169
rect 26878 11160 26884 11172
rect 26936 11160 26942 11212
rect 26513 11135 26571 11141
rect 26513 11132 26525 11135
rect 25700 11104 26525 11132
rect 25593 11095 25651 11101
rect 26513 11101 26525 11104
rect 26559 11101 26571 11135
rect 26513 11095 26571 11101
rect 19852 11036 22324 11064
rect 22364 11067 22422 11073
rect 19852 11024 19858 11036
rect 22364 11033 22376 11067
rect 22410 11064 22422 11067
rect 22462 11064 22468 11076
rect 22410 11036 22468 11064
rect 22410 11033 22422 11036
rect 22364 11027 22422 11033
rect 22462 11024 22468 11036
rect 22520 11024 22526 11076
rect 23290 11024 23296 11076
rect 23348 11064 23354 11076
rect 24964 11064 24992 11095
rect 23348 11036 24992 11064
rect 23348 11024 23354 11036
rect 25038 11024 25044 11076
rect 25096 11064 25102 11076
rect 25424 11064 25452 11095
rect 26326 11064 26332 11076
rect 25096 11036 25360 11064
rect 25424 11036 26332 11064
rect 25096 11024 25102 11036
rect 18046 10996 18052 11008
rect 17512 10968 18052 10996
rect 18046 10956 18052 10968
rect 18104 10956 18110 11008
rect 18230 10956 18236 11008
rect 18288 10996 18294 11008
rect 20898 10996 20904 11008
rect 18288 10968 20904 10996
rect 18288 10956 18294 10968
rect 20898 10956 20904 10968
rect 20956 10956 20962 11008
rect 20990 10956 20996 11008
rect 21048 10996 21054 11008
rect 21266 10996 21272 11008
rect 21048 10968 21272 10996
rect 21048 10956 21054 10968
rect 21266 10956 21272 10968
rect 21324 10956 21330 11008
rect 23477 10999 23535 11005
rect 23477 10965 23489 10999
rect 23523 10996 23535 10999
rect 23842 10996 23848 11008
rect 23523 10968 23848 10996
rect 23523 10965 23535 10968
rect 23477 10959 23535 10965
rect 23842 10956 23848 10968
rect 23900 10956 23906 11008
rect 24118 10956 24124 11008
rect 24176 10996 24182 11008
rect 24486 10996 24492 11008
rect 24176 10968 24492 10996
rect 24176 10956 24182 10968
rect 24486 10956 24492 10968
rect 24544 10956 24550 11008
rect 25332 10996 25360 11036
rect 26326 11024 26332 11036
rect 26384 11024 26390 11076
rect 25590 10996 25596 11008
rect 25332 10968 25596 10996
rect 25590 10956 25596 10968
rect 25648 10956 25654 11008
rect 1104 10906 28060 10928
rect 1104 10854 9935 10906
rect 9987 10854 9999 10906
rect 10051 10854 10063 10906
rect 10115 10854 10127 10906
rect 10179 10854 10191 10906
rect 10243 10854 18920 10906
rect 18972 10854 18984 10906
rect 19036 10854 19048 10906
rect 19100 10854 19112 10906
rect 19164 10854 19176 10906
rect 19228 10854 28060 10906
rect 1104 10832 28060 10854
rect 2038 10752 2044 10804
rect 2096 10792 2102 10804
rect 2225 10795 2283 10801
rect 2225 10792 2237 10795
rect 2096 10764 2237 10792
rect 2096 10752 2102 10764
rect 2225 10761 2237 10764
rect 2271 10761 2283 10795
rect 2225 10755 2283 10761
rect 3878 10752 3884 10804
rect 3936 10792 3942 10804
rect 3936 10764 5672 10792
rect 3936 10752 3942 10764
rect 1857 10727 1915 10733
rect 1857 10693 1869 10727
rect 1903 10724 1915 10727
rect 3053 10727 3111 10733
rect 3053 10724 3065 10727
rect 1903 10696 3065 10724
rect 1903 10693 1915 10696
rect 1857 10687 1915 10693
rect 3053 10693 3065 10696
rect 3099 10693 3111 10727
rect 3418 10724 3424 10736
rect 3053 10687 3111 10693
rect 3252 10696 3424 10724
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10656 2099 10659
rect 2130 10656 2136 10668
rect 2087 10628 2136 10656
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 2130 10616 2136 10628
rect 2188 10616 2194 10668
rect 3252 10665 3280 10696
rect 3418 10684 3424 10696
rect 3476 10684 3482 10736
rect 4982 10724 4988 10736
rect 4540 10696 4988 10724
rect 3237 10659 3295 10665
rect 3237 10625 3249 10659
rect 3283 10625 3295 10659
rect 3237 10619 3295 10625
rect 3326 10616 3332 10668
rect 3384 10656 3390 10668
rect 4540 10665 4568 10696
rect 4982 10684 4988 10696
rect 5040 10684 5046 10736
rect 5534 10724 5540 10736
rect 5495 10696 5540 10724
rect 5534 10684 5540 10696
rect 5592 10684 5598 10736
rect 5644 10724 5672 10764
rect 5718 10752 5724 10804
rect 5776 10792 5782 10804
rect 6546 10792 6552 10804
rect 5776 10764 6552 10792
rect 5776 10752 5782 10764
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 7006 10752 7012 10804
rect 7064 10792 7070 10804
rect 8757 10795 8815 10801
rect 8757 10792 8769 10795
rect 7064 10764 8769 10792
rect 7064 10752 7070 10764
rect 8757 10761 8769 10764
rect 8803 10761 8815 10795
rect 8757 10755 8815 10761
rect 9214 10752 9220 10804
rect 9272 10792 9278 10804
rect 10781 10795 10839 10801
rect 9272 10764 10640 10792
rect 9272 10752 9278 10764
rect 10134 10724 10140 10736
rect 5644 10696 10140 10724
rect 10134 10684 10140 10696
rect 10192 10684 10198 10736
rect 10612 10733 10640 10764
rect 10781 10761 10793 10795
rect 10827 10792 10839 10795
rect 11790 10792 11796 10804
rect 10827 10764 11796 10792
rect 10827 10761 10839 10764
rect 10781 10755 10839 10761
rect 11790 10752 11796 10764
rect 11848 10752 11854 10804
rect 12069 10795 12127 10801
rect 12069 10761 12081 10795
rect 12115 10792 12127 10795
rect 12342 10792 12348 10804
rect 12115 10764 12348 10792
rect 12115 10761 12127 10764
rect 12069 10755 12127 10761
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 13906 10752 13912 10804
rect 13964 10792 13970 10804
rect 14829 10795 14887 10801
rect 14829 10792 14841 10795
rect 13964 10764 14841 10792
rect 13964 10752 13970 10764
rect 14829 10761 14841 10764
rect 14875 10761 14887 10795
rect 14829 10755 14887 10761
rect 15838 10752 15844 10804
rect 15896 10792 15902 10804
rect 16390 10792 16396 10804
rect 15896 10764 16396 10792
rect 15896 10752 15902 10764
rect 16390 10752 16396 10764
rect 16448 10752 16454 10804
rect 17310 10752 17316 10804
rect 17368 10792 17374 10804
rect 17368 10764 20300 10792
rect 17368 10752 17374 10764
rect 10597 10727 10655 10733
rect 10597 10693 10609 10727
rect 10643 10693 10655 10727
rect 10597 10687 10655 10693
rect 14366 10684 14372 10736
rect 14424 10724 14430 10736
rect 16936 10727 16994 10733
rect 14424 10696 15976 10724
rect 14424 10684 14430 10696
rect 3605 10659 3663 10665
rect 3384 10628 3429 10656
rect 3384 10616 3390 10628
rect 3605 10625 3617 10659
rect 3651 10625 3663 10659
rect 3605 10619 3663 10625
rect 4525 10659 4583 10665
rect 4525 10625 4537 10659
rect 4571 10625 4583 10659
rect 4525 10619 4583 10625
rect 4617 10659 4675 10665
rect 4617 10625 4629 10659
rect 4663 10625 4675 10659
rect 5258 10656 5264 10668
rect 5219 10628 5264 10656
rect 4617 10619 4675 10625
rect 2222 10548 2228 10600
rect 2280 10588 2286 10600
rect 3620 10588 3648 10619
rect 2280 10560 3648 10588
rect 4632 10588 4660 10619
rect 5258 10616 5264 10628
rect 5316 10616 5322 10668
rect 5350 10616 5356 10668
rect 5408 10656 5414 10668
rect 5445 10659 5503 10665
rect 5445 10656 5457 10659
rect 5408 10628 5457 10656
rect 5408 10616 5414 10628
rect 5445 10625 5457 10628
rect 5491 10625 5503 10659
rect 5445 10619 5503 10625
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10656 5687 10659
rect 6549 10659 6607 10665
rect 5675 10628 5948 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 5920 10588 5948 10628
rect 6549 10625 6561 10659
rect 6595 10656 6607 10659
rect 6638 10656 6644 10668
rect 6595 10628 6644 10656
rect 6595 10625 6607 10628
rect 6549 10619 6607 10625
rect 6638 10616 6644 10628
rect 6696 10616 6702 10668
rect 6822 10665 6828 10668
rect 6816 10656 6828 10665
rect 6783 10628 6828 10656
rect 6816 10619 6828 10628
rect 6822 10616 6828 10619
rect 6880 10616 6886 10668
rect 7374 10616 7380 10668
rect 7432 10656 7438 10668
rect 7558 10656 7564 10668
rect 7432 10628 7564 10656
rect 7432 10616 7438 10628
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 7650 10616 7656 10668
rect 7708 10616 7714 10668
rect 8110 10616 8116 10668
rect 8168 10656 8174 10668
rect 8573 10659 8631 10665
rect 8573 10656 8585 10659
rect 8168 10628 8585 10656
rect 8168 10616 8174 10628
rect 8573 10625 8585 10628
rect 8619 10625 8631 10659
rect 8573 10619 8631 10625
rect 9861 10659 9919 10665
rect 9861 10625 9873 10659
rect 9907 10656 9919 10659
rect 9950 10656 9956 10668
rect 9907 10628 9956 10656
rect 9907 10625 9919 10628
rect 9861 10619 9919 10625
rect 9950 10616 9956 10628
rect 10008 10616 10014 10668
rect 10045 10659 10103 10665
rect 10045 10625 10057 10659
rect 10091 10656 10103 10659
rect 10091 10628 10640 10656
rect 10091 10625 10103 10628
rect 10045 10619 10103 10625
rect 5994 10588 6000 10600
rect 4632 10560 5856 10588
rect 5920 10560 6000 10588
rect 2280 10548 2286 10560
rect 4982 10520 4988 10532
rect 2746 10492 4988 10520
rect 1394 10412 1400 10464
rect 1452 10452 1458 10464
rect 2746 10452 2774 10492
rect 4982 10480 4988 10492
rect 5040 10480 5046 10532
rect 5828 10529 5856 10560
rect 5994 10548 6000 10560
rect 6052 10588 6058 10600
rect 6052 10560 6592 10588
rect 6052 10548 6058 10560
rect 6564 10532 6592 10560
rect 5813 10523 5871 10529
rect 5813 10489 5825 10523
rect 5859 10489 5871 10523
rect 5813 10483 5871 10489
rect 6546 10480 6552 10532
rect 6604 10480 6610 10532
rect 7668 10520 7696 10616
rect 8386 10588 8392 10600
rect 8347 10560 8392 10588
rect 8386 10548 8392 10560
rect 8444 10548 8450 10600
rect 10137 10591 10195 10597
rect 10137 10557 10149 10591
rect 10183 10588 10195 10591
rect 10318 10588 10324 10600
rect 10183 10560 10324 10588
rect 10183 10557 10195 10560
rect 10137 10551 10195 10557
rect 10318 10548 10324 10560
rect 10376 10548 10382 10600
rect 7484 10492 7696 10520
rect 7484 10464 7512 10492
rect 1452 10424 2774 10452
rect 3513 10455 3571 10461
rect 1452 10412 1458 10424
rect 3513 10421 3525 10455
rect 3559 10452 3571 10455
rect 3970 10452 3976 10464
rect 3559 10424 3976 10452
rect 3559 10421 3571 10424
rect 3513 10415 3571 10421
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 4798 10452 4804 10464
rect 4759 10424 4804 10452
rect 4798 10412 4804 10424
rect 4856 10412 4862 10464
rect 7466 10412 7472 10464
rect 7524 10412 7530 10464
rect 7558 10412 7564 10464
rect 7616 10452 7622 10464
rect 10612 10461 10640 10628
rect 10686 10616 10692 10668
rect 10744 10656 10750 10668
rect 10873 10659 10931 10665
rect 10873 10656 10885 10659
rect 10744 10628 10885 10656
rect 10744 10616 10750 10628
rect 10873 10625 10885 10628
rect 10919 10625 10931 10659
rect 10873 10619 10931 10625
rect 11146 10616 11152 10668
rect 11204 10656 11210 10668
rect 11885 10659 11943 10665
rect 11885 10656 11897 10659
rect 11204 10628 11897 10656
rect 11204 10616 11210 10628
rect 11885 10625 11897 10628
rect 11931 10656 11943 10659
rect 11974 10656 11980 10668
rect 11931 10628 11980 10656
rect 11931 10625 11943 10628
rect 11885 10619 11943 10625
rect 11974 10616 11980 10628
rect 12032 10616 12038 10668
rect 12161 10659 12219 10665
rect 12161 10625 12173 10659
rect 12207 10656 12219 10659
rect 12342 10656 12348 10668
rect 12207 10628 12348 10656
rect 12207 10625 12219 10628
rect 12161 10619 12219 10625
rect 12342 10616 12348 10628
rect 12400 10616 12406 10668
rect 12526 10616 12532 10668
rect 12584 10656 12590 10668
rect 12621 10659 12679 10665
rect 12621 10656 12633 10659
rect 12584 10628 12633 10656
rect 12584 10616 12590 10628
rect 12621 10625 12633 10628
rect 12667 10625 12679 10659
rect 13538 10656 13544 10668
rect 12621 10619 12679 10625
rect 13464 10628 13544 10656
rect 11698 10548 11704 10600
rect 11756 10588 11762 10600
rect 13464 10597 13492 10628
rect 13538 10616 13544 10628
rect 13596 10616 13602 10668
rect 13716 10659 13774 10665
rect 13716 10625 13728 10659
rect 13762 10656 13774 10659
rect 14090 10656 14096 10668
rect 13762 10628 14096 10656
rect 13762 10625 13774 10628
rect 13716 10619 13774 10625
rect 14090 10616 14096 10628
rect 14148 10616 14154 10668
rect 15654 10656 15660 10668
rect 15615 10628 15660 10656
rect 15654 10616 15660 10628
rect 15712 10616 15718 10668
rect 15838 10656 15844 10668
rect 15799 10628 15844 10656
rect 15838 10616 15844 10628
rect 15896 10616 15902 10668
rect 15948 10665 15976 10696
rect 16936 10693 16948 10727
rect 16982 10724 16994 10727
rect 19972 10727 20030 10733
rect 16982 10696 19932 10724
rect 16982 10693 16994 10696
rect 16936 10687 16994 10693
rect 15933 10659 15991 10665
rect 15933 10625 15945 10659
rect 15979 10656 15991 10659
rect 16390 10656 16396 10668
rect 15979 10628 16396 10656
rect 15979 10625 15991 10628
rect 15933 10619 15991 10625
rect 16390 10616 16396 10628
rect 16448 10616 16454 10668
rect 16666 10656 16672 10668
rect 16579 10628 16672 10656
rect 13449 10591 13507 10597
rect 13449 10588 13461 10591
rect 11756 10560 13461 10588
rect 11756 10548 11762 10560
rect 13449 10557 13461 10560
rect 13495 10557 13507 10591
rect 13449 10551 13507 10557
rect 15010 10548 15016 10600
rect 15068 10588 15074 10600
rect 16592 10588 16620 10628
rect 16666 10616 16672 10628
rect 16724 10616 16730 10668
rect 19061 10659 19119 10665
rect 16776 10628 19012 10656
rect 16776 10588 16804 10628
rect 15068 10560 16620 10588
rect 16684 10560 16804 10588
rect 15068 10548 15074 10560
rect 12805 10523 12863 10529
rect 12805 10489 12817 10523
rect 12851 10520 12863 10523
rect 13078 10520 13084 10532
rect 12851 10492 13084 10520
rect 12851 10489 12863 10492
rect 12805 10483 12863 10489
rect 13078 10480 13084 10492
rect 13136 10480 13142 10532
rect 15654 10480 15660 10532
rect 15712 10520 15718 10532
rect 16684 10520 16712 10560
rect 17862 10548 17868 10600
rect 17920 10588 17926 10600
rect 18877 10591 18935 10597
rect 18877 10588 18889 10591
rect 17920 10560 18889 10588
rect 17920 10548 17926 10560
rect 18877 10557 18889 10560
rect 18923 10557 18935 10591
rect 18877 10551 18935 10557
rect 18046 10520 18052 10532
rect 15712 10492 16712 10520
rect 18007 10492 18052 10520
rect 15712 10480 15718 10492
rect 18046 10480 18052 10492
rect 18104 10480 18110 10532
rect 7929 10455 7987 10461
rect 7929 10452 7941 10455
rect 7616 10424 7941 10452
rect 7616 10412 7622 10424
rect 7929 10421 7941 10424
rect 7975 10421 7987 10455
rect 7929 10415 7987 10421
rect 10597 10455 10655 10461
rect 10597 10421 10609 10455
rect 10643 10452 10655 10455
rect 11054 10452 11060 10464
rect 10643 10424 11060 10452
rect 10643 10421 10655 10424
rect 10597 10415 10655 10421
rect 11054 10412 11060 10424
rect 11112 10412 11118 10464
rect 11882 10452 11888 10464
rect 11843 10424 11888 10452
rect 11882 10412 11888 10424
rect 11940 10412 11946 10464
rect 15286 10412 15292 10464
rect 15344 10452 15350 10464
rect 15473 10455 15531 10461
rect 15473 10452 15485 10455
rect 15344 10424 15485 10452
rect 15344 10412 15350 10424
rect 15473 10421 15485 10424
rect 15519 10421 15531 10455
rect 18984 10452 19012 10628
rect 19061 10625 19073 10659
rect 19107 10656 19119 10659
rect 19518 10656 19524 10668
rect 19107 10628 19524 10656
rect 19107 10625 19119 10628
rect 19061 10619 19119 10625
rect 19518 10616 19524 10628
rect 19576 10616 19582 10668
rect 19702 10656 19708 10668
rect 19663 10628 19708 10656
rect 19702 10616 19708 10628
rect 19760 10616 19766 10668
rect 19904 10656 19932 10696
rect 19972 10693 19984 10727
rect 20018 10724 20030 10727
rect 20162 10724 20168 10736
rect 20018 10696 20168 10724
rect 20018 10693 20030 10696
rect 19972 10687 20030 10693
rect 20162 10684 20168 10696
rect 20220 10684 20226 10736
rect 20272 10724 20300 10764
rect 20714 10752 20720 10804
rect 20772 10792 20778 10804
rect 21085 10795 21143 10801
rect 21085 10792 21097 10795
rect 20772 10764 21097 10792
rect 20772 10752 20778 10764
rect 21085 10761 21097 10764
rect 21131 10761 21143 10795
rect 21085 10755 21143 10761
rect 21450 10752 21456 10804
rect 21508 10792 21514 10804
rect 21508 10764 22327 10792
rect 21508 10752 21514 10764
rect 20898 10724 20904 10736
rect 20272 10696 20904 10724
rect 20898 10684 20904 10696
rect 20956 10684 20962 10736
rect 22299 10724 22327 10764
rect 22370 10752 22376 10804
rect 22428 10792 22434 10804
rect 26326 10792 26332 10804
rect 22428 10764 25360 10792
rect 26287 10764 26332 10792
rect 22428 10752 22434 10764
rect 22299 10696 23152 10724
rect 21358 10656 21364 10668
rect 19904 10628 21364 10656
rect 21358 10616 21364 10628
rect 21416 10616 21422 10668
rect 21910 10616 21916 10668
rect 21968 10656 21974 10668
rect 22189 10659 22247 10665
rect 22189 10656 22201 10659
rect 21968 10628 22201 10656
rect 21968 10616 21974 10628
rect 22189 10625 22201 10628
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 22922 10616 22928 10668
rect 22980 10656 22986 10668
rect 23017 10659 23075 10665
rect 23017 10656 23029 10659
rect 22980 10628 23029 10656
rect 22980 10616 22986 10628
rect 23017 10625 23029 10628
rect 23063 10625 23075 10659
rect 23017 10619 23075 10625
rect 19150 10548 19156 10600
rect 19208 10588 19214 10600
rect 23124 10597 23152 10696
rect 24854 10684 24860 10736
rect 24912 10724 24918 10736
rect 25194 10727 25252 10733
rect 25194 10724 25206 10727
rect 24912 10696 25206 10724
rect 24912 10684 24918 10696
rect 25194 10693 25206 10696
rect 25240 10693 25252 10727
rect 25332 10724 25360 10764
rect 26326 10752 26332 10764
rect 26384 10752 26390 10804
rect 27798 10724 27804 10736
rect 25332 10696 27804 10724
rect 25194 10687 25252 10693
rect 27798 10684 27804 10696
rect 27856 10684 27862 10736
rect 23290 10616 23296 10668
rect 23348 10656 23354 10668
rect 23569 10659 23627 10665
rect 23569 10656 23581 10659
rect 23348 10628 23581 10656
rect 23348 10616 23354 10628
rect 23569 10625 23581 10628
rect 23615 10625 23627 10659
rect 23842 10656 23848 10668
rect 23803 10628 23848 10656
rect 23569 10619 23627 10625
rect 23842 10616 23848 10628
rect 23900 10616 23906 10668
rect 24210 10656 24216 10668
rect 24171 10628 24216 10656
rect 24210 10616 24216 10628
rect 24268 10616 24274 10668
rect 24762 10616 24768 10668
rect 24820 10656 24826 10668
rect 24949 10659 25007 10665
rect 24949 10656 24961 10659
rect 24820 10628 24961 10656
rect 24820 10616 24826 10628
rect 24949 10625 24961 10628
rect 24995 10625 25007 10659
rect 24949 10619 25007 10625
rect 25498 10616 25504 10668
rect 25556 10656 25562 10668
rect 27157 10659 27215 10665
rect 27157 10656 27169 10659
rect 25556 10628 27169 10656
rect 25556 10616 25562 10628
rect 27157 10625 27169 10628
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 19245 10591 19303 10597
rect 19245 10588 19257 10591
rect 19208 10560 19257 10588
rect 19208 10548 19214 10560
rect 19245 10557 19257 10560
rect 19291 10557 19303 10591
rect 19245 10551 19303 10557
rect 23109 10591 23167 10597
rect 23109 10557 23121 10591
rect 23155 10588 23167 10591
rect 23934 10588 23940 10600
rect 23155 10560 23940 10588
rect 23155 10557 23167 10560
rect 23109 10551 23167 10557
rect 23934 10548 23940 10560
rect 23992 10548 23998 10600
rect 20622 10452 20628 10464
rect 18984 10424 20628 10452
rect 15473 10415 15531 10421
rect 20622 10412 20628 10424
rect 20680 10412 20686 10464
rect 22005 10455 22063 10461
rect 22005 10421 22017 10455
rect 22051 10452 22063 10455
rect 22830 10452 22836 10464
rect 22051 10424 22836 10452
rect 22051 10421 22063 10424
rect 22005 10415 22063 10421
rect 22830 10412 22836 10424
rect 22888 10412 22894 10464
rect 26326 10412 26332 10464
rect 26384 10452 26390 10464
rect 26973 10455 27031 10461
rect 26973 10452 26985 10455
rect 26384 10424 26985 10452
rect 26384 10412 26390 10424
rect 26973 10421 26985 10424
rect 27019 10421 27031 10455
rect 26973 10415 27031 10421
rect 1104 10362 28060 10384
rect 1104 10310 5442 10362
rect 5494 10310 5506 10362
rect 5558 10310 5570 10362
rect 5622 10310 5634 10362
rect 5686 10310 5698 10362
rect 5750 10310 14428 10362
rect 14480 10310 14492 10362
rect 14544 10310 14556 10362
rect 14608 10310 14620 10362
rect 14672 10310 14684 10362
rect 14736 10310 23413 10362
rect 23465 10310 23477 10362
rect 23529 10310 23541 10362
rect 23593 10310 23605 10362
rect 23657 10310 23669 10362
rect 23721 10310 28060 10362
rect 1104 10288 28060 10310
rect 2590 10208 2596 10260
rect 2648 10248 2654 10260
rect 2866 10248 2872 10260
rect 2648 10220 2872 10248
rect 2648 10208 2654 10220
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 3326 10208 3332 10260
rect 3384 10248 3390 10260
rect 4617 10251 4675 10257
rect 4617 10248 4629 10251
rect 3384 10220 4629 10248
rect 3384 10208 3390 10220
rect 4617 10217 4629 10220
rect 4663 10217 4675 10251
rect 6914 10248 6920 10260
rect 4617 10211 4675 10217
rect 6012 10220 6920 10248
rect 3053 10183 3111 10189
rect 1780 10152 2774 10180
rect 1780 10053 1808 10152
rect 2746 10112 2774 10152
rect 3053 10149 3065 10183
rect 3099 10180 3111 10183
rect 4338 10180 4344 10192
rect 3099 10152 4344 10180
rect 3099 10149 3111 10152
rect 3053 10143 3111 10149
rect 4338 10140 4344 10152
rect 4396 10140 4402 10192
rect 6012 10180 6040 10220
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 8110 10248 8116 10260
rect 8071 10220 8116 10248
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 11517 10251 11575 10257
rect 11517 10248 11529 10251
rect 9508 10220 11529 10248
rect 4632 10152 6040 10180
rect 6089 10183 6147 10189
rect 4632 10112 4660 10152
rect 6089 10149 6101 10183
rect 6135 10149 6147 10183
rect 6089 10143 6147 10149
rect 2746 10084 4660 10112
rect 4709 10115 4767 10121
rect 4709 10081 4721 10115
rect 4755 10112 4767 10115
rect 6104 10112 6132 10143
rect 4755 10084 6040 10112
rect 6104 10084 6776 10112
rect 4755 10081 4767 10084
rect 4709 10075 4767 10081
rect 1765 10047 1823 10053
rect 1765 10013 1777 10047
rect 1811 10013 1823 10047
rect 1765 10007 1823 10013
rect 2409 10047 2467 10053
rect 2409 10013 2421 10047
rect 2455 10044 2467 10047
rect 2866 10044 2872 10056
rect 2455 10016 2872 10044
rect 2455 10013 2467 10016
rect 2409 10007 2467 10013
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10044 3295 10047
rect 4798 10044 4804 10056
rect 3283 10016 4804 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 4798 10004 4804 10016
rect 4856 10004 4862 10056
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10044 4951 10047
rect 5258 10044 5264 10056
rect 4939 10016 5264 10044
rect 4939 10013 4951 10016
rect 4893 10007 4951 10013
rect 5258 10004 5264 10016
rect 5316 10004 5322 10056
rect 5534 10044 5540 10056
rect 5495 10016 5540 10044
rect 5534 10004 5540 10016
rect 5592 10004 5598 10056
rect 5813 10047 5871 10053
rect 5813 10044 5825 10047
rect 5644 10016 5825 10044
rect 3973 9979 4031 9985
rect 3973 9945 3985 9979
rect 4019 9976 4031 9979
rect 4019 9948 4200 9976
rect 4019 9945 4031 9948
rect 3973 9939 4031 9945
rect 1578 9908 1584 9920
rect 1539 9880 1584 9908
rect 1578 9868 1584 9880
rect 1636 9868 1642 9920
rect 2222 9908 2228 9920
rect 2183 9880 2228 9908
rect 2222 9868 2228 9880
rect 2280 9868 2286 9920
rect 3418 9868 3424 9920
rect 3476 9908 3482 9920
rect 4065 9911 4123 9917
rect 4065 9908 4077 9911
rect 3476 9880 4077 9908
rect 3476 9868 3482 9880
rect 4065 9877 4077 9880
rect 4111 9877 4123 9911
rect 4172 9908 4200 9948
rect 4246 9936 4252 9988
rect 4304 9976 4310 9988
rect 4617 9979 4675 9985
rect 4617 9976 4629 9979
rect 4304 9948 4629 9976
rect 4304 9936 4310 9948
rect 4617 9945 4629 9948
rect 4663 9945 4675 9979
rect 4617 9939 4675 9945
rect 4982 9936 4988 9988
rect 5040 9976 5046 9988
rect 5644 9976 5672 10016
rect 5813 10013 5825 10016
rect 5859 10013 5871 10047
rect 5813 10007 5871 10013
rect 5905 10047 5963 10053
rect 5905 10013 5917 10047
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 5040 9948 5672 9976
rect 5040 9936 5046 9948
rect 5718 9936 5724 9988
rect 5776 9976 5782 9988
rect 5776 9948 5821 9976
rect 5776 9936 5782 9948
rect 4338 9908 4344 9920
rect 4172 9880 4344 9908
rect 4065 9871 4123 9877
rect 4338 9868 4344 9880
rect 4396 9868 4402 9920
rect 5077 9911 5135 9917
rect 5077 9877 5089 9911
rect 5123 9908 5135 9911
rect 5350 9908 5356 9920
rect 5123 9880 5356 9908
rect 5123 9877 5135 9880
rect 5077 9871 5135 9877
rect 5350 9868 5356 9880
rect 5408 9868 5414 9920
rect 5920 9908 5948 10007
rect 6012 9976 6040 10084
rect 6454 10004 6460 10056
rect 6512 10044 6518 10056
rect 6748 10053 6776 10084
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 8110 10112 8116 10124
rect 6972 10084 8116 10112
rect 6972 10072 6978 10084
rect 8110 10072 8116 10084
rect 8168 10072 8174 10124
rect 9508 10112 9536 10220
rect 11517 10217 11529 10220
rect 11563 10248 11575 10251
rect 11790 10248 11796 10260
rect 11563 10220 11796 10248
rect 11563 10217 11575 10220
rect 11517 10211 11575 10217
rect 11790 10208 11796 10220
rect 11848 10208 11854 10260
rect 11974 10208 11980 10260
rect 12032 10248 12038 10260
rect 14090 10248 14096 10260
rect 12032 10220 12664 10248
rect 14051 10220 14096 10248
rect 12032 10208 12038 10220
rect 10134 10112 10140 10124
rect 9416 10084 9536 10112
rect 10095 10084 10140 10112
rect 6549 10047 6607 10053
rect 6549 10044 6561 10047
rect 6512 10016 6561 10044
rect 6512 10004 6518 10016
rect 6549 10013 6561 10016
rect 6595 10013 6607 10047
rect 6549 10007 6607 10013
rect 6733 10047 6791 10053
rect 6733 10013 6745 10047
rect 6779 10013 6791 10047
rect 7558 10044 7564 10056
rect 7471 10016 7564 10044
rect 6733 10007 6791 10013
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10044 7987 10047
rect 8294 10044 8300 10056
rect 7975 10016 8300 10044
rect 7975 10013 7987 10016
rect 7929 10007 7987 10013
rect 8294 10004 8300 10016
rect 8352 10004 8358 10056
rect 9214 10044 9220 10056
rect 9175 10016 9220 10044
rect 9214 10004 9220 10016
rect 9272 10004 9278 10056
rect 9416 10053 9444 10084
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 12158 10072 12164 10124
rect 12216 10112 12222 10124
rect 12437 10115 12495 10121
rect 12437 10112 12449 10115
rect 12216 10084 12449 10112
rect 12216 10072 12222 10084
rect 12437 10081 12449 10084
rect 12483 10081 12495 10115
rect 12636 10112 12664 10220
rect 14090 10208 14096 10220
rect 14148 10208 14154 10260
rect 14182 10208 14188 10260
rect 14240 10248 14246 10260
rect 16390 10248 16396 10260
rect 14240 10220 15976 10248
rect 16351 10220 16396 10248
rect 14240 10208 14246 10220
rect 12710 10140 12716 10192
rect 12768 10180 12774 10192
rect 12897 10183 12955 10189
rect 12897 10180 12909 10183
rect 12768 10152 12909 10180
rect 12768 10140 12774 10152
rect 12897 10149 12909 10152
rect 12943 10149 12955 10183
rect 15948 10180 15976 10220
rect 16390 10208 16396 10220
rect 16448 10208 16454 10260
rect 17221 10251 17279 10257
rect 17221 10217 17233 10251
rect 17267 10248 17279 10251
rect 18230 10248 18236 10260
rect 17267 10220 18236 10248
rect 17267 10217 17279 10220
rect 17221 10211 17279 10217
rect 18230 10208 18236 10220
rect 18288 10208 18294 10260
rect 18414 10208 18420 10260
rect 18472 10248 18478 10260
rect 18601 10251 18659 10257
rect 18601 10248 18613 10251
rect 18472 10220 18613 10248
rect 18472 10208 18478 10220
rect 18601 10217 18613 10220
rect 18647 10217 18659 10251
rect 18601 10211 18659 10217
rect 19518 10208 19524 10260
rect 19576 10248 19582 10260
rect 19797 10251 19855 10257
rect 19797 10248 19809 10251
rect 19576 10220 19809 10248
rect 19576 10208 19582 10220
rect 19797 10217 19809 10220
rect 19843 10217 19855 10251
rect 19797 10211 19855 10217
rect 20349 10251 20407 10257
rect 20349 10217 20361 10251
rect 20395 10248 20407 10251
rect 20438 10248 20444 10260
rect 20395 10220 20444 10248
rect 20395 10217 20407 10220
rect 20349 10211 20407 10217
rect 20438 10208 20444 10220
rect 20496 10208 20502 10260
rect 20993 10251 21051 10257
rect 20993 10217 21005 10251
rect 21039 10248 21051 10251
rect 22462 10248 22468 10260
rect 21039 10220 22468 10248
rect 21039 10217 21051 10220
rect 20993 10211 21051 10217
rect 22462 10208 22468 10220
rect 22520 10208 22526 10260
rect 22922 10208 22928 10260
rect 22980 10248 22986 10260
rect 25133 10251 25191 10257
rect 25133 10248 25145 10251
rect 22980 10220 25145 10248
rect 22980 10208 22986 10220
rect 25133 10217 25145 10220
rect 25179 10217 25191 10251
rect 25133 10211 25191 10217
rect 15948 10152 22094 10180
rect 12897 10143 12955 10149
rect 12912 10112 12940 10143
rect 14642 10112 14648 10124
rect 12636 10084 12756 10112
rect 12912 10084 14648 10112
rect 12437 10075 12495 10081
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10013 9459 10047
rect 9401 10007 9459 10013
rect 9493 10047 9551 10053
rect 9493 10013 9505 10047
rect 9539 10044 9551 10047
rect 9674 10044 9680 10056
rect 9539 10016 9680 10044
rect 9539 10013 9551 10016
rect 9493 10007 9551 10013
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 10404 10047 10462 10053
rect 10404 10013 10416 10047
rect 10450 10044 10462 10047
rect 10962 10044 10968 10056
rect 10450 10016 10968 10044
rect 10450 10013 10462 10016
rect 10404 10007 10462 10013
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 11330 10004 11336 10056
rect 11388 10044 11394 10056
rect 12621 10047 12679 10053
rect 12621 10044 12633 10047
rect 11388 10016 12633 10044
rect 11388 10004 11394 10016
rect 12621 10013 12633 10016
rect 12667 10013 12679 10047
rect 12728 10044 12756 10084
rect 14642 10072 14648 10084
rect 14700 10072 14706 10124
rect 15010 10112 15016 10124
rect 14971 10084 15016 10112
rect 15010 10072 15016 10084
rect 15068 10072 15074 10124
rect 16114 10072 16120 10124
rect 16172 10112 16178 10124
rect 22066 10112 22094 10152
rect 23658 10140 23664 10192
rect 23716 10180 23722 10192
rect 23845 10183 23903 10189
rect 23845 10180 23857 10183
rect 23716 10152 23857 10180
rect 23716 10140 23722 10152
rect 23845 10149 23857 10152
rect 23891 10180 23903 10183
rect 24762 10180 24768 10192
rect 23891 10152 24768 10180
rect 23891 10149 23903 10152
rect 23845 10143 23903 10149
rect 24762 10140 24768 10152
rect 24820 10180 24826 10192
rect 24820 10152 26004 10180
rect 24820 10140 24826 10152
rect 25976 10121 26004 10152
rect 25961 10115 26019 10121
rect 16172 10084 21772 10112
rect 22066 10084 24164 10112
rect 16172 10072 16178 10084
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 12728 10016 14105 10044
rect 12621 10007 12679 10013
rect 14093 10013 14105 10016
rect 14139 10013 14151 10047
rect 14093 10007 14151 10013
rect 14274 10004 14280 10056
rect 14332 10044 14338 10056
rect 15286 10053 15292 10056
rect 14369 10047 14427 10053
rect 14369 10044 14381 10047
rect 14332 10016 14381 10044
rect 14332 10004 14338 10016
rect 14369 10013 14381 10016
rect 14415 10013 14427 10047
rect 15280 10044 15292 10053
rect 15247 10016 15292 10044
rect 14369 10007 14427 10013
rect 15280 10007 15292 10016
rect 15286 10004 15292 10007
rect 15344 10004 15350 10056
rect 16482 10004 16488 10056
rect 16540 10044 16546 10056
rect 16853 10047 16911 10053
rect 16853 10044 16865 10047
rect 16540 10016 16865 10044
rect 16540 10004 16546 10016
rect 16853 10013 16865 10016
rect 16899 10013 16911 10047
rect 16853 10007 16911 10013
rect 17037 10047 17095 10053
rect 17037 10013 17049 10047
rect 17083 10013 17095 10047
rect 17037 10007 17095 10013
rect 7576 9976 7604 10004
rect 6012 9948 7604 9976
rect 7745 9979 7803 9985
rect 7745 9945 7757 9979
rect 7791 9945 7803 9979
rect 7745 9939 7803 9945
rect 6546 9908 6552 9920
rect 5920 9880 6552 9908
rect 6546 9868 6552 9880
rect 6604 9868 6610 9920
rect 6917 9911 6975 9917
rect 6917 9877 6929 9911
rect 6963 9908 6975 9911
rect 7006 9908 7012 9920
rect 6963 9880 7012 9908
rect 6963 9877 6975 9880
rect 6917 9871 6975 9877
rect 7006 9868 7012 9880
rect 7064 9868 7070 9920
rect 7558 9868 7564 9920
rect 7616 9908 7622 9920
rect 7760 9908 7788 9939
rect 7834 9936 7840 9988
rect 7892 9976 7898 9988
rect 7892 9948 7937 9976
rect 10888 9948 12011 9976
rect 7892 9936 7898 9948
rect 7616 9880 7788 9908
rect 7616 9868 7622 9880
rect 8478 9868 8484 9920
rect 8536 9908 8542 9920
rect 9033 9911 9091 9917
rect 9033 9908 9045 9911
rect 8536 9880 9045 9908
rect 8536 9868 8542 9880
rect 9033 9877 9045 9880
rect 9079 9877 9091 9911
rect 9033 9871 9091 9877
rect 9490 9868 9496 9920
rect 9548 9908 9554 9920
rect 10888 9908 10916 9948
rect 9548 9880 10916 9908
rect 9548 9868 9554 9880
rect 10962 9868 10968 9920
rect 11020 9908 11026 9920
rect 11882 9908 11888 9920
rect 11020 9880 11888 9908
rect 11020 9868 11026 9880
rect 11882 9868 11888 9880
rect 11940 9868 11946 9920
rect 11983 9908 12011 9948
rect 12250 9936 12256 9988
rect 12308 9976 12314 9988
rect 12989 9979 13047 9985
rect 12989 9976 13001 9979
rect 12308 9948 13001 9976
rect 12308 9936 12314 9948
rect 12989 9945 13001 9948
rect 13035 9945 13047 9979
rect 12989 9939 13047 9945
rect 12526 9908 12532 9920
rect 11983 9880 12532 9908
rect 12526 9868 12532 9880
rect 12584 9868 12590 9920
rect 13004 9908 13032 9939
rect 13078 9936 13084 9988
rect 13136 9976 13142 9988
rect 13136 9948 14412 9976
rect 13136 9936 13142 9948
rect 13906 9908 13912 9920
rect 13004 9880 13912 9908
rect 13906 9868 13912 9880
rect 13964 9868 13970 9920
rect 14182 9868 14188 9920
rect 14240 9908 14246 9920
rect 14277 9911 14335 9917
rect 14277 9908 14289 9911
rect 14240 9880 14289 9908
rect 14240 9868 14246 9880
rect 14277 9877 14289 9880
rect 14323 9877 14335 9911
rect 14384 9908 14412 9948
rect 15654 9936 15660 9988
rect 15712 9976 15718 9988
rect 17052 9976 17080 10007
rect 17310 10004 17316 10056
rect 17368 10044 17374 10056
rect 17586 10044 17592 10056
rect 17368 10016 17592 10044
rect 17368 10004 17374 10016
rect 17586 10004 17592 10016
rect 17644 10004 17650 10056
rect 17678 10004 17684 10056
rect 17736 10004 17742 10056
rect 17862 10044 17868 10056
rect 17823 10016 17868 10044
rect 17862 10004 17868 10016
rect 17920 10004 17926 10056
rect 18524 10053 18552 10084
rect 18509 10047 18567 10053
rect 18509 10013 18521 10047
rect 18555 10013 18567 10047
rect 18509 10007 18567 10013
rect 19245 10047 19303 10053
rect 19245 10013 19257 10047
rect 19291 10013 19303 10047
rect 19245 10007 19303 10013
rect 15712 9948 17080 9976
rect 17696 9976 17724 10004
rect 18598 9976 18604 9988
rect 17696 9948 18604 9976
rect 15712 9936 15718 9948
rect 18598 9936 18604 9948
rect 18656 9936 18662 9988
rect 19260 9976 19288 10007
rect 19334 10004 19340 10056
rect 19392 10044 19398 10056
rect 19613 10047 19671 10053
rect 19613 10044 19625 10047
rect 19392 10016 19625 10044
rect 19392 10004 19398 10016
rect 19613 10013 19625 10016
rect 19659 10013 19671 10047
rect 19613 10007 19671 10013
rect 20533 10047 20591 10053
rect 20533 10013 20545 10047
rect 20579 10044 20591 10047
rect 20898 10044 20904 10056
rect 20579 10016 20904 10044
rect 20579 10013 20591 10016
rect 20533 10007 20591 10013
rect 20898 10004 20904 10016
rect 20956 10004 20962 10056
rect 21744 10053 21772 10084
rect 21177 10047 21235 10053
rect 21177 10013 21189 10047
rect 21223 10013 21235 10047
rect 21177 10007 21235 10013
rect 21729 10047 21787 10053
rect 21729 10013 21741 10047
rect 21775 10013 21787 10047
rect 21729 10007 21787 10013
rect 21913 10047 21971 10053
rect 21913 10013 21925 10047
rect 21959 10044 21971 10047
rect 23106 10044 23112 10056
rect 21959 10016 23112 10044
rect 21959 10013 21971 10016
rect 21913 10007 21971 10013
rect 19426 9976 19432 9988
rect 19260 9948 19334 9976
rect 19387 9948 19432 9976
rect 16390 9908 16396 9920
rect 14384 9880 16396 9908
rect 14277 9871 14335 9877
rect 16390 9868 16396 9880
rect 16448 9868 16454 9920
rect 17586 9868 17592 9920
rect 17644 9908 17650 9920
rect 17681 9911 17739 9917
rect 17681 9908 17693 9911
rect 17644 9880 17693 9908
rect 17644 9868 17650 9880
rect 17681 9877 17693 9880
rect 17727 9877 17739 9911
rect 19306 9908 19334 9948
rect 19426 9936 19432 9948
rect 19484 9936 19490 9988
rect 19521 9979 19579 9985
rect 19521 9945 19533 9979
rect 19567 9976 19579 9979
rect 20990 9976 20996 9988
rect 19567 9948 20996 9976
rect 19567 9945 19579 9948
rect 19521 9939 19579 9945
rect 20990 9936 20996 9948
rect 21048 9936 21054 9988
rect 20714 9908 20720 9920
rect 19306 9880 20720 9908
rect 17681 9871 17739 9877
rect 20714 9868 20720 9880
rect 20772 9868 20778 9920
rect 21192 9908 21220 10007
rect 23106 10004 23112 10016
rect 23164 10044 23170 10056
rect 23661 10047 23719 10053
rect 23661 10044 23673 10047
rect 23164 10016 23673 10044
rect 23164 10004 23170 10016
rect 23661 10013 23673 10016
rect 23707 10013 23719 10047
rect 23661 10007 23719 10013
rect 22738 9976 22744 9988
rect 22699 9948 22744 9976
rect 22738 9936 22744 9948
rect 22796 9936 22802 9988
rect 22646 9908 22652 9920
rect 21192 9880 22652 9908
rect 22646 9868 22652 9880
rect 22704 9868 22710 9920
rect 22833 9911 22891 9917
rect 22833 9877 22845 9911
rect 22879 9908 22891 9911
rect 23290 9908 23296 9920
rect 22879 9880 23296 9908
rect 22879 9877 22891 9880
rect 22833 9871 22891 9877
rect 23290 9868 23296 9880
rect 23348 9868 23354 9920
rect 24136 9908 24164 10084
rect 25961 10081 25973 10115
rect 26007 10081 26019 10115
rect 25961 10075 26019 10081
rect 24210 10004 24216 10056
rect 24268 10044 24274 10056
rect 24397 10047 24455 10053
rect 24397 10044 24409 10047
rect 24268 10016 24409 10044
rect 24268 10004 24274 10016
rect 24397 10013 24409 10016
rect 24443 10013 24455 10047
rect 24397 10007 24455 10013
rect 24670 10004 24676 10056
rect 24728 10044 24734 10056
rect 25317 10047 25375 10053
rect 25317 10044 25329 10047
rect 24728 10016 25329 10044
rect 24728 10004 24734 10016
rect 25317 10013 25329 10016
rect 25363 10013 25375 10047
rect 25317 10007 25375 10013
rect 26228 9979 26286 9985
rect 26228 9945 26240 9979
rect 26274 9976 26286 9979
rect 26694 9976 26700 9988
rect 26274 9948 26700 9976
rect 26274 9945 26286 9948
rect 26228 9939 26286 9945
rect 26694 9936 26700 9948
rect 26752 9936 26758 9988
rect 24581 9911 24639 9917
rect 24581 9908 24593 9911
rect 24136 9880 24593 9908
rect 24581 9877 24593 9880
rect 24627 9908 24639 9911
rect 25774 9908 25780 9920
rect 24627 9880 25780 9908
rect 24627 9877 24639 9880
rect 24581 9871 24639 9877
rect 25774 9868 25780 9880
rect 25832 9868 25838 9920
rect 26878 9868 26884 9920
rect 26936 9908 26942 9920
rect 27341 9911 27399 9917
rect 27341 9908 27353 9911
rect 26936 9880 27353 9908
rect 26936 9868 26942 9880
rect 27341 9877 27353 9880
rect 27387 9877 27399 9911
rect 27341 9871 27399 9877
rect 1104 9818 28060 9840
rect 1104 9766 9935 9818
rect 9987 9766 9999 9818
rect 10051 9766 10063 9818
rect 10115 9766 10127 9818
rect 10179 9766 10191 9818
rect 10243 9766 18920 9818
rect 18972 9766 18984 9818
rect 19036 9766 19048 9818
rect 19100 9766 19112 9818
rect 19164 9766 19176 9818
rect 19228 9766 28060 9818
rect 1104 9744 28060 9766
rect 1578 9664 1584 9716
rect 1636 9704 1642 9716
rect 8110 9704 8116 9716
rect 1636 9676 8116 9704
rect 1636 9664 1642 9676
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 9030 9664 9036 9716
rect 9088 9704 9094 9716
rect 9490 9704 9496 9716
rect 9088 9676 9496 9704
rect 9088 9664 9094 9676
rect 9490 9664 9496 9676
rect 9548 9664 9554 9716
rect 11882 9704 11888 9716
rect 10612 9676 11100 9704
rect 2032 9639 2090 9645
rect 2032 9605 2044 9639
rect 2078 9636 2090 9639
rect 2222 9636 2228 9648
rect 2078 9608 2228 9636
rect 2078 9605 2090 9608
rect 2032 9599 2090 9605
rect 2222 9596 2228 9608
rect 2280 9596 2286 9648
rect 4338 9596 4344 9648
rect 4396 9636 4402 9648
rect 4396 9608 5672 9636
rect 4396 9596 4402 9608
rect 3326 9528 3332 9580
rect 3384 9568 3390 9580
rect 4137 9571 4195 9577
rect 4137 9568 4149 9571
rect 3384 9540 4149 9568
rect 3384 9528 3390 9540
rect 4137 9537 4149 9540
rect 4183 9537 4195 9571
rect 4137 9531 4195 9537
rect 1578 9460 1584 9512
rect 1636 9500 1642 9512
rect 1765 9503 1823 9509
rect 1765 9500 1777 9503
rect 1636 9472 1777 9500
rect 1636 9460 1642 9472
rect 1765 9469 1777 9472
rect 1811 9469 1823 9503
rect 1765 9463 1823 9469
rect 3786 9460 3792 9512
rect 3844 9500 3850 9512
rect 3881 9503 3939 9509
rect 3881 9500 3893 9503
rect 3844 9472 3893 9500
rect 3844 9460 3850 9472
rect 3881 9469 3893 9472
rect 3927 9469 3939 9503
rect 3881 9463 3939 9469
rect 5534 9392 5540 9444
rect 5592 9392 5598 9444
rect 5644 9432 5672 9608
rect 5718 9596 5724 9648
rect 5776 9636 5782 9648
rect 6638 9636 6644 9648
rect 5776 9608 6644 9636
rect 5776 9596 5782 9608
rect 6638 9596 6644 9608
rect 6696 9596 6702 9648
rect 7558 9596 7564 9648
rect 7616 9636 7622 9648
rect 10612 9645 10640 9676
rect 10597 9639 10655 9645
rect 10597 9636 10609 9639
rect 7616 9608 10609 9636
rect 7616 9596 7622 9608
rect 10597 9605 10609 9608
rect 10643 9605 10655 9639
rect 10597 9599 10655 9605
rect 10689 9639 10747 9645
rect 10689 9605 10701 9639
rect 10735 9636 10747 9639
rect 10962 9636 10968 9648
rect 10735 9608 10968 9636
rect 10735 9605 10747 9608
rect 10689 9599 10747 9605
rect 10962 9596 10968 9608
rect 11020 9596 11026 9648
rect 11072 9636 11100 9676
rect 11716 9676 11888 9704
rect 11716 9636 11744 9676
rect 11882 9664 11888 9676
rect 11940 9664 11946 9716
rect 12912 9676 15240 9704
rect 11072 9608 11744 9636
rect 11790 9596 11796 9648
rect 11848 9636 11854 9648
rect 12161 9639 12219 9645
rect 12161 9636 12173 9639
rect 11848 9608 12173 9636
rect 11848 9596 11854 9608
rect 12161 9605 12173 9608
rect 12207 9605 12219 9639
rect 12161 9599 12219 9605
rect 6546 9528 6552 9580
rect 6604 9568 6610 9580
rect 7009 9571 7067 9577
rect 7009 9568 7021 9571
rect 6604 9540 7021 9568
rect 6604 9528 6610 9540
rect 7009 9537 7021 9540
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 7834 9528 7840 9580
rect 7892 9568 7898 9580
rect 8113 9571 8171 9577
rect 8113 9568 8125 9571
rect 7892 9540 8125 9568
rect 7892 9528 7898 9540
rect 8113 9537 8125 9540
rect 8159 9537 8171 9571
rect 8113 9531 8171 9537
rect 8478 9528 8484 9580
rect 8536 9568 8542 9580
rect 8757 9571 8815 9577
rect 8757 9568 8769 9571
rect 8536 9540 8769 9568
rect 8536 9528 8542 9540
rect 8757 9537 8769 9540
rect 8803 9537 8815 9571
rect 8757 9531 8815 9537
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9568 9091 9571
rect 9398 9568 9404 9580
rect 9079 9540 9404 9568
rect 9079 9537 9091 9540
rect 9033 9531 9091 9537
rect 9398 9528 9404 9540
rect 9456 9528 9462 9580
rect 9490 9528 9496 9580
rect 9548 9568 9554 9580
rect 9769 9571 9827 9577
rect 9769 9568 9781 9571
rect 9548 9540 9781 9568
rect 9548 9528 9554 9540
rect 9769 9537 9781 9540
rect 9815 9537 9827 9571
rect 9769 9531 9827 9537
rect 9858 9528 9864 9580
rect 9916 9568 9922 9580
rect 10413 9571 10471 9577
rect 10413 9568 10425 9571
rect 9916 9540 10425 9568
rect 9916 9528 9922 9540
rect 10413 9537 10425 9540
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 6733 9503 6791 9509
rect 6733 9469 6745 9503
rect 6779 9500 6791 9503
rect 7852 9500 7880 9528
rect 8294 9500 8300 9512
rect 6779 9472 7880 9500
rect 8207 9472 8300 9500
rect 6779 9469 6791 9472
rect 6733 9463 6791 9469
rect 8294 9460 8300 9472
rect 8352 9500 8358 9512
rect 10796 9500 10824 9531
rect 11054 9528 11060 9580
rect 11112 9568 11118 9580
rect 11977 9571 12035 9577
rect 11977 9568 11989 9571
rect 11112 9540 11989 9568
rect 11112 9528 11118 9540
rect 11977 9537 11989 9540
rect 12023 9537 12035 9571
rect 12912 9568 12940 9676
rect 15105 9639 15163 9645
rect 15105 9636 15117 9639
rect 11977 9531 12035 9537
rect 12084 9540 12940 9568
rect 13004 9608 15117 9636
rect 12084 9500 12112 9540
rect 8352 9472 12112 9500
rect 8352 9460 8358 9472
rect 12158 9460 12164 9512
rect 12216 9500 12222 9512
rect 13004 9500 13032 9608
rect 15105 9605 15117 9608
rect 15151 9605 15163 9639
rect 15212 9636 15240 9676
rect 17034 9664 17040 9716
rect 17092 9704 17098 9716
rect 17678 9704 17684 9716
rect 17092 9676 17684 9704
rect 17092 9664 17098 9676
rect 17678 9664 17684 9676
rect 17736 9664 17742 9716
rect 17770 9664 17776 9716
rect 17828 9704 17834 9716
rect 19518 9704 19524 9716
rect 17828 9676 18828 9704
rect 17828 9664 17834 9676
rect 16666 9636 16672 9648
rect 15212 9608 16672 9636
rect 15105 9599 15163 9605
rect 16666 9596 16672 9608
rect 16724 9596 16730 9648
rect 18800 9645 18828 9676
rect 18892 9676 19524 9704
rect 18892 9645 18920 9676
rect 19518 9664 19524 9676
rect 19576 9664 19582 9716
rect 23201 9707 23259 9713
rect 23201 9673 23213 9707
rect 23247 9673 23259 9707
rect 23201 9667 23259 9673
rect 18785 9639 18843 9645
rect 18432 9608 18700 9636
rect 13440 9571 13498 9577
rect 13440 9537 13452 9571
rect 13486 9568 13498 9571
rect 13486 9540 14596 9568
rect 13486 9537 13498 9540
rect 13440 9531 13498 9537
rect 13170 9500 13176 9512
rect 12216 9472 13032 9500
rect 13131 9472 13176 9500
rect 12216 9460 12222 9472
rect 13170 9460 13176 9472
rect 13228 9460 13234 9512
rect 14568 9500 14596 9540
rect 14642 9528 14648 9580
rect 14700 9568 14706 9580
rect 15013 9571 15071 9577
rect 15013 9568 15025 9571
rect 14700 9540 15025 9568
rect 14700 9528 14706 9540
rect 15013 9537 15025 9540
rect 15059 9537 15071 9571
rect 15838 9568 15844 9580
rect 15799 9540 15844 9568
rect 15013 9531 15071 9537
rect 15838 9528 15844 9540
rect 15896 9528 15902 9580
rect 16853 9571 16911 9577
rect 16853 9537 16865 9571
rect 16899 9568 16911 9571
rect 17034 9568 17040 9580
rect 16899 9540 17040 9568
rect 16899 9537 16911 9540
rect 16853 9531 16911 9537
rect 17034 9528 17040 9540
rect 17092 9528 17098 9580
rect 18049 9571 18107 9577
rect 18049 9537 18061 9571
rect 18095 9568 18107 9571
rect 18230 9568 18236 9580
rect 18095 9540 18236 9568
rect 18095 9537 18107 9540
rect 18049 9531 18107 9537
rect 18230 9528 18236 9540
rect 18288 9528 18294 9580
rect 14568 9472 15700 9500
rect 5644 9404 8340 9432
rect 2958 9324 2964 9376
rect 3016 9364 3022 9376
rect 3145 9367 3203 9373
rect 3145 9364 3157 9367
rect 3016 9336 3157 9364
rect 3016 9324 3022 9336
rect 3145 9333 3157 9336
rect 3191 9364 3203 9367
rect 4246 9364 4252 9376
rect 3191 9336 4252 9364
rect 3191 9333 3203 9336
rect 3145 9327 3203 9333
rect 4246 9324 4252 9336
rect 4304 9324 4310 9376
rect 5261 9367 5319 9373
rect 5261 9333 5273 9367
rect 5307 9364 5319 9367
rect 5552 9364 5580 9392
rect 5810 9364 5816 9376
rect 5307 9336 5816 9364
rect 5307 9333 5319 9336
rect 5261 9327 5319 9333
rect 5810 9324 5816 9336
rect 5868 9324 5874 9376
rect 8312 9364 8340 9404
rect 8386 9392 8392 9444
rect 8444 9432 8450 9444
rect 10226 9432 10232 9444
rect 8444 9404 10232 9432
rect 8444 9392 8450 9404
rect 8849 9367 8907 9373
rect 8849 9364 8861 9367
rect 8312 9336 8861 9364
rect 8849 9333 8861 9336
rect 8895 9364 8907 9367
rect 9030 9364 9036 9376
rect 8895 9336 9036 9364
rect 8895 9333 8907 9336
rect 8849 9327 8907 9333
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 9876 9373 9904 9404
rect 10226 9392 10232 9404
rect 10284 9392 10290 9444
rect 10502 9392 10508 9444
rect 10560 9432 10566 9444
rect 10965 9435 11023 9441
rect 10965 9432 10977 9435
rect 10560 9404 10977 9432
rect 10560 9392 10566 9404
rect 10965 9401 10977 9404
rect 11011 9401 11023 9435
rect 12250 9432 12256 9444
rect 10965 9395 11023 9401
rect 11072 9404 12256 9432
rect 9861 9367 9919 9373
rect 9861 9333 9873 9367
rect 9907 9333 9919 9367
rect 9861 9327 9919 9333
rect 9950 9324 9956 9376
rect 10008 9364 10014 9376
rect 11072 9364 11100 9404
rect 12250 9392 12256 9404
rect 12308 9392 12314 9444
rect 12526 9432 12532 9444
rect 12406 9404 12532 9432
rect 10008 9336 11100 9364
rect 10008 9324 10014 9336
rect 11146 9324 11152 9376
rect 11204 9364 11210 9376
rect 12406 9364 12434 9404
rect 12526 9392 12532 9404
rect 12584 9392 12590 9444
rect 15672 9441 15700 9472
rect 16666 9460 16672 9512
rect 16724 9500 16730 9512
rect 16942 9500 16948 9512
rect 16724 9472 16948 9500
rect 16724 9460 16730 9472
rect 16942 9460 16948 9472
rect 17000 9460 17006 9512
rect 15657 9435 15715 9441
rect 14476 9404 15608 9432
rect 11204 9336 12434 9364
rect 11204 9324 11210 9336
rect 12894 9324 12900 9376
rect 12952 9364 12958 9376
rect 14476 9364 14504 9404
rect 12952 9336 14504 9364
rect 14553 9367 14611 9373
rect 12952 9324 12958 9336
rect 14553 9333 14565 9367
rect 14599 9364 14611 9367
rect 14826 9364 14832 9376
rect 14599 9336 14832 9364
rect 14599 9333 14611 9336
rect 14553 9327 14611 9333
rect 14826 9324 14832 9336
rect 14884 9324 14890 9376
rect 15580 9364 15608 9404
rect 15657 9401 15669 9435
rect 15703 9401 15715 9435
rect 17770 9432 17776 9444
rect 15657 9395 15715 9401
rect 16546 9404 17776 9432
rect 16546 9364 16574 9404
rect 17770 9392 17776 9404
rect 17828 9392 17834 9444
rect 15580 9336 16574 9364
rect 16669 9367 16727 9373
rect 16669 9333 16681 9367
rect 16715 9364 16727 9367
rect 16942 9364 16948 9376
rect 16715 9336 16948 9364
rect 16715 9333 16727 9336
rect 16669 9327 16727 9333
rect 16942 9324 16948 9336
rect 17000 9324 17006 9376
rect 17865 9367 17923 9373
rect 17865 9333 17877 9367
rect 17911 9364 17923 9367
rect 18046 9364 18052 9376
rect 17911 9336 18052 9364
rect 17911 9333 17923 9336
rect 17865 9327 17923 9333
rect 18046 9324 18052 9336
rect 18104 9324 18110 9376
rect 18432 9364 18460 9608
rect 18672 9577 18700 9608
rect 18785 9605 18797 9639
rect 18831 9605 18843 9639
rect 18785 9599 18843 9605
rect 18873 9639 18931 9645
rect 18873 9605 18885 9639
rect 18919 9605 18931 9639
rect 19334 9636 19340 9648
rect 18873 9599 18931 9605
rect 19076 9608 19340 9636
rect 18647 9571 18705 9577
rect 18647 9537 18659 9571
rect 18693 9537 18705 9571
rect 18647 9531 18705 9537
rect 18969 9571 19027 9577
rect 18969 9537 18981 9571
rect 19015 9558 19027 9571
rect 19076 9558 19104 9608
rect 19334 9596 19340 9608
rect 19392 9596 19398 9648
rect 23216 9636 23244 9667
rect 23290 9664 23296 9716
rect 23348 9704 23354 9716
rect 27338 9704 27344 9716
rect 23348 9676 27344 9704
rect 23348 9664 23354 9676
rect 25222 9636 25228 9648
rect 19444 9608 25228 9636
rect 19015 9537 19104 9558
rect 18969 9531 19104 9537
rect 18984 9530 19104 9531
rect 19444 9432 19472 9608
rect 25222 9596 25228 9608
rect 25280 9596 25286 9648
rect 19518 9528 19524 9580
rect 19576 9568 19582 9580
rect 19613 9571 19671 9577
rect 19613 9568 19625 9571
rect 19576 9540 19625 9568
rect 19576 9528 19582 9540
rect 19613 9537 19625 9540
rect 19659 9537 19671 9571
rect 19794 9568 19800 9580
rect 19755 9540 19800 9568
rect 19613 9531 19671 9537
rect 19794 9528 19800 9540
rect 19852 9528 19858 9580
rect 19886 9528 19892 9580
rect 19944 9568 19950 9580
rect 20625 9571 20683 9577
rect 20625 9568 20637 9571
rect 19944 9540 20637 9568
rect 19944 9528 19950 9540
rect 20625 9537 20637 9540
rect 20671 9568 20683 9571
rect 20714 9568 20720 9580
rect 20671 9540 20720 9568
rect 20671 9537 20683 9540
rect 20625 9531 20683 9537
rect 20714 9528 20720 9540
rect 20772 9528 20778 9580
rect 21266 9568 21272 9580
rect 21227 9540 21272 9568
rect 21266 9528 21272 9540
rect 21324 9528 21330 9580
rect 22094 9577 22100 9580
rect 22088 9531 22100 9577
rect 22152 9568 22158 9580
rect 23658 9568 23664 9580
rect 22152 9540 22188 9568
rect 23619 9540 23664 9568
rect 22094 9528 22100 9531
rect 22152 9528 22158 9540
rect 23658 9528 23664 9540
rect 23716 9528 23722 9580
rect 25700 9577 25728 9676
rect 27338 9664 27344 9676
rect 27396 9664 27402 9716
rect 25869 9639 25927 9645
rect 25869 9605 25881 9639
rect 25915 9636 25927 9639
rect 26418 9636 26424 9648
rect 25915 9608 26424 9636
rect 25915 9605 25927 9608
rect 25869 9599 25927 9605
rect 26418 9596 26424 9608
rect 26476 9596 26482 9648
rect 23928 9571 23986 9577
rect 23928 9537 23940 9571
rect 23974 9568 23986 9571
rect 25685 9571 25743 9577
rect 23974 9540 25544 9568
rect 23974 9537 23986 9540
rect 23928 9531 23986 9537
rect 19981 9503 20039 9509
rect 19981 9469 19993 9503
rect 20027 9500 20039 9503
rect 20806 9500 20812 9512
rect 20027 9472 20812 9500
rect 20027 9469 20039 9472
rect 19981 9463 20039 9469
rect 20806 9460 20812 9472
rect 20864 9460 20870 9512
rect 21821 9503 21879 9509
rect 21821 9469 21833 9503
rect 21867 9469 21879 9503
rect 21821 9463 21879 9469
rect 18672 9404 19472 9432
rect 18672 9364 18700 9404
rect 18432 9336 18700 9364
rect 19153 9367 19211 9373
rect 19153 9333 19165 9367
rect 19199 9364 19211 9367
rect 19702 9364 19708 9376
rect 19199 9336 19708 9364
rect 19199 9333 19211 9336
rect 19153 9327 19211 9333
rect 19702 9324 19708 9336
rect 19760 9324 19766 9376
rect 20438 9364 20444 9376
rect 20399 9336 20444 9364
rect 20438 9324 20444 9336
rect 20496 9324 20502 9376
rect 21085 9367 21143 9373
rect 21085 9333 21097 9367
rect 21131 9364 21143 9367
rect 21358 9364 21364 9376
rect 21131 9336 21364 9364
rect 21131 9333 21143 9336
rect 21085 9327 21143 9333
rect 21358 9324 21364 9336
rect 21416 9324 21422 9376
rect 21836 9364 21864 9463
rect 23658 9392 23664 9444
rect 23716 9392 23722 9444
rect 24854 9392 24860 9444
rect 24912 9432 24918 9444
rect 25314 9432 25320 9444
rect 24912 9404 25320 9432
rect 24912 9392 24918 9404
rect 25314 9392 25320 9404
rect 25372 9392 25378 9444
rect 25516 9432 25544 9540
rect 25685 9537 25697 9571
rect 25731 9537 25743 9571
rect 25685 9531 25743 9537
rect 25774 9528 25780 9580
rect 25832 9568 25838 9580
rect 25961 9571 26019 9577
rect 25961 9568 25973 9571
rect 25832 9540 25973 9568
rect 25832 9528 25838 9540
rect 25961 9537 25973 9540
rect 26007 9537 26019 9571
rect 25961 9531 26019 9537
rect 25976 9500 26004 9531
rect 26050 9528 26056 9580
rect 26108 9568 26114 9580
rect 27065 9571 27123 9577
rect 27065 9568 27077 9571
rect 26108 9540 27077 9568
rect 26108 9528 26114 9540
rect 27065 9537 27077 9540
rect 27111 9537 27123 9571
rect 27065 9531 27123 9537
rect 27154 9500 27160 9512
rect 25976 9472 27160 9500
rect 27154 9460 27160 9472
rect 27212 9460 27218 9512
rect 27062 9432 27068 9444
rect 25516 9404 27068 9432
rect 27062 9392 27068 9404
rect 27120 9392 27126 9444
rect 23676 9364 23704 9392
rect 21836 9336 23704 9364
rect 23842 9324 23848 9376
rect 23900 9364 23906 9376
rect 25041 9367 25099 9373
rect 25041 9364 25053 9367
rect 23900 9336 25053 9364
rect 23900 9324 23906 9336
rect 25041 9333 25053 9336
rect 25087 9333 25099 9367
rect 25498 9364 25504 9376
rect 25459 9336 25504 9364
rect 25041 9327 25099 9333
rect 25498 9324 25504 9336
rect 25556 9324 25562 9376
rect 27249 9367 27307 9373
rect 27249 9333 27261 9367
rect 27295 9364 27307 9367
rect 27614 9364 27620 9376
rect 27295 9336 27620 9364
rect 27295 9333 27307 9336
rect 27249 9327 27307 9333
rect 27614 9324 27620 9336
rect 27672 9324 27678 9376
rect 1104 9274 28060 9296
rect 1104 9222 5442 9274
rect 5494 9222 5506 9274
rect 5558 9222 5570 9274
rect 5622 9222 5634 9274
rect 5686 9222 5698 9274
rect 5750 9222 14428 9274
rect 14480 9222 14492 9274
rect 14544 9222 14556 9274
rect 14608 9222 14620 9274
rect 14672 9222 14684 9274
rect 14736 9222 23413 9274
rect 23465 9222 23477 9274
rect 23529 9222 23541 9274
rect 23593 9222 23605 9274
rect 23657 9222 23669 9274
rect 23721 9222 28060 9274
rect 1104 9200 28060 9222
rect 9950 9160 9956 9172
rect 1504 9132 9956 9160
rect 1504 8965 1532 9132
rect 9950 9120 9956 9132
rect 10008 9120 10014 9172
rect 12342 9160 12348 9172
rect 10336 9132 12348 9160
rect 1857 9095 1915 9101
rect 1857 9061 1869 9095
rect 1903 9092 1915 9095
rect 3145 9095 3203 9101
rect 1903 9064 3096 9092
rect 1903 9061 1915 9064
rect 1857 9055 1915 9061
rect 2590 9024 2596 9036
rect 1596 8996 2596 9024
rect 1596 8965 1624 8996
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 2682 8984 2688 9036
rect 2740 9024 2746 9036
rect 3068 9024 3096 9064
rect 3145 9061 3157 9095
rect 3191 9092 3203 9095
rect 3970 9092 3976 9104
rect 3191 9064 3976 9092
rect 3191 9061 3203 9064
rect 3145 9055 3203 9061
rect 3970 9052 3976 9064
rect 4028 9092 4034 9104
rect 5997 9095 6055 9101
rect 4028 9064 4292 9092
rect 4028 9052 4034 9064
rect 4264 9033 4292 9064
rect 5997 9061 6009 9095
rect 6043 9092 6055 9095
rect 7558 9092 7564 9104
rect 6043 9064 7564 9092
rect 6043 9061 6055 9064
rect 5997 9055 6055 9061
rect 7558 9052 7564 9064
rect 7616 9052 7622 9104
rect 4249 9027 4307 9033
rect 2740 8984 2774 9024
rect 3068 8996 3924 9024
rect 1489 8959 1547 8965
rect 1489 8925 1501 8959
rect 1535 8925 1547 8959
rect 1489 8919 1547 8925
rect 1581 8959 1639 8965
rect 1581 8925 1593 8959
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 1762 8956 1768 8968
rect 1719 8928 1768 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 1762 8916 1768 8928
rect 1820 8916 1826 8968
rect 2746 8956 2774 8984
rect 2869 8959 2927 8965
rect 2869 8956 2881 8959
rect 2746 8928 2881 8956
rect 2869 8925 2881 8928
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 2958 8916 2964 8968
rect 3016 8956 3022 8968
rect 3237 8959 3295 8965
rect 3016 8928 3061 8956
rect 3016 8916 3022 8928
rect 3237 8925 3249 8959
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 2314 8848 2320 8900
rect 2372 8888 2378 8900
rect 3252 8888 3280 8919
rect 2372 8860 3280 8888
rect 2372 8848 2378 8860
rect 2590 8780 2596 8832
rect 2648 8820 2654 8832
rect 2685 8823 2743 8829
rect 2685 8820 2697 8823
rect 2648 8792 2697 8820
rect 2648 8780 2654 8792
rect 2685 8789 2697 8792
rect 2731 8789 2743 8823
rect 3896 8820 3924 8996
rect 4249 8993 4261 9027
rect 4295 8993 4307 9027
rect 4249 8987 4307 8993
rect 5902 8984 5908 9036
rect 5960 9024 5966 9036
rect 6457 9027 6515 9033
rect 6457 9024 6469 9027
rect 5960 8996 6469 9024
rect 5960 8984 5966 8996
rect 6457 8993 6469 8996
rect 6503 8993 6515 9027
rect 6457 8987 6515 8993
rect 6638 8984 6644 9036
rect 6696 9024 6702 9036
rect 6733 9027 6791 9033
rect 6733 9024 6745 9027
rect 6696 8996 6745 9024
rect 6696 8984 6702 8996
rect 6733 8993 6745 8996
rect 6779 8993 6791 9027
rect 9398 9024 9404 9036
rect 6733 8987 6791 8993
rect 8036 8996 9404 9024
rect 3973 8959 4031 8965
rect 3973 8925 3985 8959
rect 4019 8956 4031 8959
rect 4338 8956 4344 8968
rect 4019 8928 4344 8956
rect 4019 8925 4031 8928
rect 3973 8919 4031 8925
rect 4338 8916 4344 8928
rect 4396 8956 4402 8968
rect 6288 8956 6500 8958
rect 8036 8956 8064 8996
rect 9398 8984 9404 8996
rect 9456 9024 9462 9036
rect 10336 9033 10364 9132
rect 12342 9120 12348 9132
rect 12400 9120 12406 9172
rect 12526 9160 12532 9172
rect 12487 9132 12532 9160
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 13357 9163 13415 9169
rect 13357 9129 13369 9163
rect 13403 9160 13415 9163
rect 15838 9160 15844 9172
rect 13403 9132 15844 9160
rect 13403 9129 13415 9132
rect 13357 9123 13415 9129
rect 15838 9120 15844 9132
rect 15896 9120 15902 9172
rect 15930 9120 15936 9172
rect 15988 9160 15994 9172
rect 17310 9160 17316 9172
rect 15988 9132 17316 9160
rect 15988 9120 15994 9132
rect 17310 9120 17316 9132
rect 17368 9160 17374 9172
rect 18049 9163 18107 9169
rect 18049 9160 18061 9163
rect 17368 9132 18061 9160
rect 17368 9120 17374 9132
rect 18049 9129 18061 9132
rect 18095 9129 18107 9163
rect 18049 9123 18107 9129
rect 18509 9163 18567 9169
rect 18509 9129 18521 9163
rect 18555 9160 18567 9163
rect 19794 9160 19800 9172
rect 18555 9132 19656 9160
rect 19755 9132 19800 9160
rect 18555 9129 18567 9132
rect 18509 9123 18567 9129
rect 13170 9052 13176 9104
rect 13228 9052 13234 9104
rect 18690 9052 18696 9104
rect 18748 9052 18754 9104
rect 19628 9092 19656 9132
rect 19794 9120 19800 9132
rect 19852 9120 19858 9172
rect 20438 9120 20444 9172
rect 20496 9160 20502 9172
rect 20496 9132 21496 9160
rect 20496 9120 20502 9132
rect 20254 9092 20260 9104
rect 19628 9064 20260 9092
rect 20254 9052 20260 9064
rect 20312 9052 20318 9104
rect 9585 9027 9643 9033
rect 9585 9024 9597 9027
rect 9456 8996 9597 9024
rect 9456 8984 9462 8996
rect 9585 8993 9597 8996
rect 9631 8993 9643 9027
rect 9585 8987 9643 8993
rect 10321 9027 10379 9033
rect 10321 8993 10333 9027
rect 10367 8993 10379 9027
rect 10321 8987 10379 8993
rect 12526 8984 12532 9036
rect 12584 9024 12590 9036
rect 12802 9024 12808 9036
rect 12584 8996 12808 9024
rect 12584 8984 12590 8996
rect 12802 8984 12808 8996
rect 12860 9024 12866 9036
rect 12989 9027 13047 9033
rect 12989 9024 13001 9027
rect 12860 8996 13001 9024
rect 12860 8984 12866 8996
rect 12989 8993 13001 8996
rect 13035 8993 13047 9027
rect 13188 9024 13216 9052
rect 14645 9027 14703 9033
rect 14645 9024 14657 9027
rect 13188 8996 14657 9024
rect 12989 8987 13047 8993
rect 14645 8993 14657 8996
rect 14691 8993 14703 9027
rect 18708 9024 18736 9052
rect 21468 9024 21496 9132
rect 21542 9120 21548 9172
rect 21600 9160 21606 9172
rect 26050 9160 26056 9172
rect 21600 9132 26056 9160
rect 21600 9120 21606 9132
rect 26050 9120 26056 9132
rect 26108 9120 26114 9172
rect 26694 9160 26700 9172
rect 26655 9132 26700 9160
rect 26694 9120 26700 9132
rect 26752 9120 26758 9172
rect 21634 9052 21640 9104
rect 21692 9092 21698 9104
rect 21821 9095 21879 9101
rect 21821 9092 21833 9095
rect 21692 9064 21833 9092
rect 21692 9052 21698 9064
rect 21821 9061 21833 9064
rect 21867 9061 21879 9095
rect 21821 9055 21879 9061
rect 21910 9052 21916 9104
rect 21968 9092 21974 9104
rect 23385 9095 23443 9101
rect 23385 9092 23397 9095
rect 21968 9064 23397 9092
rect 21968 9052 21974 9064
rect 23385 9061 23397 9064
rect 23431 9092 23443 9095
rect 23431 9064 24348 9092
rect 23431 9061 23443 9064
rect 23385 9055 23443 9061
rect 23842 9024 23848 9036
rect 18708 8996 19564 9024
rect 21468 8996 22094 9024
rect 14645 8987 14703 8993
rect 9214 8956 9220 8968
rect 4396 8930 8064 8956
rect 4396 8928 6316 8930
rect 6472 8928 8064 8930
rect 8128 8928 9220 8956
rect 4396 8916 4402 8928
rect 5813 8891 5871 8897
rect 5813 8857 5825 8891
rect 5859 8888 5871 8891
rect 5902 8888 5908 8900
rect 5859 8860 5908 8888
rect 5859 8857 5871 8860
rect 5813 8851 5871 8857
rect 5902 8848 5908 8860
rect 5960 8848 5966 8900
rect 8128 8888 8156 8928
rect 9214 8916 9220 8928
rect 9272 8916 9278 8968
rect 10502 8956 10508 8968
rect 10463 8928 10508 8956
rect 10502 8916 10508 8928
rect 10560 8916 10566 8968
rect 10689 8959 10747 8965
rect 10689 8925 10701 8959
rect 10735 8956 10747 8959
rect 11054 8956 11060 8968
rect 10735 8928 11060 8956
rect 10735 8925 10747 8928
rect 10689 8919 10747 8925
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 11149 8959 11207 8965
rect 11149 8925 11161 8959
rect 11195 8956 11207 8959
rect 11698 8956 11704 8968
rect 11195 8928 11704 8956
rect 11195 8925 11207 8928
rect 11149 8919 11207 8925
rect 11698 8916 11704 8928
rect 11756 8916 11762 8968
rect 11882 8916 11888 8968
rect 11940 8956 11946 8968
rect 12894 8956 12900 8968
rect 11940 8928 12900 8956
rect 11940 8916 11946 8928
rect 12894 8916 12900 8928
rect 12952 8916 12958 8968
rect 13170 8956 13176 8968
rect 13131 8928 13176 8956
rect 13170 8916 13176 8928
rect 13228 8916 13234 8968
rect 14660 8956 14688 8987
rect 16942 8965 16948 8968
rect 16669 8959 16727 8965
rect 16669 8956 16681 8959
rect 14660 8928 16681 8956
rect 16669 8925 16681 8928
rect 16715 8925 16727 8959
rect 16936 8956 16948 8965
rect 16903 8928 16948 8956
rect 16669 8919 16727 8925
rect 16936 8919 16948 8928
rect 6564 8860 8156 8888
rect 8205 8891 8263 8897
rect 6564 8820 6592 8860
rect 8205 8857 8217 8891
rect 8251 8888 8263 8891
rect 8386 8888 8392 8900
rect 8251 8860 8392 8888
rect 8251 8857 8263 8860
rect 8205 8851 8263 8857
rect 8386 8848 8392 8860
rect 8444 8848 8450 8900
rect 8478 8848 8484 8900
rect 8536 8888 8542 8900
rect 9401 8891 9459 8897
rect 9401 8888 9413 8891
rect 8536 8860 9413 8888
rect 8536 8848 8542 8860
rect 9401 8857 9413 8860
rect 9447 8857 9459 8891
rect 9401 8851 9459 8857
rect 9582 8848 9588 8900
rect 9640 8888 9646 8900
rect 11416 8891 11474 8897
rect 9640 8860 10824 8888
rect 9640 8848 9646 8860
rect 3896 8792 6592 8820
rect 2685 8783 2743 8789
rect 6638 8780 6644 8832
rect 6696 8820 6702 8832
rect 8294 8820 8300 8832
rect 6696 8792 8300 8820
rect 6696 8780 6702 8792
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 9030 8780 9036 8832
rect 9088 8820 9094 8832
rect 9214 8820 9220 8832
rect 9088 8792 9220 8820
rect 9088 8780 9094 8792
rect 9214 8780 9220 8792
rect 9272 8780 9278 8832
rect 10796 8820 10824 8860
rect 11416 8857 11428 8891
rect 11462 8888 11474 8891
rect 13630 8888 13636 8900
rect 11462 8860 13636 8888
rect 11462 8857 11474 8860
rect 11416 8851 11474 8857
rect 13630 8848 13636 8860
rect 13688 8848 13694 8900
rect 14912 8891 14970 8897
rect 14912 8857 14924 8891
rect 14958 8888 14970 8891
rect 15102 8888 15108 8900
rect 14958 8860 15108 8888
rect 14958 8857 14970 8860
rect 14912 8851 14970 8857
rect 15102 8848 15108 8860
rect 15160 8848 15166 8900
rect 12158 8820 12164 8832
rect 10796 8792 12164 8820
rect 12158 8780 12164 8792
rect 12216 8780 12222 8832
rect 12526 8780 12532 8832
rect 12584 8820 12590 8832
rect 13354 8820 13360 8832
rect 12584 8792 13360 8820
rect 12584 8780 12590 8792
rect 13354 8780 13360 8792
rect 13412 8820 13418 8832
rect 14826 8820 14832 8832
rect 13412 8792 14832 8820
rect 13412 8780 13418 8792
rect 14826 8780 14832 8792
rect 14884 8780 14890 8832
rect 15470 8780 15476 8832
rect 15528 8820 15534 8832
rect 16025 8823 16083 8829
rect 16025 8820 16037 8823
rect 15528 8792 16037 8820
rect 15528 8780 15534 8792
rect 16025 8789 16037 8792
rect 16071 8789 16083 8823
rect 16684 8820 16712 8919
rect 16942 8916 16948 8919
rect 17000 8916 17006 8968
rect 18693 8959 18751 8965
rect 18693 8925 18705 8959
rect 18739 8925 18751 8959
rect 19242 8956 19248 8968
rect 19203 8928 19248 8956
rect 18693 8919 18751 8925
rect 17310 8820 17316 8832
rect 16684 8792 17316 8820
rect 16025 8783 16083 8789
rect 17310 8780 17316 8792
rect 17368 8820 17374 8832
rect 17770 8820 17776 8832
rect 17368 8792 17776 8820
rect 17368 8780 17374 8792
rect 17770 8780 17776 8792
rect 17828 8780 17834 8832
rect 18708 8820 18736 8919
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 19426 8956 19432 8968
rect 19387 8928 19432 8956
rect 19426 8916 19432 8928
rect 19484 8916 19490 8968
rect 19536 8965 19564 8996
rect 19521 8959 19579 8965
rect 19521 8925 19533 8959
rect 19567 8925 19579 8959
rect 19521 8919 19579 8925
rect 19613 8959 19671 8965
rect 19613 8925 19625 8959
rect 19659 8925 19671 8959
rect 19613 8919 19671 8925
rect 19334 8848 19340 8900
rect 19392 8888 19398 8900
rect 19628 8888 19656 8919
rect 19886 8916 19892 8968
rect 19944 8956 19950 8968
rect 20441 8959 20499 8965
rect 20441 8956 20453 8959
rect 19944 8928 20453 8956
rect 19944 8916 19950 8928
rect 20441 8925 20453 8928
rect 20487 8925 20499 8959
rect 20441 8919 20499 8925
rect 20708 8959 20766 8965
rect 20708 8925 20720 8959
rect 20754 8956 20766 8959
rect 21082 8956 21088 8968
rect 20754 8928 21088 8956
rect 20754 8925 20766 8928
rect 20708 8919 20766 8925
rect 21082 8916 21088 8928
rect 21140 8916 21146 8968
rect 19392 8860 19656 8888
rect 19392 8848 19398 8860
rect 20070 8848 20076 8900
rect 20128 8888 20134 8900
rect 21542 8888 21548 8900
rect 20128 8860 21548 8888
rect 20128 8848 20134 8860
rect 21542 8848 21548 8860
rect 21600 8848 21606 8900
rect 22066 8888 22094 8996
rect 23032 8996 23520 9024
rect 22370 8916 22376 8968
rect 22428 8956 22434 8968
rect 23032 8965 23060 8996
rect 22465 8959 22523 8965
rect 22465 8956 22477 8959
rect 22428 8928 22477 8956
rect 22428 8916 22434 8928
rect 22465 8925 22477 8928
rect 22511 8925 22523 8959
rect 22465 8919 22523 8925
rect 23017 8959 23075 8965
rect 23017 8925 23029 8959
rect 23063 8925 23075 8959
rect 23198 8956 23204 8968
rect 23159 8928 23204 8956
rect 23017 8919 23075 8925
rect 23198 8916 23204 8928
rect 23256 8916 23262 8968
rect 23382 8888 23388 8900
rect 22066 8860 23388 8888
rect 23382 8848 23388 8860
rect 23440 8848 23446 8900
rect 23492 8888 23520 8996
rect 23584 8996 23848 9024
rect 23584 8965 23612 8996
rect 23842 8984 23848 8996
rect 23900 8984 23906 9036
rect 23569 8959 23627 8965
rect 23569 8925 23581 8959
rect 23615 8925 23627 8959
rect 23569 8919 23627 8925
rect 23753 8959 23811 8965
rect 23753 8925 23765 8959
rect 23799 8956 23811 8959
rect 24210 8956 24216 8968
rect 23799 8928 24216 8956
rect 23799 8925 23811 8928
rect 23753 8919 23811 8925
rect 24210 8916 24216 8928
rect 24268 8916 24274 8968
rect 24320 8956 24348 9064
rect 24762 8984 24768 9036
rect 24820 9024 24826 9036
rect 24857 9027 24915 9033
rect 24857 9024 24869 9027
rect 24820 8996 24869 9024
rect 24820 8984 24826 8996
rect 24857 8993 24869 8996
rect 24903 8993 24915 9027
rect 27338 9024 27344 9036
rect 24857 8987 24915 8993
rect 26896 8996 27344 9024
rect 25124 8959 25182 8965
rect 24320 8928 24992 8956
rect 24854 8888 24860 8900
rect 23492 8860 24860 8888
rect 24854 8848 24860 8860
rect 24912 8848 24918 8900
rect 24964 8888 24992 8928
rect 25124 8925 25136 8959
rect 25170 8952 25182 8959
rect 25498 8956 25504 8968
rect 25240 8952 25504 8956
rect 25170 8928 25504 8952
rect 25170 8925 25268 8928
rect 25124 8924 25268 8925
rect 25124 8919 25182 8924
rect 25498 8916 25504 8928
rect 25556 8916 25562 8968
rect 26694 8916 26700 8968
rect 26752 8956 26758 8968
rect 26896 8965 26924 8996
rect 27338 8984 27344 8996
rect 27396 8984 27402 9036
rect 26881 8959 26939 8965
rect 26881 8956 26893 8959
rect 26752 8928 26893 8956
rect 26752 8916 26758 8928
rect 26881 8925 26893 8928
rect 26927 8925 26939 8959
rect 27154 8956 27160 8968
rect 27115 8928 27160 8956
rect 26881 8919 26939 8925
rect 27154 8916 27160 8928
rect 27212 8916 27218 8968
rect 26602 8888 26608 8900
rect 24964 8860 26608 8888
rect 26602 8848 26608 8860
rect 26660 8848 26666 8900
rect 20898 8820 20904 8832
rect 18708 8792 20904 8820
rect 20898 8780 20904 8792
rect 20956 8780 20962 8832
rect 20990 8780 20996 8832
rect 21048 8820 21054 8832
rect 21910 8820 21916 8832
rect 21048 8792 21916 8820
rect 21048 8780 21054 8792
rect 21910 8780 21916 8792
rect 21968 8780 21974 8832
rect 22281 8823 22339 8829
rect 22281 8789 22293 8823
rect 22327 8820 22339 8823
rect 23934 8820 23940 8832
rect 22327 8792 23940 8820
rect 22327 8789 22339 8792
rect 22281 8783 22339 8789
rect 23934 8780 23940 8792
rect 23992 8780 23998 8832
rect 26237 8823 26295 8829
rect 26237 8789 26249 8823
rect 26283 8820 26295 8823
rect 26418 8820 26424 8832
rect 26283 8792 26424 8820
rect 26283 8789 26295 8792
rect 26237 8783 26295 8789
rect 26418 8780 26424 8792
rect 26476 8780 26482 8832
rect 26878 8780 26884 8832
rect 26936 8820 26942 8832
rect 27065 8823 27123 8829
rect 27065 8820 27077 8823
rect 26936 8792 27077 8820
rect 26936 8780 26942 8792
rect 27065 8789 27077 8792
rect 27111 8789 27123 8823
rect 27065 8783 27123 8789
rect 1104 8730 28060 8752
rect 1104 8678 9935 8730
rect 9987 8678 9999 8730
rect 10051 8678 10063 8730
rect 10115 8678 10127 8730
rect 10179 8678 10191 8730
rect 10243 8678 18920 8730
rect 18972 8678 18984 8730
rect 19036 8678 19048 8730
rect 19100 8678 19112 8730
rect 19164 8678 19176 8730
rect 19228 8678 28060 8730
rect 1104 8656 28060 8678
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 2961 8619 3019 8625
rect 2961 8616 2973 8619
rect 2924 8588 2973 8616
rect 2924 8576 2930 8588
rect 2961 8585 2973 8588
rect 3007 8585 3019 8619
rect 6546 8616 6552 8628
rect 2961 8579 3019 8585
rect 4448 8588 6552 8616
rect 2590 8548 2596 8560
rect 2551 8520 2596 8548
rect 2590 8508 2596 8520
rect 2648 8508 2654 8560
rect 2777 8551 2835 8557
rect 2777 8517 2789 8551
rect 2823 8548 2835 8551
rect 4448 8548 4476 8588
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 6638 8576 6644 8628
rect 6696 8616 6702 8628
rect 8297 8619 8355 8625
rect 8297 8616 8309 8619
rect 6696 8588 8309 8616
rect 6696 8576 6702 8588
rect 8297 8585 8309 8588
rect 8343 8585 8355 8619
rect 8297 8579 8355 8585
rect 10502 8576 10508 8628
rect 10560 8616 10566 8628
rect 12069 8619 12127 8625
rect 12069 8616 12081 8619
rect 10560 8588 12081 8616
rect 10560 8576 10566 8588
rect 12069 8585 12081 8588
rect 12115 8585 12127 8619
rect 13170 8616 13176 8628
rect 13131 8588 13176 8616
rect 12069 8579 12127 8585
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 13630 8616 13636 8628
rect 13591 8588 13636 8616
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 15930 8616 15936 8628
rect 15488 8588 15936 8616
rect 4614 8548 4620 8560
rect 2823 8520 4476 8548
rect 4575 8520 4620 8548
rect 2823 8517 2835 8520
rect 2777 8511 2835 8517
rect 4614 8508 4620 8520
rect 4672 8508 4678 8560
rect 8849 8551 8907 8557
rect 8849 8517 8861 8551
rect 8895 8548 8907 8551
rect 9490 8548 9496 8560
rect 8895 8520 9496 8548
rect 8895 8517 8907 8520
rect 8849 8511 8907 8517
rect 9490 8508 9496 8520
rect 9548 8508 9554 8560
rect 11606 8508 11612 8560
rect 11664 8548 11670 8560
rect 11701 8551 11759 8557
rect 11701 8548 11713 8551
rect 11664 8520 11713 8548
rect 11664 8508 11670 8520
rect 11701 8517 11713 8520
rect 11747 8517 11759 8551
rect 11701 8511 11759 8517
rect 12710 8508 12716 8560
rect 12768 8548 12774 8560
rect 12805 8551 12863 8557
rect 12805 8548 12817 8551
rect 12768 8520 12817 8548
rect 12768 8508 12774 8520
rect 12805 8517 12817 8520
rect 12851 8517 12863 8551
rect 12805 8511 12863 8517
rect 12897 8551 12955 8557
rect 12897 8517 12909 8551
rect 12943 8548 12955 8551
rect 15194 8548 15200 8560
rect 12943 8520 15200 8548
rect 12943 8517 12955 8520
rect 12897 8511 12955 8517
rect 15194 8508 15200 8520
rect 15252 8508 15258 8560
rect 2038 8480 2044 8492
rect 1999 8452 2044 8480
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8480 3663 8483
rect 3970 8480 3976 8492
rect 3651 8452 3976 8480
rect 3651 8449 3663 8452
rect 3605 8443 3663 8449
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 5258 8480 5264 8492
rect 5219 8452 5264 8480
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 5537 8483 5595 8489
rect 5537 8449 5549 8483
rect 5583 8480 5595 8483
rect 6638 8480 6644 8492
rect 5583 8452 6644 8480
rect 5583 8449 5595 8452
rect 5537 8443 5595 8449
rect 6638 8440 6644 8452
rect 6696 8440 6702 8492
rect 7184 8483 7242 8489
rect 7184 8449 7196 8483
rect 7230 8480 7242 8483
rect 8386 8480 8392 8492
rect 7230 8452 8392 8480
rect 7230 8449 7242 8452
rect 7184 8443 7242 8449
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 8662 8440 8668 8492
rect 8720 8480 8726 8492
rect 8757 8483 8815 8489
rect 8757 8480 8769 8483
rect 8720 8452 8769 8480
rect 8720 8440 8726 8452
rect 8757 8449 8769 8452
rect 8803 8480 8815 8483
rect 9030 8480 9036 8492
rect 8803 8452 9036 8480
rect 8803 8449 8815 8452
rect 8757 8443 8815 8449
rect 9030 8440 9036 8452
rect 9088 8440 9094 8492
rect 11054 8480 11060 8492
rect 9692 8452 11060 8480
rect 5350 8412 5356 8424
rect 5311 8384 5356 8412
rect 5350 8372 5356 8384
rect 5408 8372 5414 8424
rect 6914 8412 6920 8424
rect 6875 8384 6920 8412
rect 6914 8372 6920 8384
rect 6972 8372 6978 8424
rect 9490 8372 9496 8424
rect 9548 8412 9554 8424
rect 9692 8421 9720 8452
rect 11054 8440 11060 8452
rect 11112 8440 11118 8492
rect 11146 8440 11152 8492
rect 11204 8480 11210 8492
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 11204 8452 11529 8480
rect 11204 8440 11210 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11790 8480 11796 8492
rect 11751 8452 11796 8480
rect 11517 8443 11575 8449
rect 11790 8440 11796 8452
rect 11848 8440 11854 8492
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8449 11943 8483
rect 11885 8443 11943 8449
rect 9677 8415 9735 8421
rect 9677 8412 9689 8415
rect 9548 8384 9689 8412
rect 9548 8372 9554 8384
rect 9677 8381 9689 8384
rect 9723 8381 9735 8415
rect 9677 8375 9735 8381
rect 9858 8372 9864 8424
rect 9916 8412 9922 8424
rect 10137 8415 10195 8421
rect 10137 8412 10149 8415
rect 9916 8384 10149 8412
rect 9916 8372 9922 8384
rect 10137 8381 10149 8384
rect 10183 8381 10195 8415
rect 10137 8375 10195 8381
rect 10413 8415 10471 8421
rect 10413 8381 10425 8415
rect 10459 8412 10471 8415
rect 11891 8412 11919 8443
rect 12526 8440 12532 8492
rect 12584 8480 12590 8492
rect 12621 8483 12679 8489
rect 12621 8480 12633 8483
rect 12584 8452 12633 8480
rect 12584 8440 12590 8452
rect 12621 8449 12633 8452
rect 12667 8449 12679 8483
rect 12621 8443 12679 8449
rect 12989 8483 13047 8489
rect 12989 8449 13001 8483
rect 13035 8478 13047 8483
rect 13170 8480 13176 8492
rect 13096 8478 13176 8480
rect 13035 8452 13176 8478
rect 13035 8450 13124 8452
rect 13035 8449 13047 8450
rect 12989 8443 13047 8449
rect 13170 8440 13176 8452
rect 13228 8440 13234 8492
rect 13446 8440 13452 8492
rect 13504 8480 13510 8492
rect 13630 8480 13636 8492
rect 13504 8452 13636 8480
rect 13504 8440 13510 8452
rect 13630 8440 13636 8452
rect 13688 8440 13694 8492
rect 13817 8483 13875 8489
rect 13817 8449 13829 8483
rect 13863 8480 13875 8483
rect 13906 8480 13912 8492
rect 13863 8452 13912 8480
rect 13863 8449 13875 8452
rect 13817 8443 13875 8449
rect 13906 8440 13912 8452
rect 13964 8440 13970 8492
rect 14461 8483 14519 8489
rect 14461 8449 14473 8483
rect 14507 8480 14519 8483
rect 14826 8480 14832 8492
rect 14507 8452 14832 8480
rect 14507 8449 14519 8452
rect 14461 8443 14519 8449
rect 14826 8440 14832 8452
rect 14884 8440 14890 8492
rect 15381 8483 15439 8489
rect 15381 8449 15393 8483
rect 15427 8480 15439 8483
rect 15488 8480 15516 8588
rect 15930 8576 15936 8588
rect 15988 8576 15994 8628
rect 17034 8616 17040 8628
rect 16995 8588 17040 8616
rect 17034 8576 17040 8588
rect 17092 8576 17098 8628
rect 18414 8616 18420 8628
rect 17604 8588 18420 8616
rect 15657 8551 15715 8557
rect 15657 8517 15669 8551
rect 15703 8548 15715 8551
rect 15838 8548 15844 8560
rect 15703 8520 15844 8548
rect 15703 8517 15715 8520
rect 15657 8511 15715 8517
rect 15838 8508 15844 8520
rect 15896 8508 15902 8560
rect 17604 8557 17632 8588
rect 18414 8576 18420 8588
rect 18472 8576 18478 8628
rect 18877 8619 18935 8625
rect 18877 8585 18889 8619
rect 18923 8616 18935 8619
rect 19518 8616 19524 8628
rect 18923 8588 19524 8616
rect 18923 8585 18935 8588
rect 18877 8579 18935 8585
rect 19518 8576 19524 8588
rect 19576 8576 19582 8628
rect 19889 8619 19947 8625
rect 19628 8588 19840 8616
rect 17589 8551 17647 8557
rect 16776 8520 16988 8548
rect 16776 8489 16804 8520
rect 15427 8452 15516 8480
rect 15565 8483 15623 8489
rect 15427 8449 15439 8452
rect 15381 8443 15439 8449
rect 15565 8449 15577 8483
rect 15611 8449 15623 8483
rect 15565 8443 15623 8449
rect 15749 8483 15807 8489
rect 15749 8449 15761 8483
rect 15795 8449 15807 8483
rect 15749 8443 15807 8449
rect 16761 8483 16819 8489
rect 16761 8449 16773 8483
rect 16807 8449 16819 8483
rect 16761 8443 16819 8449
rect 16853 8483 16911 8489
rect 16853 8449 16865 8483
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 12342 8412 12348 8424
rect 10459 8384 12348 8412
rect 10459 8381 10471 8384
rect 10413 8375 10471 8381
rect 12342 8372 12348 8384
rect 12400 8372 12406 8424
rect 14277 8415 14335 8421
rect 14277 8381 14289 8415
rect 14323 8381 14335 8415
rect 14277 8375 14335 8381
rect 2130 8304 2136 8356
rect 2188 8344 2194 8356
rect 3421 8347 3479 8353
rect 3421 8344 3433 8347
rect 2188 8316 3433 8344
rect 2188 8304 2194 8316
rect 3421 8313 3433 8316
rect 3467 8313 3479 8347
rect 3421 8307 3479 8313
rect 5721 8347 5779 8353
rect 5721 8313 5733 8347
rect 5767 8344 5779 8347
rect 6730 8344 6736 8356
rect 5767 8316 6736 8344
rect 5767 8313 5779 8316
rect 5721 8307 5779 8313
rect 6730 8304 6736 8316
rect 6788 8304 6794 8356
rect 8294 8304 8300 8356
rect 8352 8344 8358 8356
rect 12526 8344 12532 8356
rect 8352 8316 12532 8344
rect 8352 8304 8358 8316
rect 12526 8304 12532 8316
rect 12584 8304 12590 8356
rect 12710 8304 12716 8356
rect 12768 8344 12774 8356
rect 14292 8344 14320 8375
rect 15580 8356 15608 8443
rect 15764 8412 15792 8443
rect 15838 8412 15844 8424
rect 15764 8384 15844 8412
rect 15838 8372 15844 8384
rect 15896 8412 15902 8424
rect 16206 8412 16212 8424
rect 15896 8384 16212 8412
rect 15896 8372 15902 8384
rect 16206 8372 16212 8384
rect 16264 8372 16270 8424
rect 14645 8347 14703 8353
rect 12768 8316 12848 8344
rect 14292 8316 14504 8344
rect 12768 8304 12774 8316
rect 1854 8276 1860 8288
rect 1815 8248 1860 8276
rect 1854 8236 1860 8248
rect 1912 8236 1918 8288
rect 4062 8236 4068 8288
rect 4120 8276 4126 8288
rect 4246 8276 4252 8288
rect 4120 8248 4252 8276
rect 4120 8236 4126 8248
rect 4246 8236 4252 8248
rect 4304 8236 4310 8288
rect 4614 8236 4620 8288
rect 4672 8276 4678 8288
rect 4709 8279 4767 8285
rect 4709 8276 4721 8279
rect 4672 8248 4721 8276
rect 4672 8236 4678 8248
rect 4709 8245 4721 8248
rect 4755 8245 4767 8279
rect 5350 8276 5356 8288
rect 5311 8248 5356 8276
rect 4709 8239 4767 8245
rect 5350 8236 5356 8248
rect 5408 8236 5414 8288
rect 6822 8236 6828 8288
rect 6880 8276 6886 8288
rect 8662 8276 8668 8288
rect 6880 8248 8668 8276
rect 6880 8236 6886 8248
rect 8662 8236 8668 8248
rect 8720 8236 8726 8288
rect 11698 8236 11704 8288
rect 11756 8276 11762 8288
rect 12820 8276 12848 8316
rect 13354 8276 13360 8288
rect 11756 8248 13360 8276
rect 11756 8236 11762 8248
rect 13354 8236 13360 8248
rect 13412 8236 13418 8288
rect 13906 8236 13912 8288
rect 13964 8276 13970 8288
rect 14476 8276 14504 8316
rect 14645 8313 14657 8347
rect 14691 8344 14703 8347
rect 15286 8344 15292 8356
rect 14691 8316 15292 8344
rect 14691 8313 14703 8316
rect 14645 8307 14703 8313
rect 15286 8304 15292 8316
rect 15344 8304 15350 8356
rect 15562 8304 15568 8356
rect 15620 8304 15626 8356
rect 15933 8347 15991 8353
rect 15933 8313 15945 8347
rect 15979 8344 15991 8347
rect 16868 8344 16896 8443
rect 16960 8424 16988 8520
rect 17589 8517 17601 8551
rect 17635 8517 17647 8551
rect 17770 8548 17776 8560
rect 17731 8520 17776 8548
rect 17589 8511 17647 8517
rect 17770 8508 17776 8520
rect 17828 8508 17834 8560
rect 19628 8548 19656 8588
rect 18432 8520 19656 8548
rect 19812 8548 19840 8588
rect 19889 8585 19901 8619
rect 19935 8616 19947 8619
rect 19978 8616 19984 8628
rect 19935 8588 19984 8616
rect 19935 8585 19947 8588
rect 19889 8579 19947 8585
rect 19978 8576 19984 8588
rect 20036 8576 20042 8628
rect 20254 8576 20260 8628
rect 20312 8616 20318 8628
rect 21634 8616 21640 8628
rect 20312 8588 21640 8616
rect 20312 8576 20318 8588
rect 21634 8576 21640 8588
rect 21692 8576 21698 8628
rect 23658 8616 23664 8628
rect 22066 8588 23664 8616
rect 22066 8548 22094 8588
rect 23658 8576 23664 8588
rect 23716 8576 23722 8628
rect 23753 8619 23811 8625
rect 23753 8585 23765 8619
rect 23799 8616 23811 8619
rect 25130 8616 25136 8628
rect 23799 8588 25136 8616
rect 23799 8585 23811 8588
rect 23753 8579 23811 8585
rect 25130 8576 25136 8588
rect 25188 8576 25194 8628
rect 25314 8576 25320 8628
rect 25372 8616 25378 8628
rect 27338 8616 27344 8628
rect 25372 8588 27344 8616
rect 25372 8576 25378 8588
rect 27338 8576 27344 8588
rect 27396 8576 27402 8628
rect 19812 8520 22094 8548
rect 22373 8551 22431 8557
rect 18432 8489 18460 8520
rect 22373 8517 22385 8551
rect 22419 8548 22431 8551
rect 22738 8548 22744 8560
rect 22419 8520 22744 8548
rect 22419 8517 22431 8520
rect 22373 8511 22431 8517
rect 22738 8508 22744 8520
rect 22796 8508 22802 8560
rect 23106 8548 23112 8560
rect 23067 8520 23112 8548
rect 23106 8508 23112 8520
rect 23164 8508 23170 8560
rect 25774 8548 25780 8560
rect 23860 8520 25780 8548
rect 18417 8483 18475 8489
rect 18417 8449 18429 8483
rect 18463 8449 18475 8483
rect 18417 8443 18475 8449
rect 19061 8483 19119 8489
rect 19061 8449 19073 8483
rect 19107 8480 19119 8483
rect 19107 8452 19656 8480
rect 19107 8449 19119 8452
rect 19061 8443 19119 8449
rect 16942 8372 16948 8424
rect 17000 8412 17006 8424
rect 19426 8412 19432 8424
rect 17000 8384 19432 8412
rect 17000 8372 17006 8384
rect 19426 8372 19432 8384
rect 19484 8412 19490 8424
rect 19521 8415 19579 8421
rect 19521 8412 19533 8415
rect 19484 8384 19533 8412
rect 19484 8372 19490 8384
rect 19521 8381 19533 8384
rect 19567 8381 19579 8415
rect 19628 8412 19656 8452
rect 19702 8440 19708 8492
rect 19760 8480 19766 8492
rect 20806 8480 20812 8492
rect 19760 8452 19805 8480
rect 20767 8452 20812 8480
rect 19760 8440 19766 8452
rect 20806 8440 20812 8452
rect 20864 8440 20870 8492
rect 20898 8440 20904 8492
rect 20956 8480 20962 8492
rect 23860 8480 23888 8520
rect 25774 8508 25780 8520
rect 25832 8508 25838 8560
rect 26050 8508 26056 8560
rect 26108 8548 26114 8560
rect 27246 8548 27252 8560
rect 26108 8520 27252 8548
rect 26108 8508 26114 8520
rect 27246 8508 27252 8520
rect 27304 8508 27310 8560
rect 20956 8452 23888 8480
rect 23937 8483 23995 8489
rect 20956 8440 20962 8452
rect 23937 8449 23949 8483
rect 23983 8480 23995 8483
rect 24118 8480 24124 8492
rect 23983 8452 24124 8480
rect 23983 8449 23995 8452
rect 23937 8443 23995 8449
rect 24118 8440 24124 8452
rect 24176 8440 24182 8492
rect 24210 8440 24216 8492
rect 24268 8480 24274 8492
rect 24581 8483 24639 8489
rect 24581 8480 24593 8483
rect 24268 8452 24593 8480
rect 24268 8440 24274 8452
rect 24581 8449 24593 8452
rect 24627 8449 24639 8483
rect 24581 8443 24639 8449
rect 25308 8483 25366 8489
rect 25308 8449 25320 8483
rect 25354 8480 25366 8483
rect 26142 8480 26148 8492
rect 25354 8452 26148 8480
rect 25354 8449 25366 8452
rect 25308 8443 25366 8449
rect 26142 8440 26148 8452
rect 26200 8440 26206 8492
rect 26786 8440 26792 8492
rect 26844 8480 26850 8492
rect 26973 8483 27031 8489
rect 26973 8480 26985 8483
rect 26844 8452 26985 8480
rect 26844 8440 26850 8452
rect 26973 8449 26985 8452
rect 27019 8449 27031 8483
rect 26973 8443 27031 8449
rect 19628 8384 23152 8412
rect 19521 8375 19579 8381
rect 15979 8316 16896 8344
rect 18233 8347 18291 8353
rect 15979 8313 15991 8316
rect 15933 8307 15991 8313
rect 18233 8313 18245 8347
rect 18279 8344 18291 8347
rect 20070 8344 20076 8356
rect 18279 8316 20076 8344
rect 18279 8313 18291 8316
rect 18233 8307 18291 8313
rect 20070 8304 20076 8316
rect 20128 8304 20134 8356
rect 20625 8347 20683 8353
rect 20625 8313 20637 8347
rect 20671 8344 20683 8347
rect 21082 8344 21088 8356
rect 20671 8316 21088 8344
rect 20671 8313 20683 8316
rect 20625 8307 20683 8313
rect 21082 8304 21088 8316
rect 21140 8304 21146 8356
rect 22557 8347 22615 8353
rect 22557 8313 22569 8347
rect 22603 8344 22615 8347
rect 22738 8344 22744 8356
rect 22603 8316 22744 8344
rect 22603 8313 22615 8316
rect 22557 8307 22615 8313
rect 22738 8304 22744 8316
rect 22796 8304 22802 8356
rect 23124 8344 23152 8384
rect 23198 8372 23204 8424
rect 23256 8412 23262 8424
rect 25041 8415 25099 8421
rect 25041 8412 25053 8415
rect 23256 8384 25053 8412
rect 23256 8372 23262 8384
rect 25041 8381 25053 8384
rect 25087 8381 25099 8415
rect 27246 8412 27252 8424
rect 25041 8375 25099 8381
rect 26252 8384 27252 8412
rect 26252 8344 26280 8384
rect 27246 8372 27252 8384
rect 27304 8372 27310 8424
rect 23124 8316 25084 8344
rect 16850 8276 16856 8288
rect 13964 8248 16856 8276
rect 13964 8236 13970 8248
rect 16850 8236 16856 8248
rect 16908 8236 16914 8288
rect 23198 8276 23204 8288
rect 23159 8248 23204 8276
rect 23198 8236 23204 8248
rect 23256 8236 23262 8288
rect 24394 8276 24400 8288
rect 24355 8248 24400 8276
rect 24394 8236 24400 8248
rect 24452 8236 24458 8288
rect 25056 8276 25084 8316
rect 25976 8316 26280 8344
rect 25976 8276 26004 8316
rect 26510 8304 26516 8356
rect 26568 8344 26574 8356
rect 27157 8347 27215 8353
rect 27157 8344 27169 8347
rect 26568 8316 27169 8344
rect 26568 8304 26574 8316
rect 27157 8313 27169 8316
rect 27203 8313 27215 8347
rect 27157 8307 27215 8313
rect 25056 8248 26004 8276
rect 26421 8279 26479 8285
rect 26421 8245 26433 8279
rect 26467 8276 26479 8279
rect 26970 8276 26976 8288
rect 26467 8248 26976 8276
rect 26467 8245 26479 8248
rect 26421 8239 26479 8245
rect 26970 8236 26976 8248
rect 27028 8236 27034 8288
rect 1104 8186 28060 8208
rect 1104 8134 5442 8186
rect 5494 8134 5506 8186
rect 5558 8134 5570 8186
rect 5622 8134 5634 8186
rect 5686 8134 5698 8186
rect 5750 8134 14428 8186
rect 14480 8134 14492 8186
rect 14544 8134 14556 8186
rect 14608 8134 14620 8186
rect 14672 8134 14684 8186
rect 14736 8134 23413 8186
rect 23465 8134 23477 8186
rect 23529 8134 23541 8186
rect 23593 8134 23605 8186
rect 23657 8134 23669 8186
rect 23721 8134 28060 8186
rect 1104 8112 28060 8134
rect 3234 8032 3240 8084
rect 3292 8072 3298 8084
rect 3970 8072 3976 8084
rect 3292 8044 3976 8072
rect 3292 8032 3298 8044
rect 3970 8032 3976 8044
rect 4028 8032 4034 8084
rect 4062 8032 4068 8084
rect 4120 8072 4126 8084
rect 5629 8075 5687 8081
rect 5629 8072 5641 8075
rect 4120 8044 5641 8072
rect 4120 8032 4126 8044
rect 5629 8041 5641 8044
rect 5675 8041 5687 8075
rect 5629 8035 5687 8041
rect 6730 8032 6736 8084
rect 6788 8072 6794 8084
rect 7926 8072 7932 8084
rect 6788 8044 7932 8072
rect 6788 8032 6794 8044
rect 7926 8032 7932 8044
rect 7984 8032 7990 8084
rect 8202 8032 8208 8084
rect 8260 8072 8266 8084
rect 9309 8075 9367 8081
rect 9309 8072 9321 8075
rect 8260 8044 9321 8072
rect 8260 8032 8266 8044
rect 9309 8041 9321 8044
rect 9355 8041 9367 8075
rect 9309 8035 9367 8041
rect 13262 8032 13268 8084
rect 13320 8072 13326 8084
rect 13446 8072 13452 8084
rect 13320 8044 13452 8072
rect 13320 8032 13326 8044
rect 13446 8032 13452 8044
rect 13504 8032 13510 8084
rect 15102 8072 15108 8084
rect 15063 8044 15108 8072
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 18693 8075 18751 8081
rect 18693 8072 18705 8075
rect 15856 8044 18705 8072
rect 2774 7964 2780 8016
rect 2832 8004 2838 8016
rect 3418 8004 3424 8016
rect 2832 7976 3424 8004
rect 2832 7964 2838 7976
rect 3418 7964 3424 7976
rect 3476 7964 3482 8016
rect 5258 7964 5264 8016
rect 5316 8004 5322 8016
rect 6089 8007 6147 8013
rect 6089 8004 6101 8007
rect 5316 7976 6101 8004
rect 5316 7964 5322 7976
rect 6089 7973 6101 7976
rect 6135 7973 6147 8007
rect 6089 7967 6147 7973
rect 7374 7964 7380 8016
rect 7432 8004 7438 8016
rect 7432 7976 8156 8004
rect 7432 7964 7438 7976
rect 5810 7936 5816 7948
rect 5771 7908 5816 7936
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 6454 7896 6460 7948
rect 6512 7936 6518 7948
rect 7653 7939 7711 7945
rect 7653 7936 7665 7939
rect 6512 7908 7665 7936
rect 6512 7896 6518 7908
rect 7653 7905 7665 7908
rect 7699 7905 7711 7939
rect 7653 7899 7711 7905
rect 8128 7880 8156 7976
rect 8938 7964 8944 8016
rect 8996 8004 9002 8016
rect 11882 8004 11888 8016
rect 8996 7976 11888 8004
rect 8996 7964 9002 7976
rect 11882 7964 11888 7976
rect 11940 7964 11946 8016
rect 12066 8004 12072 8016
rect 12027 7976 12072 8004
rect 12066 7964 12072 7976
rect 12124 7964 12130 8016
rect 13538 8004 13544 8016
rect 12820 7976 13544 8004
rect 10597 7939 10655 7945
rect 10597 7905 10609 7939
rect 10643 7936 10655 7939
rect 11698 7936 11704 7948
rect 10643 7908 11704 7936
rect 10643 7905 10655 7908
rect 10597 7899 10655 7905
rect 11698 7896 11704 7908
rect 11756 7896 11762 7948
rect 1578 7868 1584 7880
rect 1539 7840 1584 7868
rect 1578 7828 1584 7840
rect 1636 7868 1642 7880
rect 3786 7868 3792 7880
rect 1636 7840 3792 7868
rect 1636 7828 1642 7840
rect 3786 7828 3792 7840
rect 3844 7868 3850 7880
rect 4614 7868 4620 7880
rect 3844 7840 4620 7868
rect 3844 7828 3850 7840
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 5905 7871 5963 7877
rect 5905 7837 5917 7871
rect 5951 7837 5963 7871
rect 6638 7868 6644 7880
rect 6599 7840 6644 7868
rect 5905 7831 5963 7837
rect 1854 7809 1860 7812
rect 1848 7800 1860 7809
rect 1815 7772 1860 7800
rect 1848 7763 1860 7772
rect 1854 7760 1860 7763
rect 1912 7760 1918 7812
rect 3418 7760 3424 7812
rect 3476 7800 3482 7812
rect 4034 7803 4092 7809
rect 4034 7800 4046 7803
rect 3476 7772 4046 7800
rect 3476 7760 3482 7772
rect 4034 7769 4046 7772
rect 4080 7769 4092 7803
rect 5629 7803 5687 7809
rect 5629 7800 5641 7803
rect 4034 7763 4092 7769
rect 4172 7772 5641 7800
rect 2961 7735 3019 7741
rect 2961 7701 2973 7735
rect 3007 7732 3019 7735
rect 3234 7732 3240 7744
rect 3007 7704 3240 7732
rect 3007 7701 3019 7704
rect 2961 7695 3019 7701
rect 3234 7692 3240 7704
rect 3292 7732 3298 7744
rect 4172 7732 4200 7772
rect 5629 7769 5641 7772
rect 5675 7769 5687 7803
rect 5629 7763 5687 7769
rect 3292 7704 4200 7732
rect 5169 7735 5227 7741
rect 3292 7692 3298 7704
rect 5169 7701 5181 7735
rect 5215 7732 5227 7735
rect 5258 7732 5264 7744
rect 5215 7704 5264 7732
rect 5215 7701 5227 7704
rect 5169 7695 5227 7701
rect 5258 7692 5264 7704
rect 5316 7732 5322 7744
rect 5920 7732 5948 7831
rect 6638 7828 6644 7840
rect 6696 7828 6702 7880
rect 6730 7828 6736 7880
rect 6788 7868 6794 7880
rect 6917 7871 6975 7877
rect 6917 7868 6929 7871
rect 6788 7840 6929 7868
rect 6788 7828 6794 7840
rect 6917 7837 6929 7840
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 6362 7760 6368 7812
rect 6420 7800 6426 7812
rect 6825 7803 6883 7809
rect 6825 7800 6837 7803
rect 6420 7772 6837 7800
rect 6420 7760 6426 7772
rect 6825 7769 6837 7772
rect 6871 7769 6883 7803
rect 7024 7800 7052 7831
rect 7852 7800 7880 7831
rect 8110 7828 8116 7880
rect 8168 7828 8174 7880
rect 10042 7828 10048 7880
rect 10100 7868 10106 7880
rect 10321 7871 10379 7877
rect 10321 7868 10333 7871
rect 10100 7840 10333 7868
rect 10100 7828 10106 7840
rect 10321 7837 10333 7840
rect 10367 7868 10379 7871
rect 10502 7868 10508 7880
rect 10367 7840 10508 7868
rect 10367 7837 10379 7840
rect 10321 7831 10379 7837
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 11054 7828 11060 7880
rect 11112 7868 11118 7880
rect 11885 7871 11943 7877
rect 11885 7868 11897 7871
rect 11112 7840 11897 7868
rect 11112 7828 11118 7840
rect 11885 7837 11897 7840
rect 11931 7868 11943 7871
rect 11974 7868 11980 7880
rect 11931 7840 11980 7868
rect 11931 7837 11943 7840
rect 11885 7831 11943 7837
rect 11974 7828 11980 7840
rect 12032 7828 12038 7880
rect 8938 7800 8944 7812
rect 6825 7763 6883 7769
rect 6932 7772 7052 7800
rect 7208 7772 7880 7800
rect 8899 7772 8944 7800
rect 5316 7704 5948 7732
rect 5316 7692 5322 7704
rect 6730 7692 6736 7744
rect 6788 7732 6794 7744
rect 6932 7732 6960 7772
rect 7208 7741 7236 7772
rect 8938 7760 8944 7772
rect 8996 7760 9002 7812
rect 9125 7803 9183 7809
rect 9125 7769 9137 7803
rect 9171 7800 9183 7803
rect 9490 7800 9496 7812
rect 9171 7772 9496 7800
rect 9171 7769 9183 7772
rect 9125 7763 9183 7769
rect 9490 7760 9496 7772
rect 9548 7760 9554 7812
rect 10134 7760 10140 7812
rect 10192 7800 10198 7812
rect 11330 7800 11336 7812
rect 10192 7772 11336 7800
rect 10192 7760 10198 7772
rect 11330 7760 11336 7772
rect 11388 7760 11394 7812
rect 12342 7760 12348 7812
rect 12400 7800 12406 7812
rect 12621 7803 12679 7809
rect 12621 7800 12633 7803
rect 12400 7772 12633 7800
rect 12400 7760 12406 7772
rect 12621 7769 12633 7772
rect 12667 7769 12679 7803
rect 12621 7763 12679 7769
rect 12710 7760 12716 7812
rect 12768 7800 12774 7812
rect 12820 7809 12848 7976
rect 13538 7964 13544 7976
rect 13596 7964 13602 8016
rect 14182 7964 14188 8016
rect 14240 8004 14246 8016
rect 14645 8007 14703 8013
rect 14240 7976 14504 8004
rect 14240 7964 14246 7976
rect 13354 7896 13360 7948
rect 13412 7936 13418 7948
rect 13412 7908 14228 7936
rect 13412 7896 13418 7908
rect 13265 7871 13323 7877
rect 13265 7837 13277 7871
rect 13311 7868 13323 7871
rect 13538 7868 13544 7880
rect 13311 7840 13544 7868
rect 13311 7837 13323 7840
rect 13265 7831 13323 7837
rect 12805 7803 12863 7809
rect 12805 7800 12817 7803
rect 12768 7772 12817 7800
rect 12768 7760 12774 7772
rect 12805 7769 12817 7772
rect 12851 7769 12863 7803
rect 12805 7763 12863 7769
rect 6788 7704 6960 7732
rect 7193 7735 7251 7741
rect 6788 7692 6794 7704
rect 7193 7701 7205 7735
rect 7239 7701 7251 7735
rect 7193 7695 7251 7701
rect 7926 7692 7932 7744
rect 7984 7732 7990 7744
rect 8021 7735 8079 7741
rect 8021 7732 8033 7735
rect 7984 7704 8033 7732
rect 7984 7692 7990 7704
rect 8021 7701 8033 7704
rect 8067 7701 8079 7735
rect 8021 7695 8079 7701
rect 11054 7692 11060 7744
rect 11112 7732 11118 7744
rect 13280 7732 13308 7831
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 14093 7871 14151 7877
rect 14093 7837 14105 7871
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 11112 7704 13308 7732
rect 14108 7732 14136 7831
rect 14200 7800 14228 7908
rect 14366 7868 14372 7880
rect 14327 7840 14372 7868
rect 14366 7828 14372 7840
rect 14424 7828 14430 7880
rect 14476 7877 14504 7976
rect 14645 7973 14657 8007
rect 14691 8004 14703 8007
rect 14826 8004 14832 8016
rect 14691 7976 14832 8004
rect 14691 7973 14703 7976
rect 14645 7967 14703 7973
rect 14826 7964 14832 7976
rect 14884 7964 14890 8016
rect 14461 7871 14519 7877
rect 14461 7837 14473 7871
rect 14507 7837 14519 7871
rect 15286 7868 15292 7880
rect 15247 7840 15292 7868
rect 14461 7831 14519 7837
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 15856 7877 15884 8044
rect 18693 8041 18705 8044
rect 18739 8072 18751 8075
rect 22002 8072 22008 8084
rect 18739 8044 22008 8072
rect 18739 8041 18751 8044
rect 18693 8035 18751 8041
rect 22002 8032 22008 8044
rect 22060 8032 22066 8084
rect 23106 8072 23112 8084
rect 22480 8044 23112 8072
rect 19242 7964 19248 8016
rect 19300 8004 19306 8016
rect 19613 8007 19671 8013
rect 19613 8004 19625 8007
rect 19300 7976 19625 8004
rect 19300 7964 19306 7976
rect 19613 7973 19625 7976
rect 19659 7973 19671 8007
rect 22480 8004 22508 8044
rect 23106 8032 23112 8044
rect 23164 8032 23170 8084
rect 26142 8032 26148 8084
rect 26200 8072 26206 8084
rect 26421 8075 26479 8081
rect 26421 8072 26433 8075
rect 26200 8044 26433 8072
rect 26200 8032 26206 8044
rect 26421 8041 26433 8044
rect 26467 8041 26479 8075
rect 26421 8035 26479 8041
rect 19613 7967 19671 7973
rect 21560 7976 22508 8004
rect 24044 7976 24532 8004
rect 17310 7936 17316 7948
rect 17271 7908 17316 7936
rect 17310 7896 17316 7908
rect 17368 7896 17374 7948
rect 18598 7896 18604 7948
rect 18656 7936 18662 7948
rect 18656 7908 20300 7936
rect 18656 7896 18662 7908
rect 15841 7871 15899 7877
rect 15841 7837 15853 7871
rect 15887 7837 15899 7871
rect 16206 7868 16212 7880
rect 16167 7840 16212 7868
rect 15841 7831 15899 7837
rect 16206 7828 16212 7840
rect 16264 7828 16270 7880
rect 17586 7877 17592 7880
rect 17580 7868 17592 7877
rect 17547 7840 17592 7868
rect 17580 7831 17592 7840
rect 17586 7828 17592 7831
rect 17644 7828 17650 7880
rect 19886 7828 19892 7880
rect 19944 7868 19950 7880
rect 20165 7871 20223 7877
rect 20165 7868 20177 7871
rect 19944 7840 20177 7868
rect 19944 7828 19950 7840
rect 20165 7837 20177 7840
rect 20211 7837 20223 7871
rect 20272 7868 20300 7908
rect 20421 7871 20479 7877
rect 20421 7868 20433 7871
rect 20272 7840 20433 7868
rect 20165 7831 20223 7837
rect 20421 7837 20433 7840
rect 20467 7837 20479 7871
rect 20421 7831 20479 7837
rect 14277 7803 14335 7809
rect 14277 7800 14289 7803
rect 14200 7772 14289 7800
rect 14277 7769 14289 7772
rect 14323 7800 14335 7803
rect 15562 7800 15568 7812
rect 14323 7772 15568 7800
rect 14323 7769 14335 7772
rect 14277 7763 14335 7769
rect 15562 7760 15568 7772
rect 15620 7800 15626 7812
rect 16025 7803 16083 7809
rect 16025 7800 16037 7803
rect 15620 7772 16037 7800
rect 15620 7760 15626 7772
rect 16025 7769 16037 7772
rect 16071 7769 16083 7803
rect 16025 7763 16083 7769
rect 16117 7803 16175 7809
rect 16117 7769 16129 7803
rect 16163 7800 16175 7803
rect 16298 7800 16304 7812
rect 16163 7772 16304 7800
rect 16163 7769 16175 7772
rect 16117 7763 16175 7769
rect 16298 7760 16304 7772
rect 16356 7760 16362 7812
rect 19242 7800 19248 7812
rect 19203 7772 19248 7800
rect 19242 7760 19248 7772
rect 19300 7760 19306 7812
rect 19334 7760 19340 7812
rect 19392 7800 19398 7812
rect 19429 7803 19487 7809
rect 19429 7800 19441 7803
rect 19392 7772 19441 7800
rect 19392 7760 19398 7772
rect 19429 7769 19441 7772
rect 19475 7769 19487 7803
rect 19429 7763 19487 7769
rect 21560 7744 21588 7976
rect 22186 7828 22192 7880
rect 22244 7868 22250 7880
rect 22465 7871 22523 7877
rect 22465 7868 22477 7871
rect 22244 7840 22477 7868
rect 22244 7828 22250 7840
rect 22465 7837 22477 7840
rect 22511 7868 22523 7871
rect 23198 7868 23204 7880
rect 22511 7840 23204 7868
rect 22511 7837 22523 7840
rect 22465 7831 22523 7837
rect 23198 7828 23204 7840
rect 23256 7868 23262 7880
rect 24044 7868 24072 7976
rect 24302 7868 24308 7880
rect 23256 7840 24072 7868
rect 24136 7840 24308 7868
rect 23256 7828 23262 7840
rect 22732 7803 22790 7809
rect 22732 7769 22744 7803
rect 22778 7800 22790 7803
rect 23290 7800 23296 7812
rect 22778 7772 23296 7800
rect 22778 7769 22790 7772
rect 22732 7763 22790 7769
rect 23290 7760 23296 7772
rect 23348 7760 23354 7812
rect 24136 7800 24164 7840
rect 24302 7828 24308 7840
rect 24360 7828 24366 7880
rect 24504 7877 24532 7976
rect 24489 7871 24547 7877
rect 24489 7837 24501 7871
rect 24535 7837 24547 7871
rect 24489 7831 24547 7837
rect 24578 7828 24584 7880
rect 24636 7868 24642 7880
rect 24745 7871 24803 7877
rect 24745 7868 24757 7871
rect 24636 7840 24757 7868
rect 24636 7828 24642 7840
rect 24745 7837 24757 7840
rect 24791 7837 24803 7871
rect 24745 7831 24803 7837
rect 25038 7828 25044 7880
rect 25096 7868 25102 7880
rect 25958 7868 25964 7880
rect 25096 7840 25964 7868
rect 25096 7828 25102 7840
rect 25958 7828 25964 7840
rect 26016 7828 26022 7880
rect 26605 7871 26663 7877
rect 26605 7837 26617 7871
rect 26651 7868 26663 7871
rect 26694 7868 26700 7880
rect 26651 7840 26700 7868
rect 26651 7837 26663 7840
rect 26605 7831 26663 7837
rect 26694 7828 26700 7840
rect 26752 7828 26758 7880
rect 26881 7871 26939 7877
rect 26881 7837 26893 7871
rect 26927 7868 26939 7871
rect 27154 7868 27160 7880
rect 26927 7840 27160 7868
rect 26927 7837 26939 7840
rect 26881 7831 26939 7837
rect 27154 7828 27160 7840
rect 27212 7828 27218 7880
rect 23676 7772 24164 7800
rect 15470 7732 15476 7744
rect 14108 7704 15476 7732
rect 11112 7692 11118 7704
rect 15470 7692 15476 7704
rect 15528 7692 15534 7744
rect 16393 7735 16451 7741
rect 16393 7701 16405 7735
rect 16439 7732 16451 7735
rect 16942 7732 16948 7744
rect 16439 7704 16948 7732
rect 16439 7701 16451 7704
rect 16393 7695 16451 7701
rect 16942 7692 16948 7704
rect 17000 7692 17006 7744
rect 17678 7692 17684 7744
rect 17736 7732 17742 7744
rect 18138 7732 18144 7744
rect 17736 7704 18144 7732
rect 17736 7692 17742 7704
rect 18138 7692 18144 7704
rect 18196 7692 18202 7744
rect 21542 7732 21548 7744
rect 21503 7704 21548 7732
rect 21542 7692 21548 7704
rect 21600 7692 21606 7744
rect 21910 7692 21916 7744
rect 21968 7732 21974 7744
rect 23676 7732 23704 7772
rect 24210 7760 24216 7812
rect 24268 7800 24274 7812
rect 27982 7800 27988 7812
rect 24268 7772 27988 7800
rect 24268 7760 24274 7772
rect 27982 7760 27988 7772
rect 28040 7760 28046 7812
rect 21968 7704 23704 7732
rect 21968 7692 21974 7704
rect 23750 7692 23756 7744
rect 23808 7732 23814 7744
rect 23845 7735 23903 7741
rect 23845 7732 23857 7735
rect 23808 7704 23857 7732
rect 23808 7692 23814 7704
rect 23845 7701 23857 7704
rect 23891 7701 23903 7735
rect 23845 7695 23903 7701
rect 24578 7692 24584 7744
rect 24636 7732 24642 7744
rect 25869 7735 25927 7741
rect 25869 7732 25881 7735
rect 24636 7704 25881 7732
rect 24636 7692 24642 7704
rect 25869 7701 25881 7704
rect 25915 7701 25927 7735
rect 25869 7695 25927 7701
rect 26789 7735 26847 7741
rect 26789 7701 26801 7735
rect 26835 7732 26847 7735
rect 26970 7732 26976 7744
rect 26835 7704 26976 7732
rect 26835 7701 26847 7704
rect 26789 7695 26847 7701
rect 26970 7692 26976 7704
rect 27028 7692 27034 7744
rect 1104 7642 28060 7664
rect 1104 7590 9935 7642
rect 9987 7590 9999 7642
rect 10051 7590 10063 7642
rect 10115 7590 10127 7642
rect 10179 7590 10191 7642
rect 10243 7590 18920 7642
rect 18972 7590 18984 7642
rect 19036 7590 19048 7642
rect 19100 7590 19112 7642
rect 19164 7590 19176 7642
rect 19228 7590 28060 7642
rect 1104 7568 28060 7590
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 2225 7531 2283 7537
rect 2225 7528 2237 7531
rect 2096 7500 2237 7528
rect 2096 7488 2102 7500
rect 2225 7497 2237 7500
rect 2271 7497 2283 7531
rect 2225 7491 2283 7497
rect 2682 7488 2688 7540
rect 2740 7528 2746 7540
rect 3786 7528 3792 7540
rect 2740 7500 3792 7528
rect 2740 7488 2746 7500
rect 3786 7488 3792 7500
rect 3844 7488 3850 7540
rect 6270 7488 6276 7540
rect 6328 7528 6334 7540
rect 10505 7531 10563 7537
rect 6328 7500 10088 7528
rect 6328 7488 6334 7500
rect 1857 7463 1915 7469
rect 1857 7429 1869 7463
rect 1903 7460 1915 7463
rect 2961 7463 3019 7469
rect 2961 7460 2973 7463
rect 1903 7432 2973 7460
rect 1903 7429 1915 7432
rect 1857 7423 1915 7429
rect 2961 7429 2973 7432
rect 3007 7429 3019 7463
rect 2961 7423 3019 7429
rect 4246 7420 4252 7472
rect 4304 7460 4310 7472
rect 5537 7463 5595 7469
rect 5537 7460 5549 7463
rect 4304 7432 5549 7460
rect 4304 7420 4310 7432
rect 5537 7429 5549 7432
rect 5583 7429 5595 7463
rect 6822 7460 6828 7472
rect 5537 7423 5595 7429
rect 5644 7432 6828 7460
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7392 2099 7395
rect 2130 7392 2136 7404
rect 2087 7364 2136 7392
rect 2087 7361 2099 7364
rect 2041 7355 2099 7361
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 2774 7392 2780 7404
rect 2746 7352 2780 7392
rect 2832 7392 2838 7404
rect 3145 7395 3203 7401
rect 3145 7392 3157 7395
rect 2832 7364 3157 7392
rect 2832 7352 2838 7364
rect 3145 7361 3157 7364
rect 3191 7361 3203 7395
rect 3145 7355 3203 7361
rect 3234 7352 3240 7404
rect 3292 7392 3298 7404
rect 3513 7395 3571 7401
rect 3292 7364 3337 7392
rect 3292 7352 3298 7364
rect 3513 7361 3525 7395
rect 3559 7392 3571 7395
rect 3694 7392 3700 7404
rect 3559 7364 3700 7392
rect 3559 7361 3571 7364
rect 3513 7355 3571 7361
rect 3694 7352 3700 7364
rect 3752 7352 3758 7404
rect 4338 7392 4344 7404
rect 4299 7364 4344 7392
rect 4338 7352 4344 7364
rect 4396 7352 4402 7404
rect 5258 7392 5264 7404
rect 5219 7364 5264 7392
rect 5258 7352 5264 7364
rect 5316 7352 5322 7404
rect 5644 7401 5672 7432
rect 6822 7420 6828 7432
rect 6880 7460 6886 7472
rect 7469 7463 7527 7469
rect 7469 7460 7481 7463
rect 6880 7432 7481 7460
rect 6880 7420 6886 7432
rect 7469 7429 7481 7432
rect 7515 7429 7527 7463
rect 7469 7423 7527 7429
rect 7742 7420 7748 7472
rect 7800 7460 7806 7472
rect 8450 7463 8508 7469
rect 8450 7460 8462 7463
rect 7800 7432 8462 7460
rect 7800 7420 7806 7432
rect 8450 7429 8462 7432
rect 8496 7429 8508 7463
rect 8450 7423 8508 7429
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 5629 7395 5687 7401
rect 5629 7361 5641 7395
rect 5675 7361 5687 7395
rect 6454 7392 6460 7404
rect 6415 7364 6460 7392
rect 5629 7355 5687 7361
rect 2590 7284 2596 7336
rect 2648 7324 2654 7336
rect 2746 7324 2774 7352
rect 2648 7296 2774 7324
rect 2648 7284 2654 7296
rect 2866 7284 2872 7336
rect 2924 7324 2930 7336
rect 5460 7324 5488 7355
rect 6454 7352 6460 7364
rect 6512 7352 6518 7404
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7392 7343 7395
rect 7834 7392 7840 7404
rect 7331 7364 7840 7392
rect 7331 7361 7343 7364
rect 7285 7355 7343 7361
rect 6362 7324 6368 7336
rect 2924 7296 4568 7324
rect 5460 7296 6368 7324
rect 2924 7284 2930 7296
rect 2774 7216 2780 7268
rect 2832 7256 2838 7268
rect 4062 7256 4068 7268
rect 2832 7228 4068 7256
rect 2832 7216 2838 7228
rect 4062 7216 4068 7228
rect 4120 7216 4126 7268
rect 3421 7191 3479 7197
rect 3421 7157 3433 7191
rect 3467 7188 3479 7191
rect 4246 7188 4252 7200
rect 3467 7160 4252 7188
rect 3467 7157 3479 7160
rect 3421 7151 3479 7157
rect 4246 7148 4252 7160
rect 4304 7188 4310 7200
rect 4433 7191 4491 7197
rect 4433 7188 4445 7191
rect 4304 7160 4445 7188
rect 4304 7148 4310 7160
rect 4433 7157 4445 7160
rect 4479 7157 4491 7191
rect 4540 7188 4568 7296
rect 6362 7284 6368 7296
rect 6420 7284 6426 7336
rect 5813 7259 5871 7265
rect 5813 7225 5825 7259
rect 5859 7256 5871 7259
rect 6564 7256 6592 7355
rect 7834 7352 7840 7364
rect 7892 7392 7898 7404
rect 9858 7392 9864 7404
rect 7892 7364 9864 7392
rect 7892 7352 7898 7364
rect 9858 7352 9864 7364
rect 9916 7352 9922 7404
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 8202 7324 8208 7336
rect 6972 7296 8208 7324
rect 6972 7284 6978 7296
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 10060 7324 10088 7500
rect 10505 7497 10517 7531
rect 10551 7528 10563 7531
rect 10594 7528 10600 7540
rect 10551 7500 10600 7528
rect 10551 7497 10563 7500
rect 10505 7491 10563 7497
rect 10594 7488 10600 7500
rect 10652 7488 10658 7540
rect 12526 7488 12532 7540
rect 12584 7528 12590 7540
rect 17129 7531 17187 7537
rect 12584 7500 16160 7528
rect 12584 7488 12590 7500
rect 10137 7463 10195 7469
rect 10137 7429 10149 7463
rect 10183 7460 10195 7463
rect 11517 7463 11575 7469
rect 11517 7460 11529 7463
rect 10183 7432 11529 7460
rect 10183 7429 10195 7432
rect 10137 7423 10195 7429
rect 11517 7429 11529 7432
rect 11563 7429 11575 7463
rect 12618 7460 12624 7472
rect 11517 7423 11575 7429
rect 11624 7432 12112 7460
rect 12579 7432 12624 7460
rect 10226 7352 10232 7404
rect 10284 7392 10290 7404
rect 10321 7395 10379 7401
rect 10321 7392 10333 7395
rect 10284 7364 10333 7392
rect 10284 7352 10290 7364
rect 10321 7361 10333 7364
rect 10367 7361 10379 7395
rect 11624 7392 11652 7432
rect 10321 7355 10379 7361
rect 10428 7364 11652 7392
rect 11701 7395 11759 7401
rect 10428 7324 10456 7364
rect 11701 7361 11713 7395
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 10060 7296 10456 7324
rect 11514 7284 11520 7336
rect 11572 7324 11578 7336
rect 11716 7324 11744 7355
rect 11790 7352 11796 7404
rect 11848 7392 11854 7404
rect 12084 7401 12112 7432
rect 12618 7420 12624 7432
rect 12676 7420 12682 7472
rect 14182 7460 14188 7472
rect 13464 7432 14188 7460
rect 13464 7401 13492 7432
rect 14182 7420 14188 7432
rect 14240 7420 14246 7472
rect 16132 7460 16160 7500
rect 17129 7497 17141 7531
rect 17175 7528 17187 7531
rect 17862 7528 17868 7540
rect 17175 7500 17868 7528
rect 17175 7497 17187 7500
rect 17129 7491 17187 7497
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 18877 7531 18935 7537
rect 18877 7497 18889 7531
rect 18923 7528 18935 7531
rect 19242 7528 19248 7540
rect 18923 7500 19248 7528
rect 18923 7497 18935 7500
rect 18877 7491 18935 7497
rect 19242 7488 19248 7500
rect 19300 7488 19306 7540
rect 20622 7488 20628 7540
rect 20680 7528 20686 7540
rect 23658 7528 23664 7540
rect 20680 7500 21680 7528
rect 20680 7488 20686 7500
rect 16132 7432 16252 7460
rect 12069 7395 12127 7401
rect 11848 7364 11893 7392
rect 11848 7352 11854 7364
rect 12069 7361 12081 7395
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 13449 7395 13507 7401
rect 13449 7361 13461 7395
rect 13495 7361 13507 7395
rect 13449 7355 13507 7361
rect 13538 7352 13544 7404
rect 13596 7392 13602 7404
rect 14093 7395 14151 7401
rect 14093 7392 14105 7395
rect 13596 7364 14105 7392
rect 13596 7352 13602 7364
rect 14093 7361 14105 7364
rect 14139 7361 14151 7395
rect 14093 7355 14151 7361
rect 14737 7395 14795 7401
rect 14737 7361 14749 7395
rect 14783 7392 14795 7395
rect 15194 7392 15200 7404
rect 14783 7364 15200 7392
rect 14783 7361 14795 7364
rect 14737 7355 14795 7361
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 15289 7395 15347 7401
rect 15289 7361 15301 7395
rect 15335 7361 15347 7395
rect 16114 7392 16120 7404
rect 16075 7364 16120 7392
rect 15289 7355 15347 7361
rect 11572 7296 11744 7324
rect 11977 7327 12035 7333
rect 11572 7284 11578 7296
rect 11977 7293 11989 7327
rect 12023 7324 12035 7327
rect 12342 7324 12348 7336
rect 12023 7296 12348 7324
rect 12023 7293 12035 7296
rect 11977 7287 12035 7293
rect 5859 7228 6592 7256
rect 5859 7225 5871 7228
rect 5813 7219 5871 7225
rect 9398 7216 9404 7268
rect 9456 7256 9462 7268
rect 11992 7256 12020 7287
rect 12342 7284 12348 7296
rect 12400 7324 12406 7336
rect 15304 7324 15332 7355
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 16224 7392 16252 7432
rect 16574 7420 16580 7472
rect 16632 7460 16638 7472
rect 17957 7463 18015 7469
rect 17957 7460 17969 7463
rect 16632 7432 17969 7460
rect 16632 7420 16638 7432
rect 17957 7429 17969 7432
rect 18003 7429 18015 7463
rect 21542 7460 21548 7472
rect 17957 7423 18015 7429
rect 19168 7432 21548 7460
rect 16758 7392 16764 7404
rect 16224 7364 16620 7392
rect 16719 7364 16764 7392
rect 12400 7296 15332 7324
rect 15473 7327 15531 7333
rect 12400 7284 12406 7296
rect 15473 7293 15485 7327
rect 15519 7324 15531 7327
rect 15654 7324 15660 7336
rect 15519 7296 15660 7324
rect 15519 7293 15531 7296
rect 15473 7287 15531 7293
rect 15654 7284 15660 7296
rect 15712 7284 15718 7336
rect 16592 7324 16620 7364
rect 16758 7352 16764 7364
rect 16816 7352 16822 7404
rect 16942 7392 16948 7404
rect 16903 7364 16948 7392
rect 16942 7352 16948 7364
rect 17000 7352 17006 7404
rect 17586 7392 17592 7404
rect 17547 7364 17592 7392
rect 17586 7352 17592 7364
rect 17644 7352 17650 7404
rect 17773 7395 17831 7401
rect 17773 7361 17785 7395
rect 17819 7361 17831 7395
rect 19058 7392 19064 7404
rect 19019 7364 19064 7392
rect 17773 7355 17831 7361
rect 17788 7324 17816 7355
rect 19058 7352 19064 7364
rect 19116 7352 19122 7404
rect 19168 7401 19196 7432
rect 21542 7420 21548 7432
rect 21600 7420 21606 7472
rect 21652 7460 21680 7500
rect 22296 7500 23664 7528
rect 22296 7469 22324 7500
rect 23658 7488 23664 7500
rect 23716 7488 23722 7540
rect 23958 7531 24016 7537
rect 23958 7497 23970 7531
rect 24004 7497 24016 7531
rect 23958 7491 24016 7497
rect 24121 7531 24179 7537
rect 24121 7497 24133 7531
rect 24167 7528 24179 7531
rect 24210 7528 24216 7540
rect 24167 7500 24216 7528
rect 24167 7497 24179 7500
rect 24121 7491 24179 7497
rect 22281 7463 22339 7469
rect 21652 7432 22232 7460
rect 19153 7395 19211 7401
rect 19153 7361 19165 7395
rect 19199 7361 19211 7395
rect 19426 7392 19432 7404
rect 19387 7364 19432 7392
rect 19153 7355 19211 7361
rect 19426 7352 19432 7364
rect 19484 7352 19490 7404
rect 19610 7352 19616 7404
rect 19668 7392 19674 7404
rect 19889 7395 19947 7401
rect 19889 7392 19901 7395
rect 19668 7364 19901 7392
rect 19668 7352 19674 7364
rect 19889 7361 19901 7364
rect 19935 7361 19947 7395
rect 19889 7355 19947 7361
rect 20073 7395 20131 7401
rect 20073 7361 20085 7395
rect 20119 7361 20131 7395
rect 20073 7355 20131 7361
rect 19334 7324 19340 7336
rect 16592 7296 19340 7324
rect 16776 7268 16804 7296
rect 19334 7284 19340 7296
rect 19392 7324 19398 7336
rect 20088 7324 20116 7355
rect 20162 7352 20168 7404
rect 20220 7392 20226 7404
rect 20438 7392 20444 7404
rect 20220 7364 20444 7392
rect 20220 7352 20226 7364
rect 20438 7352 20444 7364
rect 20496 7352 20502 7404
rect 20898 7392 20904 7404
rect 20859 7364 20904 7392
rect 20898 7352 20904 7364
rect 20956 7352 20962 7404
rect 19392 7296 20116 7324
rect 19392 7284 19398 7296
rect 9456 7228 12020 7256
rect 13265 7259 13323 7265
rect 9456 7216 9462 7228
rect 13265 7225 13277 7259
rect 13311 7256 13323 7259
rect 16298 7256 16304 7268
rect 13311 7228 16304 7256
rect 13311 7225 13323 7228
rect 13265 7219 13323 7225
rect 16298 7216 16304 7228
rect 16356 7216 16362 7268
rect 16758 7216 16764 7268
rect 16816 7216 16822 7268
rect 17862 7216 17868 7268
rect 17920 7256 17926 7268
rect 20257 7259 20315 7265
rect 20257 7256 20269 7259
rect 17920 7228 20269 7256
rect 17920 7216 17926 7228
rect 20257 7225 20269 7228
rect 20303 7225 20315 7259
rect 20257 7219 20315 7225
rect 6733 7191 6791 7197
rect 6733 7188 6745 7191
rect 4540 7160 6745 7188
rect 4433 7151 4491 7157
rect 6733 7157 6745 7160
rect 6779 7157 6791 7191
rect 9582 7188 9588 7200
rect 9543 7160 9588 7188
rect 6733 7151 6791 7157
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 12526 7148 12532 7200
rect 12584 7188 12590 7200
rect 12713 7191 12771 7197
rect 12713 7188 12725 7191
rect 12584 7160 12725 7188
rect 12584 7148 12590 7160
rect 12713 7157 12725 7160
rect 12759 7157 12771 7191
rect 13906 7188 13912 7200
rect 13867 7160 13912 7188
rect 12713 7151 12771 7157
rect 13906 7148 13912 7160
rect 13964 7148 13970 7200
rect 14553 7191 14611 7197
rect 14553 7157 14565 7191
rect 14599 7188 14611 7191
rect 15286 7188 15292 7200
rect 14599 7160 15292 7188
rect 14599 7157 14611 7160
rect 14553 7151 14611 7157
rect 15286 7148 15292 7160
rect 15344 7148 15350 7200
rect 15470 7148 15476 7200
rect 15528 7188 15534 7200
rect 15933 7191 15991 7197
rect 15933 7188 15945 7191
rect 15528 7160 15945 7188
rect 15528 7148 15534 7160
rect 15933 7157 15945 7160
rect 15979 7157 15991 7191
rect 15933 7151 15991 7157
rect 16390 7148 16396 7200
rect 16448 7188 16454 7200
rect 19058 7188 19064 7200
rect 16448 7160 19064 7188
rect 16448 7148 16454 7160
rect 19058 7148 19064 7160
rect 19116 7148 19122 7200
rect 19334 7188 19340 7200
rect 19295 7160 19340 7188
rect 19334 7148 19340 7160
rect 19392 7148 19398 7200
rect 20438 7148 20444 7200
rect 20496 7188 20502 7200
rect 20717 7191 20775 7197
rect 20717 7188 20729 7191
rect 20496 7160 20729 7188
rect 20496 7148 20502 7160
rect 20717 7157 20729 7160
rect 20763 7157 20775 7191
rect 22204 7188 22232 7432
rect 22281 7429 22293 7463
rect 22327 7429 22339 7463
rect 23750 7460 23756 7472
rect 23711 7432 23756 7460
rect 22281 7423 22339 7429
rect 23750 7420 23756 7432
rect 23808 7420 23814 7472
rect 23973 7460 24001 7491
rect 24210 7488 24216 7500
rect 24268 7488 24274 7540
rect 24949 7531 25007 7537
rect 24949 7497 24961 7531
rect 24995 7497 25007 7531
rect 24949 7491 25007 7497
rect 24302 7460 24308 7472
rect 23973 7432 24308 7460
rect 24302 7420 24308 7432
rect 24360 7420 24366 7472
rect 24578 7460 24584 7472
rect 24539 7432 24584 7460
rect 24578 7420 24584 7432
rect 24636 7420 24642 7472
rect 24811 7429 24869 7435
rect 23106 7352 23112 7404
rect 23164 7392 23170 7404
rect 24811 7395 24823 7429
rect 24857 7395 24869 7429
rect 24964 7404 24992 7491
rect 25958 7488 25964 7540
rect 26016 7528 26022 7540
rect 26421 7531 26479 7537
rect 26421 7528 26433 7531
rect 26016 7500 26433 7528
rect 26016 7488 26022 7500
rect 26421 7497 26433 7500
rect 26467 7497 26479 7531
rect 27154 7528 27160 7540
rect 27212 7537 27218 7540
rect 27212 7531 27241 7537
rect 26421 7491 26479 7497
rect 26528 7500 27160 7528
rect 26053 7463 26111 7469
rect 26053 7429 26065 7463
rect 26099 7429 26111 7463
rect 26053 7423 26111 7429
rect 23164 7364 23209 7392
rect 24811 7389 24869 7395
rect 23164 7352 23170 7364
rect 24302 7284 24308 7336
rect 24360 7324 24366 7336
rect 24812 7324 24840 7389
rect 24946 7352 24952 7404
rect 25004 7352 25010 7404
rect 25498 7352 25504 7404
rect 25556 7392 25562 7404
rect 25593 7395 25651 7401
rect 25593 7392 25605 7395
rect 25556 7364 25605 7392
rect 25556 7352 25562 7364
rect 25593 7361 25605 7364
rect 25639 7361 25651 7395
rect 26068 7392 26096 7423
rect 26142 7420 26148 7472
rect 26200 7460 26206 7472
rect 26269 7463 26327 7469
rect 26269 7460 26281 7463
rect 26200 7432 26281 7460
rect 26200 7420 26206 7432
rect 26269 7429 26281 7432
rect 26315 7460 26327 7463
rect 26528 7460 26556 7500
rect 27154 7488 27160 7500
rect 27229 7528 27241 7531
rect 27522 7528 27528 7540
rect 27229 7500 27528 7528
rect 27229 7497 27241 7500
rect 27212 7491 27241 7497
rect 27212 7488 27218 7491
rect 27522 7488 27528 7500
rect 27580 7488 27586 7540
rect 26315 7432 26556 7460
rect 26315 7429 26327 7432
rect 26269 7423 26327 7429
rect 26878 7420 26884 7472
rect 26936 7460 26942 7472
rect 26973 7463 27031 7469
rect 26973 7460 26985 7463
rect 26936 7432 26985 7460
rect 26936 7420 26942 7432
rect 26973 7429 26985 7432
rect 27019 7429 27031 7463
rect 26973 7423 27031 7429
rect 26694 7392 26700 7404
rect 26068 7364 26700 7392
rect 25593 7355 25651 7361
rect 26694 7352 26700 7364
rect 26752 7392 26758 7404
rect 27338 7392 27344 7404
rect 26752 7364 27344 7392
rect 26752 7352 26758 7364
rect 27338 7352 27344 7364
rect 27396 7352 27402 7404
rect 26142 7324 26148 7336
rect 24360 7296 26148 7324
rect 24360 7284 24366 7296
rect 26142 7284 26148 7296
rect 26200 7284 26206 7336
rect 22462 7216 22468 7268
rect 22520 7256 22526 7268
rect 24210 7256 24216 7268
rect 22520 7228 24216 7256
rect 22520 7216 22526 7228
rect 24210 7216 24216 7228
rect 24268 7216 24274 7268
rect 27062 7216 27068 7268
rect 27120 7256 27126 7268
rect 27341 7259 27399 7265
rect 27341 7256 27353 7259
rect 27120 7228 27353 7256
rect 27120 7216 27126 7228
rect 27341 7225 27353 7228
rect 27387 7225 27399 7259
rect 27341 7219 27399 7225
rect 22373 7191 22431 7197
rect 22373 7188 22385 7191
rect 22204 7160 22385 7188
rect 20717 7151 20775 7157
rect 22373 7157 22385 7160
rect 22419 7157 22431 7191
rect 22373 7151 22431 7157
rect 22925 7191 22983 7197
rect 22925 7157 22937 7191
rect 22971 7188 22983 7191
rect 23198 7188 23204 7200
rect 22971 7160 23204 7188
rect 22971 7157 22983 7160
rect 22925 7151 22983 7157
rect 23198 7148 23204 7160
rect 23256 7148 23262 7200
rect 23937 7191 23995 7197
rect 23937 7157 23949 7191
rect 23983 7188 23995 7191
rect 24765 7191 24823 7197
rect 24765 7188 24777 7191
rect 23983 7160 24777 7188
rect 23983 7157 23995 7160
rect 23937 7151 23995 7157
rect 24765 7157 24777 7160
rect 24811 7188 24823 7191
rect 24854 7188 24860 7200
rect 24811 7160 24860 7188
rect 24811 7157 24823 7160
rect 24765 7151 24823 7157
rect 24854 7148 24860 7160
rect 24912 7148 24918 7200
rect 25038 7148 25044 7200
rect 25096 7188 25102 7200
rect 25409 7191 25467 7197
rect 25409 7188 25421 7191
rect 25096 7160 25421 7188
rect 25096 7148 25102 7160
rect 25409 7157 25421 7160
rect 25455 7157 25467 7191
rect 26234 7188 26240 7200
rect 26147 7160 26240 7188
rect 25409 7151 25467 7157
rect 26234 7148 26240 7160
rect 26292 7188 26298 7200
rect 27157 7191 27215 7197
rect 27157 7188 27169 7191
rect 26292 7160 27169 7188
rect 26292 7148 26298 7160
rect 27157 7157 27169 7160
rect 27203 7188 27215 7191
rect 27430 7188 27436 7200
rect 27203 7160 27436 7188
rect 27203 7157 27215 7160
rect 27157 7151 27215 7157
rect 27430 7148 27436 7160
rect 27488 7148 27494 7200
rect 1104 7098 28060 7120
rect 1104 7046 5442 7098
rect 5494 7046 5506 7098
rect 5558 7046 5570 7098
rect 5622 7046 5634 7098
rect 5686 7046 5698 7098
rect 5750 7046 14428 7098
rect 14480 7046 14492 7098
rect 14544 7046 14556 7098
rect 14608 7046 14620 7098
rect 14672 7046 14684 7098
rect 14736 7046 23413 7098
rect 23465 7046 23477 7098
rect 23529 7046 23541 7098
rect 23593 7046 23605 7098
rect 23657 7046 23669 7098
rect 23721 7046 28060 7098
rect 1104 7024 28060 7046
rect 2590 6944 2596 6996
rect 2648 6984 2654 6996
rect 2958 6984 2964 6996
rect 2648 6956 2964 6984
rect 2648 6944 2654 6956
rect 2958 6944 2964 6956
rect 3016 6944 3022 6996
rect 6362 6944 6368 6996
rect 6420 6984 6426 6996
rect 6733 6987 6791 6993
rect 6733 6984 6745 6987
rect 6420 6956 6745 6984
rect 6420 6944 6426 6956
rect 6733 6953 6745 6956
rect 6779 6953 6791 6987
rect 11054 6984 11060 6996
rect 6733 6947 6791 6953
rect 8220 6956 11060 6984
rect 7006 6916 7012 6928
rect 3988 6888 7012 6916
rect 3602 6808 3608 6860
rect 3660 6848 3666 6860
rect 3789 6851 3847 6857
rect 3789 6848 3801 6851
rect 3660 6820 3801 6848
rect 3660 6808 3666 6820
rect 3789 6817 3801 6820
rect 3835 6817 3847 6851
rect 3789 6811 3847 6817
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6780 3295 6783
rect 3988 6780 4016 6888
rect 7006 6876 7012 6888
rect 7064 6876 7070 6928
rect 7742 6848 7748 6860
rect 7576 6820 7748 6848
rect 3283 6752 4016 6780
rect 4065 6783 4123 6789
rect 3283 6749 3295 6752
rect 3237 6743 3295 6749
rect 4065 6749 4077 6783
rect 4111 6780 4123 6783
rect 5261 6783 5319 6789
rect 5261 6780 5273 6783
rect 4111 6752 5273 6780
rect 4111 6749 4123 6752
rect 4065 6743 4123 6749
rect 5261 6749 5273 6752
rect 5307 6749 5319 6783
rect 5261 6743 5319 6749
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6780 6147 6783
rect 6564 6780 6776 6796
rect 7576 6789 7604 6820
rect 7742 6808 7748 6820
rect 7800 6848 7806 6860
rect 8220 6848 8248 6956
rect 11054 6944 11060 6956
rect 11112 6944 11118 6996
rect 12710 6984 12716 6996
rect 12623 6956 12716 6984
rect 12710 6944 12716 6956
rect 12768 6984 12774 6996
rect 13538 6984 13544 6996
rect 12768 6956 13544 6984
rect 12768 6944 12774 6956
rect 13538 6944 13544 6956
rect 13596 6944 13602 6996
rect 14918 6944 14924 6996
rect 14976 6984 14982 6996
rect 15746 6984 15752 6996
rect 14976 6956 15752 6984
rect 14976 6944 14982 6956
rect 15746 6944 15752 6956
rect 15804 6944 15810 6996
rect 21174 6984 21180 6996
rect 20548 6956 21180 6984
rect 9214 6916 9220 6928
rect 8956 6888 9220 6916
rect 8956 6857 8984 6888
rect 9214 6876 9220 6888
rect 9272 6876 9278 6928
rect 9490 6876 9496 6928
rect 9548 6916 9554 6928
rect 10226 6916 10232 6928
rect 9548 6888 10232 6916
rect 9548 6876 9554 6888
rect 10226 6876 10232 6888
rect 10284 6876 10290 6928
rect 12986 6876 12992 6928
rect 13044 6916 13050 6928
rect 13354 6916 13360 6928
rect 13044 6888 13360 6916
rect 13044 6876 13050 6888
rect 13354 6876 13360 6888
rect 13412 6876 13418 6928
rect 19334 6876 19340 6928
rect 19392 6916 19398 6928
rect 19705 6919 19763 6925
rect 19705 6916 19717 6919
rect 19392 6888 19717 6916
rect 19392 6876 19398 6888
rect 19705 6885 19717 6888
rect 19751 6885 19763 6919
rect 19705 6879 19763 6885
rect 7800 6820 8248 6848
rect 8941 6851 8999 6857
rect 7800 6808 7806 6820
rect 8941 6817 8953 6851
rect 8987 6817 8999 6851
rect 10410 6848 10416 6860
rect 8941 6811 8999 6817
rect 9048 6820 10416 6848
rect 7561 6783 7619 6789
rect 6135 6768 7512 6780
rect 6135 6752 6592 6768
rect 6748 6752 7512 6768
rect 6135 6749 6147 6752
rect 6089 6743 6147 6749
rect 1946 6712 1952 6724
rect 1907 6684 1952 6712
rect 1946 6672 1952 6684
rect 2004 6672 2010 6724
rect 2133 6715 2191 6721
rect 2133 6681 2145 6715
rect 2179 6712 2191 6715
rect 3602 6712 3608 6724
rect 2179 6684 3608 6712
rect 2179 6681 2191 6684
rect 2133 6675 2191 6681
rect 3602 6672 3608 6684
rect 3660 6712 3666 6724
rect 4080 6712 4108 6743
rect 5074 6712 5080 6724
rect 3660 6684 4108 6712
rect 5035 6684 5080 6712
rect 3660 6672 3666 6684
rect 5074 6672 5080 6684
rect 5132 6672 5138 6724
rect 5445 6715 5503 6721
rect 5445 6681 5457 6715
rect 5491 6712 5503 6715
rect 6546 6712 6552 6724
rect 5491 6684 6552 6712
rect 5491 6681 5503 6684
rect 5445 6675 5503 6681
rect 6546 6672 6552 6684
rect 6604 6672 6610 6724
rect 6641 6715 6699 6721
rect 6641 6681 6653 6715
rect 6687 6712 6699 6715
rect 7006 6712 7012 6724
rect 6687 6684 7012 6712
rect 6687 6681 6699 6684
rect 6641 6675 6699 6681
rect 7006 6672 7012 6684
rect 7064 6712 7070 6724
rect 7484 6712 7512 6752
rect 7561 6749 7573 6783
rect 7607 6749 7619 6783
rect 7834 6780 7840 6792
rect 7795 6752 7840 6780
rect 7561 6743 7619 6749
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 8202 6740 8208 6792
rect 8260 6780 8266 6792
rect 9048 6780 9076 6820
rect 10410 6808 10416 6820
rect 10468 6808 10474 6860
rect 13722 6848 13728 6860
rect 12820 6820 13728 6848
rect 9214 6780 9220 6792
rect 8260 6752 9076 6780
rect 9175 6752 9220 6780
rect 8260 6740 8266 6752
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 10680 6783 10738 6789
rect 10680 6749 10692 6783
rect 10726 6780 10738 6783
rect 12342 6780 12348 6792
rect 10726 6752 12348 6780
rect 10726 6749 10738 6752
rect 10680 6743 10738 6749
rect 12342 6740 12348 6752
rect 12400 6740 12406 6792
rect 12618 6789 12624 6792
rect 12437 6783 12495 6789
rect 12437 6749 12449 6783
rect 12483 6749 12495 6783
rect 12437 6743 12495 6749
rect 12589 6783 12624 6789
rect 12589 6749 12601 6783
rect 12589 6743 12624 6749
rect 11698 6712 11704 6724
rect 7064 6684 7144 6712
rect 7484 6684 11704 6712
rect 7064 6672 7070 6684
rect 2314 6644 2320 6656
rect 2275 6616 2320 6644
rect 2314 6604 2320 6616
rect 2372 6604 2378 6656
rect 3053 6647 3111 6653
rect 3053 6613 3065 6647
rect 3099 6644 3111 6647
rect 3326 6644 3332 6656
rect 3099 6616 3332 6644
rect 3099 6613 3111 6616
rect 3053 6607 3111 6613
rect 3326 6604 3332 6616
rect 3384 6604 3390 6656
rect 5902 6644 5908 6656
rect 5863 6616 5908 6644
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 7116 6644 7144 6684
rect 11698 6672 11704 6684
rect 11756 6672 11762 6724
rect 12452 6712 12480 6743
rect 12618 6740 12624 6743
rect 12676 6740 12682 6792
rect 12820 6789 12848 6820
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 19245 6851 19303 6857
rect 19245 6817 19257 6851
rect 19291 6848 19303 6851
rect 19610 6848 19616 6860
rect 19291 6820 19616 6848
rect 19291 6817 19303 6820
rect 19245 6811 19303 6817
rect 19610 6808 19616 6820
rect 19668 6808 19674 6860
rect 20548 6848 20576 6956
rect 21174 6944 21180 6956
rect 21232 6944 21238 6996
rect 24394 6944 24400 6996
rect 24452 6984 24458 6996
rect 24581 6987 24639 6993
rect 24581 6984 24593 6987
rect 24452 6956 24593 6984
rect 24452 6944 24458 6956
rect 24581 6953 24593 6956
rect 24627 6984 24639 6987
rect 24670 6984 24676 6996
rect 24627 6956 24676 6984
rect 24627 6953 24639 6956
rect 24581 6947 24639 6953
rect 24670 6944 24676 6956
rect 24728 6944 24734 6996
rect 24854 6944 24860 6996
rect 24912 6984 24918 6996
rect 26234 6984 26240 6996
rect 24912 6956 26240 6984
rect 24912 6944 24918 6956
rect 26234 6944 26240 6956
rect 26292 6944 26298 6996
rect 27338 6984 27344 6996
rect 27299 6956 27344 6984
rect 27338 6944 27344 6956
rect 27396 6944 27402 6996
rect 22646 6876 22652 6928
rect 22704 6916 22710 6928
rect 24765 6919 24823 6925
rect 24765 6916 24777 6919
rect 22704 6888 24777 6916
rect 22704 6876 22710 6888
rect 24765 6885 24777 6888
rect 24811 6885 24823 6919
rect 24765 6879 24823 6885
rect 19812 6820 20576 6848
rect 12805 6783 12863 6789
rect 12805 6749 12817 6783
rect 12851 6749 12863 6783
rect 12805 6743 12863 6749
rect 12894 6740 12900 6792
rect 12952 6780 12958 6792
rect 13449 6783 13507 6789
rect 13449 6780 13461 6783
rect 12952 6752 13461 6780
rect 12952 6740 12958 6752
rect 13449 6749 13461 6752
rect 13495 6749 13507 6783
rect 13449 6743 13507 6749
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 14918 6780 14924 6792
rect 14599 6752 14924 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 14918 6740 14924 6752
rect 14976 6740 14982 6792
rect 15013 6783 15071 6789
rect 15013 6749 15025 6783
rect 15059 6780 15071 6783
rect 17221 6783 17279 6789
rect 17221 6780 17233 6783
rect 15059 6752 17233 6780
rect 15059 6749 15071 6752
rect 15013 6743 15071 6749
rect 17221 6749 17233 6752
rect 17267 6780 17279 6783
rect 17310 6780 17316 6792
rect 17267 6752 17316 6780
rect 17267 6749 17279 6752
rect 17221 6743 17279 6749
rect 12710 6712 12716 6724
rect 12452 6684 12716 6712
rect 12710 6672 12716 6684
rect 12768 6672 12774 6724
rect 14274 6672 14280 6724
rect 14332 6712 14338 6724
rect 15028 6712 15056 6743
rect 17310 6740 17316 6752
rect 17368 6740 17374 6792
rect 17494 6789 17500 6792
rect 17488 6743 17500 6789
rect 17552 6780 17558 6792
rect 17552 6752 17588 6780
rect 17494 6740 17500 6743
rect 17552 6740 17558 6752
rect 19058 6740 19064 6792
rect 19116 6780 19122 6792
rect 19429 6783 19487 6789
rect 19429 6780 19441 6783
rect 19116 6752 19441 6780
rect 19116 6740 19122 6752
rect 19429 6749 19441 6752
rect 19475 6749 19487 6783
rect 19429 6743 19487 6749
rect 19521 6783 19579 6789
rect 19521 6749 19533 6783
rect 19567 6780 19579 6783
rect 19702 6780 19708 6792
rect 19567 6752 19708 6780
rect 19567 6749 19579 6752
rect 19521 6743 19579 6749
rect 19702 6740 19708 6752
rect 19760 6740 19766 6792
rect 19812 6789 19840 6820
rect 21634 6808 21640 6860
rect 21692 6848 21698 6860
rect 21692 6820 22876 6848
rect 21692 6808 21698 6820
rect 19797 6783 19855 6789
rect 19797 6749 19809 6783
rect 19843 6749 19855 6783
rect 19797 6743 19855 6749
rect 19886 6740 19892 6792
rect 19944 6780 19950 6792
rect 20533 6783 20591 6789
rect 20533 6780 20545 6783
rect 19944 6752 20545 6780
rect 19944 6740 19950 6752
rect 20533 6749 20545 6752
rect 20579 6780 20591 6783
rect 22186 6780 22192 6792
rect 20579 6752 22192 6780
rect 20579 6749 20591 6752
rect 20533 6743 20591 6749
rect 22186 6740 22192 6752
rect 22244 6740 22250 6792
rect 22848 6789 22876 6820
rect 25498 6808 25504 6860
rect 25556 6848 25562 6860
rect 25961 6851 26019 6857
rect 25961 6848 25973 6851
rect 25556 6820 25973 6848
rect 25556 6808 25562 6820
rect 25961 6817 25973 6820
rect 26007 6817 26019 6851
rect 25961 6811 26019 6817
rect 22833 6783 22891 6789
rect 22833 6749 22845 6783
rect 22879 6749 22891 6783
rect 22833 6743 22891 6749
rect 23569 6783 23627 6789
rect 23569 6749 23581 6783
rect 23615 6780 23627 6783
rect 24026 6780 24032 6792
rect 23615 6752 24032 6780
rect 23615 6749 23627 6752
rect 23569 6743 23627 6749
rect 24026 6740 24032 6752
rect 24084 6740 24090 6792
rect 24210 6740 24216 6792
rect 24268 6780 24274 6792
rect 25225 6783 25283 6789
rect 25225 6780 25237 6783
rect 24268 6752 25237 6780
rect 24268 6740 24274 6752
rect 25225 6749 25237 6752
rect 25271 6749 25283 6783
rect 25225 6743 25283 6749
rect 15286 6721 15292 6724
rect 15280 6712 15292 6721
rect 14332 6684 15056 6712
rect 15247 6684 15292 6712
rect 14332 6672 14338 6684
rect 15280 6675 15292 6684
rect 15286 6672 15292 6675
rect 15344 6672 15350 6724
rect 15562 6672 15568 6724
rect 15620 6712 15626 6724
rect 20778 6715 20836 6721
rect 20778 6712 20790 6715
rect 15620 6684 20790 6712
rect 15620 6672 15626 6684
rect 20778 6681 20790 6684
rect 20824 6681 20836 6715
rect 20778 6675 20836 6681
rect 21818 6672 21824 6724
rect 21876 6712 21882 6724
rect 24394 6712 24400 6724
rect 21876 6684 24164 6712
rect 24355 6684 24400 6712
rect 21876 6672 21882 6684
rect 10594 6644 10600 6656
rect 7116 6616 10600 6644
rect 10594 6604 10600 6616
rect 10652 6604 10658 6656
rect 11790 6644 11796 6656
rect 11751 6616 11796 6644
rect 11790 6604 11796 6616
rect 11848 6604 11854 6656
rect 12253 6647 12311 6653
rect 12253 6613 12265 6647
rect 12299 6644 12311 6647
rect 12434 6644 12440 6656
rect 12299 6616 12440 6644
rect 12299 6613 12311 6616
rect 12253 6607 12311 6613
rect 12434 6604 12440 6616
rect 12492 6604 12498 6656
rect 13262 6644 13268 6656
rect 13223 6616 13268 6644
rect 13262 6604 13268 6616
rect 13320 6604 13326 6656
rect 14369 6647 14427 6653
rect 14369 6613 14381 6647
rect 14415 6644 14427 6647
rect 14918 6644 14924 6656
rect 14415 6616 14924 6644
rect 14415 6613 14427 6616
rect 14369 6607 14427 6613
rect 14918 6604 14924 6616
rect 14976 6604 14982 6656
rect 15930 6604 15936 6656
rect 15988 6644 15994 6656
rect 16393 6647 16451 6653
rect 16393 6644 16405 6647
rect 15988 6616 16405 6644
rect 15988 6604 15994 6616
rect 16393 6613 16405 6616
rect 16439 6613 16451 6647
rect 16393 6607 16451 6613
rect 17862 6604 17868 6656
rect 17920 6644 17926 6656
rect 18601 6647 18659 6653
rect 18601 6644 18613 6647
rect 17920 6616 18613 6644
rect 17920 6604 17926 6616
rect 18601 6613 18613 6616
rect 18647 6613 18659 6647
rect 18601 6607 18659 6613
rect 21913 6647 21971 6653
rect 21913 6613 21925 6647
rect 21959 6644 21971 6647
rect 22002 6644 22008 6656
rect 21959 6616 22008 6644
rect 21959 6613 21971 6616
rect 21913 6607 21971 6613
rect 22002 6604 22008 6616
rect 22060 6604 22066 6656
rect 23014 6644 23020 6656
rect 22975 6616 23020 6644
rect 23014 6604 23020 6616
rect 23072 6604 23078 6656
rect 23753 6647 23811 6653
rect 23753 6613 23765 6647
rect 23799 6644 23811 6647
rect 24026 6644 24032 6656
rect 23799 6616 24032 6644
rect 23799 6613 23811 6616
rect 23753 6607 23811 6613
rect 24026 6604 24032 6616
rect 24084 6604 24090 6656
rect 24136 6644 24164 6684
rect 24394 6672 24400 6684
rect 24452 6672 24458 6724
rect 26206 6715 26264 6721
rect 26206 6712 26218 6715
rect 24504 6684 26218 6712
rect 24504 6644 24532 6684
rect 26206 6681 26218 6684
rect 26252 6681 26264 6715
rect 26206 6675 26264 6681
rect 24136 6616 24532 6644
rect 24607 6647 24665 6653
rect 24607 6613 24619 6647
rect 24653 6644 24665 6647
rect 24762 6644 24768 6656
rect 24653 6616 24768 6644
rect 24653 6613 24665 6616
rect 24607 6607 24665 6613
rect 24762 6604 24768 6616
rect 24820 6604 24826 6656
rect 24946 6604 24952 6656
rect 25004 6644 25010 6656
rect 25409 6647 25467 6653
rect 25409 6644 25421 6647
rect 25004 6616 25421 6644
rect 25004 6604 25010 6616
rect 25409 6613 25421 6616
rect 25455 6613 25467 6647
rect 25409 6607 25467 6613
rect 1104 6554 28060 6576
rect 1104 6502 9935 6554
rect 9987 6502 9999 6554
rect 10051 6502 10063 6554
rect 10115 6502 10127 6554
rect 10179 6502 10191 6554
rect 10243 6502 18920 6554
rect 18972 6502 18984 6554
rect 19036 6502 19048 6554
rect 19100 6502 19112 6554
rect 19164 6502 19176 6554
rect 19228 6502 28060 6554
rect 1104 6480 28060 6502
rect 3329 6443 3387 6449
rect 3329 6440 3341 6443
rect 3160 6412 3341 6440
rect 1756 6375 1814 6381
rect 1756 6341 1768 6375
rect 1802 6372 1814 6375
rect 3160 6372 3188 6412
rect 3329 6409 3341 6412
rect 3375 6409 3387 6443
rect 3329 6403 3387 6409
rect 5350 6400 5356 6452
rect 5408 6440 5414 6452
rect 5445 6443 5503 6449
rect 5445 6440 5457 6443
rect 5408 6412 5457 6440
rect 5408 6400 5414 6412
rect 5445 6409 5457 6412
rect 5491 6409 5503 6443
rect 5445 6403 5503 6409
rect 8938 6400 8944 6452
rect 8996 6440 9002 6452
rect 9125 6443 9183 6449
rect 9125 6440 9137 6443
rect 8996 6412 9137 6440
rect 8996 6400 9002 6412
rect 9125 6409 9137 6412
rect 9171 6409 9183 6443
rect 9125 6403 9183 6409
rect 9674 6400 9680 6452
rect 9732 6440 9738 6452
rect 10505 6443 10563 6449
rect 10505 6440 10517 6443
rect 9732 6412 10517 6440
rect 9732 6400 9738 6412
rect 10505 6409 10517 6412
rect 10551 6409 10563 6443
rect 10505 6403 10563 6409
rect 15286 6400 15292 6452
rect 15344 6440 15350 6452
rect 16025 6443 16083 6449
rect 16025 6440 16037 6443
rect 15344 6412 16037 6440
rect 15344 6400 15350 6412
rect 16025 6409 16037 6412
rect 16071 6409 16083 6443
rect 16025 6403 16083 6409
rect 16666 6400 16672 6452
rect 16724 6400 16730 6452
rect 16945 6443 17003 6449
rect 16945 6409 16957 6443
rect 16991 6440 17003 6443
rect 17586 6440 17592 6452
rect 16991 6412 17592 6440
rect 16991 6409 17003 6412
rect 16945 6403 17003 6409
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 17862 6400 17868 6452
rect 17920 6440 17926 6452
rect 22554 6440 22560 6452
rect 17920 6412 22560 6440
rect 17920 6400 17926 6412
rect 22554 6400 22560 6412
rect 22612 6400 22618 6452
rect 24302 6440 24308 6452
rect 23860 6412 24072 6440
rect 24263 6412 24308 6440
rect 6914 6372 6920 6384
rect 1802 6344 3188 6372
rect 6380 6344 6920 6372
rect 1802 6341 1814 6344
rect 1756 6335 1814 6341
rect 1578 6304 1584 6316
rect 1504 6276 1584 6304
rect 1394 6196 1400 6248
rect 1452 6236 1458 6248
rect 1504 6245 1532 6276
rect 1578 6264 1584 6276
rect 1636 6264 1642 6316
rect 2314 6264 2320 6316
rect 2372 6304 2378 6316
rect 3513 6307 3571 6313
rect 3513 6304 3525 6307
rect 2372 6276 3525 6304
rect 2372 6264 2378 6276
rect 3513 6273 3525 6276
rect 3559 6273 3571 6307
rect 3513 6267 3571 6273
rect 4332 6307 4390 6313
rect 4332 6273 4344 6307
rect 4378 6304 4390 6307
rect 6270 6304 6276 6316
rect 4378 6276 6276 6304
rect 4378 6273 4390 6276
rect 4332 6267 4390 6273
rect 6270 6264 6276 6276
rect 6328 6264 6334 6316
rect 6380 6313 6408 6344
rect 6914 6332 6920 6344
rect 6972 6332 6978 6384
rect 8478 6372 8484 6384
rect 8439 6344 8484 6372
rect 8478 6332 8484 6344
rect 8536 6332 8542 6384
rect 11054 6372 11060 6384
rect 8956 6344 9720 6372
rect 8956 6316 8984 6344
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6273 6423 6307
rect 6621 6307 6679 6313
rect 6621 6304 6633 6307
rect 6365 6267 6423 6273
rect 6472 6276 6633 6304
rect 1489 6239 1547 6245
rect 1489 6236 1501 6239
rect 1452 6208 1501 6236
rect 1452 6196 1458 6208
rect 1489 6205 1501 6208
rect 1535 6205 1547 6239
rect 1489 6199 1547 6205
rect 2682 6196 2688 6248
rect 2740 6236 2746 6248
rect 4065 6239 4123 6245
rect 4065 6236 4077 6239
rect 2740 6208 4077 6236
rect 2740 6196 2746 6208
rect 4065 6205 4077 6208
rect 4111 6205 4123 6239
rect 4065 6199 4123 6205
rect 5810 6196 5816 6248
rect 5868 6236 5874 6248
rect 6472 6236 6500 6276
rect 6621 6273 6633 6276
rect 6667 6273 6679 6307
rect 6621 6267 6679 6273
rect 8938 6264 8944 6316
rect 8996 6264 9002 6316
rect 9214 6264 9220 6316
rect 9272 6304 9278 6316
rect 9309 6307 9367 6313
rect 9309 6304 9321 6307
rect 9272 6276 9321 6304
rect 9272 6264 9278 6276
rect 9309 6273 9321 6276
rect 9355 6273 9367 6307
rect 9309 6267 9367 6273
rect 9401 6307 9459 6313
rect 9401 6273 9413 6307
rect 9447 6304 9459 6307
rect 9582 6304 9588 6316
rect 9447 6276 9588 6304
rect 9447 6273 9459 6276
rect 9401 6267 9459 6273
rect 5868 6208 6500 6236
rect 5868 6196 5874 6208
rect 8478 6196 8484 6248
rect 8536 6236 8542 6248
rect 9324 6236 9352 6267
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 9692 6313 9720 6344
rect 9784 6344 11060 6372
rect 9677 6307 9735 6313
rect 9677 6273 9689 6307
rect 9723 6273 9735 6307
rect 9677 6267 9735 6273
rect 9784 6236 9812 6344
rect 11054 6332 11060 6344
rect 11112 6372 11118 6384
rect 11514 6372 11520 6384
rect 11112 6344 11520 6372
rect 11112 6332 11118 6344
rect 11514 6332 11520 6344
rect 11572 6332 11578 6384
rect 12526 6372 12532 6384
rect 12268 6344 12532 6372
rect 9858 6264 9864 6316
rect 9916 6304 9922 6316
rect 10137 6307 10195 6313
rect 10137 6304 10149 6307
rect 9916 6276 10149 6304
rect 9916 6264 9922 6276
rect 10137 6273 10149 6276
rect 10183 6273 10195 6307
rect 10137 6267 10195 6273
rect 10321 6307 10379 6313
rect 10321 6273 10333 6307
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 8536 6208 9812 6236
rect 8536 6196 8542 6208
rect 9490 6128 9496 6180
rect 9548 6168 9554 6180
rect 10336 6168 10364 6267
rect 10410 6264 10416 6316
rect 10468 6304 10474 6316
rect 12268 6304 12296 6344
rect 12526 6332 12532 6344
rect 12584 6372 12590 6384
rect 13072 6375 13130 6381
rect 12584 6344 12848 6372
rect 12584 6332 12590 6344
rect 12820 6313 12848 6344
rect 13072 6341 13084 6375
rect 13118 6372 13130 6375
rect 13262 6372 13268 6384
rect 13118 6344 13268 6372
rect 13118 6341 13130 6344
rect 13072 6335 13130 6341
rect 13262 6332 13268 6344
rect 13320 6332 13326 6384
rect 13354 6332 13360 6384
rect 13412 6372 13418 6384
rect 13906 6372 13912 6384
rect 13412 6344 13912 6372
rect 13412 6332 13418 6344
rect 13906 6332 13912 6344
rect 13964 6332 13970 6384
rect 14645 6375 14703 6381
rect 14645 6341 14657 6375
rect 14691 6372 14703 6375
rect 15657 6375 15715 6381
rect 15657 6372 15669 6375
rect 14691 6344 15669 6372
rect 14691 6341 14703 6344
rect 14645 6335 14703 6341
rect 15657 6341 15669 6344
rect 15703 6341 15715 6375
rect 16206 6372 16212 6384
rect 15657 6335 15715 6341
rect 15764 6344 16212 6372
rect 10468 6276 12296 6304
rect 12805 6307 12863 6313
rect 10468 6264 10474 6276
rect 12805 6273 12817 6307
rect 12851 6273 12863 6307
rect 14826 6304 14832 6316
rect 14787 6276 14832 6304
rect 12805 6267 12863 6273
rect 14826 6264 14832 6276
rect 14884 6264 14890 6316
rect 14921 6307 14979 6313
rect 14921 6273 14933 6307
rect 14967 6273 14979 6307
rect 14921 6267 14979 6273
rect 15179 6308 15237 6313
rect 15179 6307 15323 6308
rect 15179 6273 15191 6307
rect 15225 6304 15323 6307
rect 15764 6304 15792 6344
rect 16206 6332 16212 6344
rect 16264 6332 16270 6384
rect 16684 6372 16712 6400
rect 17954 6372 17960 6384
rect 16684 6344 17264 6372
rect 15225 6280 15792 6304
rect 15225 6276 15240 6280
rect 15295 6276 15792 6280
rect 15841 6307 15899 6313
rect 15225 6273 15237 6276
rect 15179 6267 15237 6273
rect 15841 6273 15853 6307
rect 15887 6273 15899 6307
rect 15841 6267 15899 6273
rect 11514 6236 11520 6248
rect 11475 6208 11520 6236
rect 11514 6196 11520 6208
rect 11572 6196 11578 6248
rect 11793 6239 11851 6245
rect 11793 6205 11805 6239
rect 11839 6236 11851 6239
rect 12710 6236 12716 6248
rect 11839 6208 12716 6236
rect 11839 6205 11851 6208
rect 11793 6199 11851 6205
rect 12710 6196 12716 6208
rect 12768 6196 12774 6248
rect 14734 6196 14740 6248
rect 14792 6236 14798 6248
rect 14936 6236 14964 6267
rect 14792 6208 14964 6236
rect 14792 6196 14798 6208
rect 15286 6196 15292 6248
rect 15344 6236 15350 6248
rect 15856 6236 15884 6267
rect 16390 6264 16396 6316
rect 16448 6304 16454 6316
rect 17236 6313 17264 6344
rect 17512 6344 17960 6372
rect 17512 6313 17540 6344
rect 17954 6332 17960 6344
rect 18012 6332 18018 6384
rect 19702 6332 19708 6384
rect 19760 6372 19766 6384
rect 20162 6381 20168 6384
rect 20156 6372 20168 6381
rect 19760 6344 20024 6372
rect 20123 6344 20168 6372
rect 19760 6332 19766 6344
rect 17129 6307 17187 6313
rect 17129 6304 17141 6307
rect 16448 6276 17141 6304
rect 16448 6264 16454 6276
rect 17129 6273 17141 6276
rect 17175 6273 17187 6307
rect 17129 6267 17187 6273
rect 17221 6307 17279 6313
rect 17221 6273 17233 6307
rect 17267 6273 17279 6307
rect 17221 6267 17279 6273
rect 17497 6307 17555 6313
rect 17497 6273 17509 6307
rect 17543 6273 17555 6307
rect 17497 6267 17555 6273
rect 17586 6264 17592 6316
rect 17644 6304 17650 6316
rect 18141 6307 18199 6313
rect 18141 6304 18153 6307
rect 17644 6276 18153 6304
rect 17644 6264 17650 6276
rect 18141 6273 18153 6276
rect 18187 6273 18199 6307
rect 18141 6267 18199 6273
rect 18414 6264 18420 6316
rect 18472 6304 18478 6316
rect 18785 6307 18843 6313
rect 18785 6304 18797 6307
rect 18472 6276 18797 6304
rect 18472 6264 18478 6276
rect 18785 6273 18797 6276
rect 18831 6273 18843 6307
rect 19426 6304 19432 6316
rect 19387 6276 19432 6304
rect 18785 6267 18843 6273
rect 19426 6264 19432 6276
rect 19484 6264 19490 6316
rect 19886 6304 19892 6316
rect 19847 6276 19892 6304
rect 19886 6264 19892 6276
rect 19944 6264 19950 6316
rect 19996 6304 20024 6344
rect 20156 6335 20168 6344
rect 20162 6332 20168 6335
rect 20220 6332 20226 6384
rect 20714 6332 20720 6384
rect 20772 6372 20778 6384
rect 21634 6372 21640 6384
rect 20772 6344 21640 6372
rect 20772 6332 20778 6344
rect 21634 6332 21640 6344
rect 21692 6332 21698 6384
rect 23860 6372 23888 6412
rect 22204 6344 23888 6372
rect 23937 6375 23995 6381
rect 22204 6316 22232 6344
rect 23937 6341 23949 6375
rect 23983 6341 23995 6375
rect 23937 6335 23995 6341
rect 22002 6304 22008 6316
rect 19996 6276 22008 6304
rect 22002 6264 22008 6276
rect 22060 6264 22066 6316
rect 22097 6307 22155 6313
rect 22097 6273 22109 6307
rect 22143 6304 22155 6307
rect 22186 6304 22192 6316
rect 22143 6276 22192 6304
rect 22143 6273 22155 6276
rect 22097 6267 22155 6273
rect 22186 6264 22192 6276
rect 22244 6264 22250 6316
rect 22364 6307 22422 6313
rect 22364 6273 22376 6307
rect 22410 6304 22422 6307
rect 22646 6304 22652 6316
rect 22410 6276 22652 6304
rect 22410 6273 22422 6276
rect 22364 6267 22422 6273
rect 22646 6264 22652 6276
rect 22704 6264 22710 6316
rect 23943 6304 23971 6335
rect 23492 6276 23971 6304
rect 24044 6304 24072 6412
rect 24302 6400 24308 6412
rect 24360 6400 24366 6452
rect 24762 6400 24768 6452
rect 24820 6400 24826 6452
rect 25222 6400 25228 6452
rect 25280 6440 25286 6452
rect 26234 6440 26240 6452
rect 25280 6412 26240 6440
rect 25280 6400 25286 6412
rect 26234 6400 26240 6412
rect 26292 6400 26298 6452
rect 27154 6400 27160 6452
rect 27212 6449 27218 6452
rect 27212 6443 27231 6449
rect 27219 6409 27231 6443
rect 27338 6440 27344 6452
rect 27299 6412 27344 6440
rect 27212 6403 27231 6409
rect 27212 6400 27218 6403
rect 27338 6400 27344 6412
rect 27396 6400 27402 6452
rect 24210 6381 24216 6384
rect 24153 6375 24216 6381
rect 24153 6341 24165 6375
rect 24199 6341 24216 6375
rect 24153 6335 24216 6341
rect 24210 6332 24216 6335
rect 24268 6372 24274 6384
rect 24780 6372 24808 6400
rect 25038 6381 25044 6384
rect 25032 6372 25044 6381
rect 24268 6344 24808 6372
rect 24999 6344 25044 6372
rect 24268 6332 24274 6344
rect 25032 6335 25044 6344
rect 25038 6332 25044 6335
rect 25096 6332 25102 6384
rect 25958 6332 25964 6384
rect 26016 6372 26022 6384
rect 26973 6375 27031 6381
rect 26973 6372 26985 6375
rect 26016 6344 26985 6372
rect 26016 6332 26022 6344
rect 26973 6341 26985 6344
rect 27019 6341 27031 6375
rect 26973 6335 27031 6341
rect 24762 6304 24768 6316
rect 24044 6276 24768 6304
rect 19334 6236 19340 6248
rect 15344 6208 15884 6236
rect 17420 6208 19340 6236
rect 15344 6196 15350 6208
rect 9548 6140 10364 6168
rect 9548 6128 9554 6140
rect 11974 6128 11980 6180
rect 12032 6128 12038 6180
rect 13740 6140 14320 6168
rect 2774 6060 2780 6112
rect 2832 6100 2838 6112
rect 2869 6103 2927 6109
rect 2869 6100 2881 6103
rect 2832 6072 2881 6100
rect 2832 6060 2838 6072
rect 2869 6069 2881 6072
rect 2915 6100 2927 6103
rect 3050 6100 3056 6112
rect 2915 6072 3056 6100
rect 2915 6069 2927 6072
rect 2869 6063 2927 6069
rect 3050 6060 3056 6072
rect 3108 6060 3114 6112
rect 7006 6060 7012 6112
rect 7064 6100 7070 6112
rect 7745 6103 7803 6109
rect 7745 6100 7757 6103
rect 7064 6072 7757 6100
rect 7064 6060 7070 6072
rect 7745 6069 7757 6072
rect 7791 6069 7803 6103
rect 7745 6063 7803 6069
rect 8202 6060 8208 6112
rect 8260 6100 8266 6112
rect 8573 6103 8631 6109
rect 8573 6100 8585 6103
rect 8260 6072 8585 6100
rect 8260 6060 8266 6072
rect 8573 6069 8585 6072
rect 8619 6100 8631 6103
rect 9398 6100 9404 6112
rect 8619 6072 9404 6100
rect 8619 6069 8631 6072
rect 8573 6063 8631 6069
rect 9398 6060 9404 6072
rect 9456 6100 9462 6112
rect 9585 6103 9643 6109
rect 9585 6100 9597 6103
rect 9456 6072 9597 6100
rect 9456 6060 9462 6072
rect 9585 6069 9597 6072
rect 9631 6069 9643 6103
rect 9585 6063 9643 6069
rect 10962 6060 10968 6112
rect 11020 6100 11026 6112
rect 11698 6100 11704 6112
rect 11020 6072 11704 6100
rect 11020 6060 11026 6072
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 11992 6100 12020 6128
rect 13740 6112 13768 6140
rect 12158 6100 12164 6112
rect 11992 6072 12164 6100
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 13538 6060 13544 6112
rect 13596 6100 13602 6112
rect 13722 6100 13728 6112
rect 13596 6072 13728 6100
rect 13596 6060 13602 6072
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 13906 6060 13912 6112
rect 13964 6100 13970 6112
rect 14185 6103 14243 6109
rect 14185 6100 14197 6103
rect 13964 6072 14197 6100
rect 13964 6060 13970 6072
rect 14185 6069 14197 6072
rect 14231 6069 14243 6103
rect 14292 6100 14320 6140
rect 15105 6103 15163 6109
rect 15105 6100 15117 6103
rect 14292 6072 15117 6100
rect 14185 6063 14243 6069
rect 15105 6069 15117 6072
rect 15151 6069 15163 6103
rect 15105 6063 15163 6069
rect 16390 6060 16396 6112
rect 16448 6100 16454 6112
rect 17420 6109 17448 6208
rect 19334 6196 19340 6208
rect 19392 6196 19398 6248
rect 18230 6128 18236 6180
rect 18288 6168 18294 6180
rect 19245 6171 19303 6177
rect 19245 6168 19257 6171
rect 18288 6140 19257 6168
rect 18288 6128 18294 6140
rect 19245 6137 19257 6140
rect 19291 6137 19303 6171
rect 19245 6131 19303 6137
rect 19702 6128 19708 6180
rect 19760 6168 19766 6180
rect 19886 6168 19892 6180
rect 19760 6140 19892 6168
rect 19760 6128 19766 6140
rect 19886 6128 19892 6140
rect 19944 6128 19950 6180
rect 17405 6103 17463 6109
rect 17405 6100 17417 6103
rect 16448 6072 17417 6100
rect 16448 6060 16454 6072
rect 17405 6069 17417 6072
rect 17451 6069 17463 6103
rect 17405 6063 17463 6069
rect 17586 6060 17592 6112
rect 17644 6100 17650 6112
rect 17957 6103 18015 6109
rect 17957 6100 17969 6103
rect 17644 6072 17969 6100
rect 17644 6060 17650 6072
rect 17957 6069 17969 6072
rect 18003 6069 18015 6103
rect 18598 6100 18604 6112
rect 18559 6072 18604 6100
rect 17957 6063 18015 6069
rect 18598 6060 18604 6072
rect 18656 6060 18662 6112
rect 20806 6060 20812 6112
rect 20864 6100 20870 6112
rect 21269 6103 21327 6109
rect 21269 6100 21281 6103
rect 20864 6072 21281 6100
rect 20864 6060 20870 6072
rect 21269 6069 21281 6072
rect 21315 6069 21327 6103
rect 21269 6063 21327 6069
rect 22094 6060 22100 6112
rect 22152 6100 22158 6112
rect 23492 6109 23520 6276
rect 24762 6264 24768 6276
rect 24820 6264 24826 6316
rect 24670 6168 24676 6180
rect 24136 6140 24676 6168
rect 24136 6109 24164 6140
rect 24670 6128 24676 6140
rect 24728 6128 24734 6180
rect 27890 6168 27896 6180
rect 25700 6140 27896 6168
rect 23477 6103 23535 6109
rect 23477 6100 23489 6103
rect 22152 6072 23489 6100
rect 22152 6060 22158 6072
rect 23477 6069 23489 6072
rect 23523 6069 23535 6103
rect 23477 6063 23535 6069
rect 24121 6103 24179 6109
rect 24121 6069 24133 6103
rect 24167 6069 24179 6103
rect 24121 6063 24179 6069
rect 24302 6060 24308 6112
rect 24360 6100 24366 6112
rect 25700 6100 25728 6140
rect 27890 6128 27896 6140
rect 27948 6128 27954 6180
rect 24360 6072 25728 6100
rect 24360 6060 24366 6072
rect 25958 6060 25964 6112
rect 26016 6100 26022 6112
rect 26145 6103 26203 6109
rect 26145 6100 26157 6103
rect 26016 6072 26157 6100
rect 26016 6060 26022 6072
rect 26145 6069 26157 6072
rect 26191 6069 26203 6103
rect 26145 6063 26203 6069
rect 27157 6103 27215 6109
rect 27157 6069 27169 6103
rect 27203 6100 27215 6103
rect 27430 6100 27436 6112
rect 27203 6072 27436 6100
rect 27203 6069 27215 6072
rect 27157 6063 27215 6069
rect 27430 6060 27436 6072
rect 27488 6060 27494 6112
rect 1104 6010 28060 6032
rect 1104 5958 5442 6010
rect 5494 5958 5506 6010
rect 5558 5958 5570 6010
rect 5622 5958 5634 6010
rect 5686 5958 5698 6010
rect 5750 5958 14428 6010
rect 14480 5958 14492 6010
rect 14544 5958 14556 6010
rect 14608 5958 14620 6010
rect 14672 5958 14684 6010
rect 14736 5958 23413 6010
rect 23465 5958 23477 6010
rect 23529 5958 23541 6010
rect 23593 5958 23605 6010
rect 23657 5958 23669 6010
rect 23721 5958 28060 6010
rect 1104 5936 28060 5958
rect 1946 5856 1952 5908
rect 2004 5896 2010 5908
rect 2685 5899 2743 5905
rect 2685 5896 2697 5899
rect 2004 5868 2697 5896
rect 2004 5856 2010 5868
rect 2685 5865 2697 5868
rect 2731 5865 2743 5899
rect 2685 5859 2743 5865
rect 3145 5899 3203 5905
rect 3145 5865 3157 5899
rect 3191 5896 3203 5899
rect 4246 5896 4252 5908
rect 3191 5868 4252 5896
rect 3191 5865 3203 5868
rect 3145 5859 3203 5865
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 5074 5896 5080 5908
rect 5035 5868 5080 5896
rect 5074 5856 5080 5868
rect 5132 5856 5138 5908
rect 5902 5856 5908 5908
rect 5960 5896 5966 5908
rect 12986 5896 12992 5908
rect 5960 5868 12992 5896
rect 5960 5856 5966 5868
rect 12986 5856 12992 5868
rect 13044 5856 13050 5908
rect 13449 5899 13507 5905
rect 13449 5865 13461 5899
rect 13495 5896 13507 5899
rect 13722 5896 13728 5908
rect 13495 5868 13728 5896
rect 13495 5865 13507 5868
rect 13449 5859 13507 5865
rect 13722 5856 13728 5868
rect 13780 5856 13786 5908
rect 20806 5896 20812 5908
rect 14108 5868 18828 5896
rect 20767 5868 20812 5896
rect 1397 5831 1455 5837
rect 1397 5797 1409 5831
rect 1443 5828 1455 5831
rect 2866 5828 2872 5840
rect 1443 5800 2872 5828
rect 1443 5797 1455 5800
rect 1397 5791 1455 5797
rect 2866 5788 2872 5800
rect 2924 5788 2930 5840
rect 2958 5788 2964 5840
rect 3016 5788 3022 5840
rect 4062 5788 4068 5840
rect 4120 5788 4126 5840
rect 4264 5828 4292 5856
rect 5537 5831 5595 5837
rect 5537 5828 5549 5831
rect 4264 5800 5549 5828
rect 5537 5797 5549 5800
rect 5583 5797 5595 5831
rect 5537 5791 5595 5797
rect 7282 5788 7288 5840
rect 7340 5828 7346 5840
rect 10226 5828 10232 5840
rect 7340 5800 10232 5828
rect 7340 5788 7346 5800
rect 10226 5788 10232 5800
rect 10284 5788 10290 5840
rect 12710 5788 12716 5840
rect 12768 5828 12774 5840
rect 12768 5800 13124 5828
rect 12768 5788 12774 5800
rect 2976 5760 3004 5788
rect 2884 5732 3004 5760
rect 1581 5695 1639 5701
rect 1581 5661 1593 5695
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5692 2283 5695
rect 2774 5692 2780 5704
rect 2271 5664 2780 5692
rect 2271 5661 2283 5664
rect 2225 5655 2283 5661
rect 1596 5624 1624 5655
rect 2774 5652 2780 5664
rect 2832 5652 2838 5704
rect 2884 5701 2912 5732
rect 3050 5720 3056 5772
rect 3108 5720 3114 5772
rect 3789 5763 3847 5769
rect 3789 5729 3801 5763
rect 3835 5760 3847 5763
rect 4080 5760 4108 5788
rect 3835 5732 4108 5760
rect 3835 5729 3847 5732
rect 3789 5723 3847 5729
rect 4890 5720 4896 5772
rect 4948 5760 4954 5772
rect 4948 5732 5672 5760
rect 4948 5720 4954 5732
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5692 3019 5695
rect 3068 5692 3096 5720
rect 3234 5692 3240 5704
rect 3007 5664 3096 5692
rect 3195 5664 3240 5692
rect 3007 5661 3019 5664
rect 2961 5655 3019 5661
rect 3234 5652 3240 5664
rect 3292 5652 3298 5704
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5692 4123 5695
rect 4246 5692 4252 5704
rect 4111 5664 4252 5692
rect 4111 5661 4123 5664
rect 4065 5655 4123 5661
rect 4246 5652 4252 5664
rect 4304 5692 4310 5704
rect 5258 5692 5264 5704
rect 4304 5664 5264 5692
rect 4304 5652 4310 5664
rect 5258 5652 5264 5664
rect 5316 5652 5322 5704
rect 5350 5652 5356 5704
rect 5408 5692 5414 5704
rect 5644 5701 5672 5732
rect 8478 5720 8484 5772
rect 8536 5760 8542 5772
rect 9398 5760 9404 5772
rect 8536 5732 9168 5760
rect 9359 5732 9404 5760
rect 8536 5720 8542 5732
rect 9140 5701 9168 5732
rect 9398 5720 9404 5732
rect 9456 5720 9462 5772
rect 10410 5720 10416 5772
rect 10468 5760 10474 5772
rect 10505 5763 10563 5769
rect 10505 5760 10517 5763
rect 10468 5732 10517 5760
rect 10468 5720 10474 5732
rect 10505 5729 10517 5732
rect 10551 5729 10563 5763
rect 10505 5723 10563 5729
rect 13096 5760 13124 5800
rect 13538 5788 13544 5840
rect 13596 5828 13602 5840
rect 14108 5828 14136 5868
rect 13596 5800 14136 5828
rect 13596 5788 13602 5800
rect 14182 5788 14188 5840
rect 14240 5828 14246 5840
rect 14737 5831 14795 5837
rect 14737 5828 14749 5831
rect 14240 5800 14749 5828
rect 14240 5788 14246 5800
rect 14737 5797 14749 5800
rect 14783 5797 14795 5831
rect 15654 5828 15660 5840
rect 15615 5800 15660 5828
rect 14737 5791 14795 5797
rect 15654 5788 15660 5800
rect 15712 5828 15718 5840
rect 16390 5828 16396 5840
rect 15712 5800 16396 5828
rect 15712 5788 15718 5800
rect 16390 5788 16396 5800
rect 16448 5828 16454 5840
rect 16669 5831 16727 5837
rect 16669 5828 16681 5831
rect 16448 5800 16681 5828
rect 16448 5788 16454 5800
rect 16669 5797 16681 5800
rect 16715 5797 16727 5831
rect 18800 5828 18828 5868
rect 20806 5856 20812 5868
rect 20864 5856 20870 5908
rect 20990 5896 20996 5908
rect 20951 5868 20996 5896
rect 20990 5856 20996 5868
rect 21048 5856 21054 5908
rect 21284 5868 21588 5896
rect 21284 5828 21312 5868
rect 18800 5800 21312 5828
rect 21453 5831 21511 5837
rect 16669 5791 16727 5797
rect 21453 5797 21465 5831
rect 21499 5797 21511 5831
rect 21560 5828 21588 5868
rect 21910 5856 21916 5908
rect 21968 5896 21974 5908
rect 22281 5899 22339 5905
rect 22281 5896 22293 5899
rect 21968 5868 22293 5896
rect 21968 5856 21974 5868
rect 22281 5865 22293 5868
rect 22327 5865 22339 5899
rect 22462 5896 22468 5908
rect 22423 5868 22468 5896
rect 22281 5859 22339 5865
rect 22462 5856 22468 5868
rect 22520 5856 22526 5908
rect 23014 5856 23020 5908
rect 23072 5896 23078 5908
rect 24581 5899 24639 5905
rect 23072 5868 24440 5896
rect 23072 5856 23078 5868
rect 23842 5828 23848 5840
rect 21560 5800 22094 5828
rect 21453 5791 21511 5797
rect 14826 5760 14832 5772
rect 13096 5732 14832 5760
rect 5629 5695 5687 5701
rect 5408 5664 5453 5692
rect 5408 5652 5414 5664
rect 5629 5661 5641 5695
rect 5675 5661 5687 5695
rect 5629 5655 5687 5661
rect 7837 5695 7895 5701
rect 7837 5661 7849 5695
rect 7883 5692 7895 5695
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 7883 5664 8953 5692
rect 7883 5661 7895 5664
rect 7837 5655 7895 5661
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 9125 5695 9183 5701
rect 9125 5661 9137 5695
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 9214 5652 9220 5704
rect 9272 5692 9278 5704
rect 9493 5695 9551 5701
rect 9272 5664 9317 5692
rect 9272 5652 9278 5664
rect 9493 5661 9505 5695
rect 9539 5692 9551 5695
rect 10772 5695 10830 5701
rect 9539 5664 9628 5692
rect 9539 5661 9551 5664
rect 9493 5655 9551 5661
rect 3050 5624 3056 5636
rect 1596 5596 3056 5624
rect 3050 5584 3056 5596
rect 3108 5584 3114 5636
rect 6638 5624 6644 5636
rect 6599 5596 6644 5624
rect 6638 5584 6644 5596
rect 6696 5584 6702 5636
rect 6825 5627 6883 5633
rect 6825 5593 6837 5627
rect 6871 5624 6883 5627
rect 8021 5627 8079 5633
rect 8021 5624 8033 5627
rect 6871 5596 8033 5624
rect 6871 5593 6883 5596
rect 6825 5587 6883 5593
rect 8021 5593 8033 5596
rect 8067 5624 8079 5627
rect 8478 5624 8484 5636
rect 8067 5596 8484 5624
rect 8067 5593 8079 5596
rect 8021 5587 8079 5593
rect 8478 5584 8484 5596
rect 8536 5624 8542 5636
rect 9600 5624 9628 5664
rect 10772 5661 10784 5695
rect 10818 5692 10830 5695
rect 11330 5692 11336 5704
rect 10818 5664 11336 5692
rect 10818 5661 10830 5664
rect 10772 5655 10830 5661
rect 11330 5652 11336 5664
rect 11388 5652 11394 5704
rect 12529 5695 12587 5701
rect 12529 5661 12541 5695
rect 12575 5692 12587 5695
rect 12710 5692 12716 5704
rect 12575 5664 12716 5692
rect 12575 5661 12587 5664
rect 12529 5655 12587 5661
rect 12710 5652 12716 5664
rect 12768 5652 12774 5704
rect 13096 5692 13124 5732
rect 14826 5720 14832 5732
rect 14884 5760 14890 5772
rect 17310 5760 17316 5772
rect 14884 5732 16436 5760
rect 17271 5732 17316 5760
rect 14884 5720 14890 5732
rect 13156 5695 13214 5701
rect 13156 5692 13168 5695
rect 13096 5664 13168 5692
rect 13156 5661 13168 5664
rect 13202 5661 13214 5695
rect 13156 5655 13214 5661
rect 13265 5695 13323 5701
rect 13265 5661 13277 5695
rect 13311 5661 13323 5695
rect 13538 5692 13544 5704
rect 13499 5664 13544 5692
rect 13265 5655 13323 5661
rect 9674 5624 9680 5636
rect 8536 5596 9536 5624
rect 9600 5596 9680 5624
rect 8536 5584 8542 5596
rect 9508 5568 9536 5596
rect 9674 5584 9680 5596
rect 9732 5584 9738 5636
rect 2041 5559 2099 5565
rect 2041 5525 2053 5559
rect 2087 5556 2099 5559
rect 3418 5556 3424 5568
rect 2087 5528 3424 5556
rect 2087 5525 2099 5528
rect 2041 5519 2099 5525
rect 3418 5516 3424 5528
rect 3476 5516 3482 5568
rect 4798 5516 4804 5568
rect 4856 5556 4862 5568
rect 7009 5559 7067 5565
rect 7009 5556 7021 5559
rect 4856 5528 7021 5556
rect 4856 5516 4862 5528
rect 7009 5525 7021 5528
rect 7055 5525 7067 5559
rect 7009 5519 7067 5525
rect 7282 5516 7288 5568
rect 7340 5556 7346 5568
rect 8205 5559 8263 5565
rect 8205 5556 8217 5559
rect 7340 5528 8217 5556
rect 7340 5516 7346 5528
rect 8205 5525 8217 5528
rect 8251 5525 8263 5559
rect 8205 5519 8263 5525
rect 8754 5516 8760 5568
rect 8812 5556 8818 5568
rect 9398 5556 9404 5568
rect 8812 5528 9404 5556
rect 8812 5516 8818 5528
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 9490 5516 9496 5568
rect 9548 5516 9554 5568
rect 11882 5556 11888 5568
rect 11843 5528 11888 5556
rect 11882 5516 11888 5528
rect 11940 5516 11946 5568
rect 12345 5559 12403 5565
rect 12345 5525 12357 5559
rect 12391 5556 12403 5559
rect 12802 5556 12808 5568
rect 12391 5528 12808 5556
rect 12391 5525 12403 5528
rect 12345 5519 12403 5525
rect 12802 5516 12808 5528
rect 12860 5516 12866 5568
rect 12986 5556 12992 5568
rect 12947 5528 12992 5556
rect 12986 5516 12992 5528
rect 13044 5516 13050 5568
rect 13280 5556 13308 5655
rect 13538 5652 13544 5664
rect 13596 5652 13602 5704
rect 15396 5701 15424 5732
rect 14369 5695 14427 5701
rect 14369 5661 14381 5695
rect 14415 5692 14427 5695
rect 15197 5695 15255 5701
rect 15197 5692 15209 5695
rect 14415 5664 15209 5692
rect 14415 5661 14427 5664
rect 14369 5655 14427 5661
rect 15197 5661 15209 5664
rect 15243 5661 15255 5695
rect 15197 5655 15255 5661
rect 15381 5695 15439 5701
rect 15381 5661 15393 5695
rect 15427 5661 15439 5695
rect 15381 5655 15439 5661
rect 15473 5695 15531 5701
rect 15473 5661 15485 5695
rect 15519 5661 15531 5695
rect 15746 5692 15752 5704
rect 15707 5664 15752 5692
rect 15473 5655 15531 5661
rect 13906 5584 13912 5636
rect 13964 5624 13970 5636
rect 14553 5627 14611 5633
rect 14553 5624 14565 5627
rect 13964 5596 14565 5624
rect 13964 5584 13970 5596
rect 14553 5593 14565 5596
rect 14599 5624 14611 5627
rect 15102 5624 15108 5636
rect 14599 5596 15108 5624
rect 14599 5593 14611 5596
rect 14553 5587 14611 5593
rect 15102 5584 15108 5596
rect 15160 5584 15166 5636
rect 15286 5584 15292 5636
rect 15344 5624 15350 5636
rect 15488 5624 15516 5655
rect 15746 5652 15752 5664
rect 15804 5652 15810 5704
rect 16408 5701 16436 5732
rect 17310 5720 17316 5732
rect 17368 5720 17374 5772
rect 19610 5720 19616 5772
rect 19668 5760 19674 5772
rect 21468 5760 21496 5791
rect 19668 5732 21496 5760
rect 19668 5720 19674 5732
rect 16393 5695 16451 5701
rect 16393 5661 16405 5695
rect 16439 5661 16451 5695
rect 16393 5655 16451 5661
rect 16485 5695 16543 5701
rect 16485 5661 16497 5695
rect 16531 5661 16543 5695
rect 16758 5692 16764 5704
rect 16719 5664 16764 5692
rect 16485 5655 16543 5661
rect 15344 5596 15516 5624
rect 16500 5624 16528 5655
rect 16758 5652 16764 5664
rect 16816 5652 16822 5704
rect 17034 5652 17040 5704
rect 17092 5692 17098 5704
rect 17569 5695 17627 5701
rect 17569 5692 17581 5695
rect 17092 5664 17581 5692
rect 17092 5652 17098 5664
rect 17569 5661 17581 5664
rect 17615 5661 17627 5695
rect 17569 5655 17627 5661
rect 19334 5652 19340 5704
rect 19392 5692 19398 5704
rect 19429 5695 19487 5701
rect 19429 5692 19441 5695
rect 19392 5664 19441 5692
rect 19392 5652 19398 5664
rect 19429 5661 19441 5664
rect 19475 5661 19487 5695
rect 20070 5692 20076 5704
rect 20031 5664 20076 5692
rect 19429 5655 19487 5661
rect 20070 5652 20076 5664
rect 20128 5652 20134 5704
rect 20180 5664 20852 5692
rect 20180 5624 20208 5664
rect 16500 5596 20208 5624
rect 20625 5627 20683 5633
rect 15344 5584 15350 5596
rect 15654 5556 15660 5568
rect 13280 5528 15660 5556
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 16206 5556 16212 5568
rect 16167 5528 16212 5556
rect 16206 5516 16212 5528
rect 16264 5516 16270 5568
rect 16758 5516 16764 5568
rect 16816 5556 16822 5568
rect 17586 5556 17592 5568
rect 16816 5528 17592 5556
rect 16816 5516 16822 5528
rect 17586 5516 17592 5528
rect 17644 5516 17650 5568
rect 18708 5565 18736 5596
rect 20625 5593 20637 5627
rect 20671 5624 20683 5627
rect 20714 5624 20720 5636
rect 20671 5596 20720 5624
rect 20671 5593 20683 5596
rect 20625 5587 20683 5593
rect 20714 5584 20720 5596
rect 20772 5584 20778 5636
rect 20824 5624 20852 5664
rect 21174 5652 21180 5704
rect 21232 5692 21238 5704
rect 21637 5695 21695 5701
rect 21637 5692 21649 5695
rect 21232 5664 21649 5692
rect 21232 5652 21238 5664
rect 21637 5661 21649 5664
rect 21683 5661 21695 5695
rect 22066 5692 22094 5800
rect 22756 5800 23848 5828
rect 22278 5720 22284 5772
rect 22336 5760 22342 5772
rect 22756 5760 22784 5800
rect 23842 5788 23848 5800
rect 23900 5788 23906 5840
rect 22336 5732 22784 5760
rect 22336 5720 22342 5732
rect 22830 5720 22836 5772
rect 22888 5760 22894 5772
rect 24412 5760 24440 5868
rect 24581 5865 24593 5899
rect 24627 5896 24639 5899
rect 24670 5896 24676 5908
rect 24627 5868 24676 5896
rect 24627 5865 24639 5868
rect 24581 5859 24639 5865
rect 24670 5856 24676 5868
rect 24728 5856 24734 5908
rect 24486 5788 24492 5840
rect 24544 5828 24550 5840
rect 25409 5831 25467 5837
rect 25409 5828 25421 5831
rect 24544 5800 25421 5828
rect 24544 5788 24550 5800
rect 25409 5797 25421 5800
rect 25455 5797 25467 5831
rect 25409 5791 25467 5797
rect 22888 5732 23612 5760
rect 24412 5732 24716 5760
rect 22888 5720 22894 5732
rect 23106 5692 23112 5704
rect 22066 5664 22324 5692
rect 23067 5664 23112 5692
rect 21637 5655 21695 5661
rect 21818 5624 21824 5636
rect 20824 5596 21824 5624
rect 21818 5584 21824 5596
rect 21876 5584 21882 5636
rect 22094 5624 22100 5636
rect 22055 5596 22100 5624
rect 22094 5584 22100 5596
rect 22152 5584 22158 5636
rect 22296 5624 22324 5664
rect 23106 5652 23112 5664
rect 23164 5652 23170 5704
rect 23584 5701 23612 5732
rect 23569 5695 23627 5701
rect 23569 5661 23581 5695
rect 23615 5661 23627 5695
rect 23569 5655 23627 5661
rect 23750 5652 23756 5704
rect 23808 5692 23814 5704
rect 23808 5664 24440 5692
rect 23808 5652 23814 5664
rect 24302 5624 24308 5636
rect 22296 5596 24308 5624
rect 24302 5584 24308 5596
rect 24360 5584 24366 5636
rect 24412 5633 24440 5664
rect 24578 5652 24584 5704
rect 24636 5652 24642 5704
rect 24688 5692 24716 5732
rect 24762 5720 24768 5772
rect 24820 5760 24826 5772
rect 25498 5760 25504 5772
rect 24820 5732 25504 5760
rect 24820 5720 24826 5732
rect 25498 5720 25504 5732
rect 25556 5760 25562 5772
rect 25961 5763 26019 5769
rect 25961 5760 25973 5763
rect 25556 5732 25973 5760
rect 25556 5720 25562 5732
rect 25961 5729 25973 5732
rect 26007 5729 26019 5763
rect 25961 5723 26019 5729
rect 25225 5695 25283 5701
rect 24688 5664 25176 5692
rect 24397 5627 24455 5633
rect 24397 5593 24409 5627
rect 24443 5593 24455 5627
rect 24596 5624 24624 5652
rect 25148 5624 25176 5664
rect 25225 5661 25237 5695
rect 25271 5692 25283 5695
rect 25682 5692 25688 5704
rect 25271 5664 25688 5692
rect 25271 5661 25283 5664
rect 25225 5655 25283 5661
rect 25682 5652 25688 5664
rect 25740 5652 25746 5704
rect 26228 5695 26286 5701
rect 26228 5661 26240 5695
rect 26274 5692 26286 5695
rect 27706 5692 27712 5704
rect 26274 5664 27712 5692
rect 26274 5661 26286 5664
rect 26228 5655 26286 5661
rect 27706 5652 27712 5664
rect 27764 5652 27770 5704
rect 28166 5624 28172 5636
rect 24596 5596 24808 5624
rect 25148 5596 28172 5624
rect 24397 5587 24455 5593
rect 18693 5559 18751 5565
rect 18693 5525 18705 5559
rect 18739 5525 18751 5559
rect 19242 5556 19248 5568
rect 19203 5528 19248 5556
rect 18693 5519 18751 5525
rect 19242 5516 19248 5528
rect 19300 5516 19306 5568
rect 19886 5556 19892 5568
rect 19847 5528 19892 5556
rect 19886 5516 19892 5528
rect 19944 5516 19950 5568
rect 20530 5516 20536 5568
rect 20588 5556 20594 5568
rect 20825 5559 20883 5565
rect 20825 5556 20837 5559
rect 20588 5528 20837 5556
rect 20588 5516 20594 5528
rect 20825 5525 20837 5528
rect 20871 5556 20883 5559
rect 22297 5559 22355 5565
rect 22297 5556 22309 5559
rect 20871 5528 22309 5556
rect 20871 5525 20883 5528
rect 20825 5519 20883 5525
rect 22297 5525 22309 5528
rect 22343 5525 22355 5559
rect 22297 5519 22355 5525
rect 22646 5516 22652 5568
rect 22704 5556 22710 5568
rect 22925 5559 22983 5565
rect 22925 5556 22937 5559
rect 22704 5528 22937 5556
rect 22704 5516 22710 5528
rect 22925 5525 22937 5528
rect 22971 5525 22983 5559
rect 22925 5519 22983 5525
rect 23753 5559 23811 5565
rect 23753 5525 23765 5559
rect 23799 5556 23811 5559
rect 23842 5556 23848 5568
rect 23799 5528 23848 5556
rect 23799 5525 23811 5528
rect 23753 5519 23811 5525
rect 23842 5516 23848 5528
rect 23900 5516 23906 5568
rect 24210 5516 24216 5568
rect 24268 5556 24274 5568
rect 24578 5556 24584 5568
rect 24636 5565 24642 5568
rect 24780 5565 24808 5596
rect 28166 5584 28172 5596
rect 28224 5584 28230 5636
rect 24636 5559 24655 5565
rect 24268 5528 24584 5556
rect 24268 5516 24274 5528
rect 24578 5516 24584 5528
rect 24643 5525 24655 5559
rect 24636 5519 24655 5525
rect 24765 5559 24823 5565
rect 24765 5525 24777 5559
rect 24811 5525 24823 5559
rect 24765 5519 24823 5525
rect 24636 5516 24642 5519
rect 26878 5516 26884 5568
rect 26936 5556 26942 5568
rect 27338 5556 27344 5568
rect 26936 5528 27344 5556
rect 26936 5516 26942 5528
rect 27338 5516 27344 5528
rect 27396 5516 27402 5568
rect 1104 5466 28060 5488
rect 1104 5414 9935 5466
rect 9987 5414 9999 5466
rect 10051 5414 10063 5466
rect 10115 5414 10127 5466
rect 10179 5414 10191 5466
rect 10243 5414 18920 5466
rect 18972 5414 18984 5466
rect 19036 5414 19048 5466
rect 19100 5414 19112 5466
rect 19164 5414 19176 5466
rect 19228 5414 28060 5466
rect 1104 5392 28060 5414
rect 3050 5352 3056 5364
rect 3011 5324 3056 5352
rect 3050 5312 3056 5324
rect 3108 5312 3114 5364
rect 3878 5312 3884 5364
rect 3936 5352 3942 5364
rect 6638 5352 6644 5364
rect 3936 5324 4384 5352
rect 6599 5324 6644 5352
rect 3936 5312 3942 5324
rect 2685 5287 2743 5293
rect 2685 5253 2697 5287
rect 2731 5284 2743 5287
rect 3789 5287 3847 5293
rect 3789 5284 3801 5287
rect 2731 5256 3801 5284
rect 2731 5253 2743 5256
rect 2685 5247 2743 5253
rect 3789 5253 3801 5256
rect 3835 5253 3847 5287
rect 4246 5284 4252 5296
rect 3789 5247 3847 5253
rect 3988 5256 4252 5284
rect 1857 5219 1915 5225
rect 1857 5185 1869 5219
rect 1903 5185 1915 5219
rect 1857 5179 1915 5185
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5216 2099 5219
rect 2869 5219 2927 5225
rect 2869 5216 2881 5219
rect 2087 5188 2881 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 2869 5185 2881 5188
rect 2915 5216 2927 5219
rect 3602 5216 3608 5228
rect 2915 5188 3608 5216
rect 2915 5185 2927 5188
rect 2869 5179 2927 5185
rect 1872 5148 1900 5179
rect 3602 5176 3608 5188
rect 3660 5216 3666 5228
rect 3988 5225 4016 5256
rect 4246 5244 4252 5256
rect 4304 5244 4310 5296
rect 3973 5219 4031 5225
rect 3660 5188 3924 5216
rect 3660 5176 3666 5188
rect 3786 5148 3792 5160
rect 1872 5120 3792 5148
rect 3786 5108 3792 5120
rect 3844 5108 3850 5160
rect 3896 5148 3924 5188
rect 3973 5185 3985 5219
rect 4019 5185 4031 5219
rect 3973 5179 4031 5185
rect 4062 5176 4068 5228
rect 4120 5216 4126 5228
rect 4356 5225 4384 5324
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 7006 5312 7012 5364
rect 7064 5312 7070 5364
rect 7558 5312 7564 5364
rect 7616 5352 7622 5364
rect 8754 5352 8760 5364
rect 7616 5324 8760 5352
rect 7616 5312 7622 5324
rect 8754 5312 8760 5324
rect 8812 5312 8818 5364
rect 9214 5352 9220 5364
rect 9175 5324 9220 5352
rect 9214 5312 9220 5324
rect 9272 5312 9278 5364
rect 9858 5312 9864 5364
rect 9916 5352 9922 5364
rect 9953 5355 10011 5361
rect 9953 5352 9965 5355
rect 9916 5324 9965 5352
rect 9916 5312 9922 5324
rect 9953 5321 9965 5324
rect 9999 5321 10011 5355
rect 11054 5352 11060 5364
rect 9953 5315 10011 5321
rect 10152 5324 11060 5352
rect 4985 5287 5043 5293
rect 4985 5253 4997 5287
rect 5031 5284 5043 5287
rect 6454 5284 6460 5296
rect 5031 5256 6460 5284
rect 5031 5253 5043 5256
rect 4985 5247 5043 5253
rect 6454 5244 6460 5256
rect 6512 5244 6518 5296
rect 7024 5284 7052 5312
rect 7282 5284 7288 5296
rect 7024 5256 7288 5284
rect 4341 5219 4399 5225
rect 4120 5188 4165 5216
rect 4120 5176 4126 5188
rect 4341 5185 4353 5219
rect 4387 5185 4399 5219
rect 4341 5179 4399 5185
rect 5169 5219 5227 5225
rect 5169 5185 5181 5219
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 5184 5148 5212 5179
rect 5258 5176 5264 5228
rect 5316 5216 5322 5228
rect 6638 5216 6644 5228
rect 5316 5188 6644 5216
rect 5316 5176 5322 5188
rect 6638 5176 6644 5188
rect 6696 5216 6702 5228
rect 6825 5219 6883 5225
rect 6825 5216 6837 5219
rect 6696 5188 6837 5216
rect 6696 5176 6702 5188
rect 6825 5185 6837 5188
rect 6871 5185 6883 5219
rect 6825 5179 6883 5185
rect 6917 5219 6975 5225
rect 6917 5185 6929 5219
rect 6963 5216 6975 5219
rect 7024 5216 7052 5256
rect 7282 5244 7288 5256
rect 7340 5244 7346 5296
rect 7190 5216 7196 5228
rect 6963 5188 7052 5216
rect 7151 5188 7196 5216
rect 6963 5185 6975 5188
rect 6917 5179 6975 5185
rect 7190 5176 7196 5188
rect 7248 5176 7254 5228
rect 7558 5176 7564 5228
rect 7616 5216 7622 5228
rect 10152 5225 10180 5324
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 12802 5312 12808 5364
rect 12860 5352 12866 5364
rect 15654 5352 15660 5364
rect 12860 5324 13584 5352
rect 15615 5324 15660 5352
rect 12860 5312 12866 5324
rect 11517 5287 11575 5293
rect 11517 5284 11529 5287
rect 10244 5256 11529 5284
rect 10244 5225 10272 5256
rect 11517 5253 11529 5256
rect 11563 5284 11575 5287
rect 11882 5284 11888 5296
rect 11563 5256 11888 5284
rect 11563 5253 11575 5256
rect 11517 5247 11575 5253
rect 11882 5244 11888 5256
rect 11940 5244 11946 5296
rect 12434 5244 12440 5296
rect 12492 5284 12498 5296
rect 12492 5256 12537 5284
rect 12492 5244 12498 5256
rect 12986 5244 12992 5296
rect 13044 5284 13050 5296
rect 13449 5287 13507 5293
rect 13449 5284 13461 5287
rect 13044 5256 13461 5284
rect 13044 5244 13050 5256
rect 13449 5253 13461 5256
rect 13495 5253 13507 5287
rect 13556 5284 13584 5324
rect 15654 5312 15660 5324
rect 15712 5312 15718 5364
rect 20622 5352 20628 5364
rect 20583 5324 20628 5352
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 20806 5312 20812 5364
rect 20864 5352 20870 5364
rect 21910 5352 21916 5364
rect 20864 5324 21916 5352
rect 20864 5312 20870 5324
rect 21910 5312 21916 5324
rect 21968 5312 21974 5364
rect 23474 5312 23480 5364
rect 23532 5352 23538 5364
rect 23937 5355 23995 5361
rect 23937 5352 23949 5355
rect 23532 5324 23949 5352
rect 23532 5312 23538 5324
rect 23937 5321 23949 5324
rect 23983 5321 23995 5355
rect 23937 5315 23995 5321
rect 24765 5355 24823 5361
rect 24765 5321 24777 5355
rect 24811 5321 24823 5355
rect 24765 5315 24823 5321
rect 14522 5287 14580 5293
rect 14522 5284 14534 5287
rect 13556 5256 14534 5284
rect 13449 5247 13507 5253
rect 14522 5253 14534 5256
rect 14568 5253 14580 5287
rect 17310 5284 17316 5296
rect 14522 5247 14580 5253
rect 16684 5256 17316 5284
rect 8093 5219 8151 5225
rect 8093 5216 8105 5219
rect 7616 5188 8105 5216
rect 7616 5176 7622 5188
rect 8093 5185 8105 5188
rect 8139 5185 8151 5219
rect 8093 5179 8151 5185
rect 10137 5219 10195 5225
rect 10137 5185 10149 5219
rect 10183 5185 10195 5219
rect 10137 5179 10195 5185
rect 10229 5219 10287 5225
rect 10229 5185 10241 5219
rect 10275 5185 10287 5219
rect 10502 5216 10508 5228
rect 10463 5188 10508 5216
rect 10229 5179 10287 5185
rect 10502 5176 10508 5188
rect 10560 5176 10566 5228
rect 11422 5176 11428 5228
rect 11480 5216 11486 5228
rect 11793 5219 11851 5225
rect 11793 5216 11805 5219
rect 11480 5188 11805 5216
rect 11480 5176 11486 5188
rect 11793 5185 11805 5188
rect 11839 5185 11851 5219
rect 11793 5179 11851 5185
rect 12250 5176 12256 5228
rect 12308 5216 12314 5228
rect 12621 5219 12679 5225
rect 12621 5216 12633 5219
rect 12308 5188 12633 5216
rect 12308 5176 12314 5188
rect 12621 5185 12633 5188
rect 12667 5185 12679 5219
rect 12621 5179 12679 5185
rect 12805 5219 12863 5225
rect 12805 5185 12817 5219
rect 12851 5216 12863 5219
rect 12894 5216 12900 5228
rect 12851 5188 12900 5216
rect 12851 5185 12863 5188
rect 12805 5179 12863 5185
rect 3896 5120 5212 5148
rect 7006 5108 7012 5160
rect 7064 5148 7070 5160
rect 7834 5148 7840 5160
rect 7064 5120 7840 5148
rect 7064 5108 7070 5120
rect 7834 5108 7840 5120
rect 7892 5108 7898 5160
rect 11514 5108 11520 5160
rect 11572 5148 11578 5160
rect 11609 5151 11667 5157
rect 11609 5148 11621 5151
rect 11572 5120 11621 5148
rect 11572 5108 11578 5120
rect 11609 5117 11621 5120
rect 11655 5117 11667 5151
rect 12636 5148 12664 5179
rect 12894 5176 12900 5188
rect 12952 5176 12958 5228
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5216 13691 5219
rect 13906 5216 13912 5228
rect 13679 5188 13912 5216
rect 13679 5185 13691 5188
rect 13633 5179 13691 5185
rect 13648 5148 13676 5179
rect 13906 5176 13912 5188
rect 13964 5176 13970 5228
rect 14274 5216 14280 5228
rect 14235 5188 14280 5216
rect 14274 5176 14280 5188
rect 14332 5176 14338 5228
rect 16684 5225 16712 5256
rect 17310 5244 17316 5256
rect 17368 5244 17374 5296
rect 18046 5244 18052 5296
rect 18104 5284 18110 5296
rect 20257 5287 20315 5293
rect 18104 5256 19564 5284
rect 18104 5244 18110 5256
rect 16669 5219 16727 5225
rect 16669 5185 16681 5219
rect 16715 5185 16727 5219
rect 16925 5219 16983 5225
rect 16925 5216 16937 5219
rect 16669 5179 16727 5185
rect 16776 5188 16937 5216
rect 12636 5120 13676 5148
rect 11609 5111 11667 5117
rect 16298 5108 16304 5160
rect 16356 5148 16362 5160
rect 16776 5148 16804 5188
rect 16925 5185 16937 5188
rect 16971 5185 16983 5219
rect 18414 5216 18420 5228
rect 16925 5179 16983 5185
rect 18064 5188 18420 5216
rect 18064 5160 18092 5188
rect 18414 5176 18420 5188
rect 18472 5216 18478 5228
rect 19536 5225 19564 5256
rect 20257 5253 20269 5287
rect 20303 5284 20315 5287
rect 20346 5284 20352 5296
rect 20303 5256 20352 5284
rect 20303 5253 20315 5256
rect 20257 5247 20315 5253
rect 20346 5244 20352 5256
rect 20404 5244 20410 5296
rect 20530 5284 20536 5296
rect 20472 5253 20536 5284
rect 18785 5219 18843 5225
rect 18785 5216 18797 5219
rect 18472 5188 18797 5216
rect 18472 5176 18478 5188
rect 18785 5185 18797 5188
rect 18831 5185 18843 5219
rect 18785 5179 18843 5185
rect 19521 5219 19579 5225
rect 20472 5222 20499 5253
rect 19521 5185 19533 5219
rect 19567 5185 19579 5219
rect 20487 5219 20499 5222
rect 20533 5244 20536 5253
rect 20588 5244 20594 5296
rect 22189 5287 22247 5293
rect 22189 5253 22201 5287
rect 22235 5284 22247 5287
rect 22462 5284 22468 5296
rect 22235 5256 22468 5284
rect 22235 5253 22247 5256
rect 22189 5247 22247 5253
rect 22462 5244 22468 5256
rect 22520 5244 22526 5296
rect 22922 5284 22928 5296
rect 22848 5256 22928 5284
rect 20533 5219 20545 5244
rect 20487 5213 20545 5219
rect 21269 5219 21327 5225
rect 19521 5179 19579 5185
rect 21269 5185 21281 5219
rect 21315 5216 21327 5219
rect 21634 5216 21640 5228
rect 21315 5188 21640 5216
rect 21315 5185 21327 5188
rect 21269 5179 21327 5185
rect 16356 5120 16804 5148
rect 16356 5108 16362 5120
rect 18046 5108 18052 5160
rect 18104 5108 18110 5160
rect 4249 5083 4307 5089
rect 4249 5049 4261 5083
rect 4295 5080 4307 5083
rect 4338 5080 4344 5092
rect 4295 5052 4344 5080
rect 4295 5049 4307 5052
rect 4249 5043 4307 5049
rect 4338 5040 4344 5052
rect 4396 5040 4402 5092
rect 4890 5040 4896 5092
rect 4948 5080 4954 5092
rect 5258 5080 5264 5092
rect 4948 5052 5264 5080
rect 4948 5040 4954 5052
rect 5258 5040 5264 5052
rect 5316 5040 5322 5092
rect 7190 5040 7196 5092
rect 7248 5080 7254 5092
rect 7466 5080 7472 5092
rect 7248 5052 7472 5080
rect 7248 5040 7254 5052
rect 7466 5040 7472 5052
rect 7524 5040 7530 5092
rect 12710 5040 12716 5092
rect 12768 5080 12774 5092
rect 13817 5083 13875 5089
rect 13817 5080 13829 5083
rect 12768 5052 13829 5080
rect 12768 5040 12774 5052
rect 13817 5049 13829 5052
rect 13863 5049 13875 5083
rect 18800 5080 18828 5179
rect 20530 5108 20536 5160
rect 20588 5148 20594 5160
rect 21284 5148 21312 5179
rect 21634 5176 21640 5188
rect 21692 5176 21698 5228
rect 22051 5220 22109 5225
rect 22051 5219 22131 5220
rect 22051 5185 22063 5219
rect 22097 5216 22131 5219
rect 22281 5219 22339 5225
rect 22097 5188 22232 5216
rect 22097 5185 22109 5188
rect 22051 5179 22109 5185
rect 20588 5120 21312 5148
rect 22204 5148 22232 5188
rect 22281 5185 22293 5219
rect 22327 5216 22339 5219
rect 22554 5216 22560 5228
rect 22327 5188 22560 5216
rect 22327 5185 22339 5188
rect 22281 5179 22339 5185
rect 22554 5176 22560 5188
rect 22612 5176 22618 5228
rect 22848 5225 22876 5256
rect 22922 5244 22928 5256
rect 22980 5244 22986 5296
rect 23569 5287 23627 5293
rect 23569 5253 23581 5287
rect 23615 5284 23627 5287
rect 23658 5284 23664 5296
rect 23615 5256 23664 5284
rect 23615 5253 23627 5256
rect 23569 5247 23627 5253
rect 23658 5244 23664 5256
rect 23716 5244 23722 5296
rect 23785 5287 23843 5293
rect 23785 5253 23797 5287
rect 23831 5284 23843 5287
rect 24210 5284 24216 5296
rect 23831 5256 24216 5284
rect 23831 5253 23843 5256
rect 23785 5247 23843 5253
rect 24210 5244 24216 5256
rect 24268 5244 24274 5296
rect 24394 5284 24400 5296
rect 24355 5256 24400 5284
rect 24394 5244 24400 5256
rect 24452 5244 24458 5296
rect 24578 5244 24584 5296
rect 24636 5293 24642 5296
rect 24636 5287 24655 5293
rect 24643 5253 24655 5287
rect 24780 5284 24808 5315
rect 24854 5284 24860 5296
rect 24780 5256 24860 5284
rect 24636 5247 24655 5253
rect 24636 5244 24642 5247
rect 24854 5244 24860 5256
rect 24912 5244 24918 5296
rect 26970 5284 26976 5296
rect 26931 5256 26976 5284
rect 26970 5244 26976 5256
rect 27028 5244 27034 5296
rect 27173 5287 27231 5293
rect 27173 5284 27185 5287
rect 27080 5256 27185 5284
rect 22833 5219 22891 5225
rect 22833 5185 22845 5219
rect 22879 5185 22891 5219
rect 27080 5216 27108 5256
rect 27173 5253 27185 5256
rect 27219 5253 27231 5287
rect 27173 5247 27231 5253
rect 22833 5179 22891 5185
rect 22940 5188 27108 5216
rect 22738 5148 22744 5160
rect 22204 5120 22744 5148
rect 20588 5108 20594 5120
rect 22738 5108 22744 5120
rect 22796 5108 22802 5160
rect 22940 5080 22968 5188
rect 26988 5160 27016 5188
rect 23014 5108 23020 5160
rect 23072 5148 23078 5160
rect 25593 5151 25651 5157
rect 25593 5148 25605 5151
rect 23072 5120 25605 5148
rect 23072 5108 23078 5120
rect 25593 5117 25605 5120
rect 25639 5117 25651 5151
rect 25593 5111 25651 5117
rect 25682 5108 25688 5160
rect 25740 5148 25746 5160
rect 25869 5151 25927 5157
rect 25869 5148 25881 5151
rect 25740 5120 25881 5148
rect 25740 5108 25746 5120
rect 25869 5117 25881 5120
rect 25915 5148 25927 5151
rect 26878 5148 26884 5160
rect 25915 5120 26884 5148
rect 25915 5117 25927 5120
rect 25869 5111 25927 5117
rect 26878 5108 26884 5120
rect 26936 5108 26942 5160
rect 26970 5108 26976 5160
rect 27028 5108 27034 5160
rect 18800 5052 22968 5080
rect 13817 5043 13875 5049
rect 26142 5040 26148 5092
rect 26200 5080 26206 5092
rect 27341 5083 27399 5089
rect 27341 5080 27353 5083
rect 26200 5052 27353 5080
rect 26200 5040 26206 5052
rect 27341 5049 27353 5052
rect 27387 5049 27399 5083
rect 27341 5043 27399 5049
rect 1854 4972 1860 5024
rect 1912 5012 1918 5024
rect 2225 5015 2283 5021
rect 2225 5012 2237 5015
rect 1912 4984 2237 5012
rect 1912 4972 1918 4984
rect 2225 4981 2237 4984
rect 2271 4981 2283 5015
rect 2225 4975 2283 4981
rect 5353 5015 5411 5021
rect 5353 4981 5365 5015
rect 5399 5012 5411 5015
rect 5810 5012 5816 5024
rect 5399 4984 5816 5012
rect 5399 4981 5411 4984
rect 5353 4975 5411 4981
rect 5810 4972 5816 4984
rect 5868 4972 5874 5024
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 7101 5015 7159 5021
rect 7101 5012 7113 5015
rect 6972 4984 7113 5012
rect 6972 4972 6978 4984
rect 7101 4981 7113 4984
rect 7147 5012 7159 5015
rect 8202 5012 8208 5024
rect 7147 4984 8208 5012
rect 7147 4981 7159 4984
rect 7101 4975 7159 4981
rect 8202 4972 8208 4984
rect 8260 5012 8266 5024
rect 10413 5015 10471 5021
rect 10413 5012 10425 5015
rect 8260 4984 10425 5012
rect 8260 4972 8266 4984
rect 10413 4981 10425 4984
rect 10459 4981 10471 5015
rect 11790 5012 11796 5024
rect 11751 4984 11796 5012
rect 10413 4975 10471 4981
rect 11790 4972 11796 4984
rect 11848 4972 11854 5024
rect 11974 5012 11980 5024
rect 11935 4984 11980 5012
rect 11974 4972 11980 4984
rect 12032 4972 12038 5024
rect 15378 4972 15384 5024
rect 15436 5012 15442 5024
rect 18049 5015 18107 5021
rect 18049 5012 18061 5015
rect 15436 4984 18061 5012
rect 15436 4972 15442 4984
rect 18049 4981 18061 4984
rect 18095 4981 18107 5015
rect 18049 4975 18107 4981
rect 18414 4972 18420 5024
rect 18472 5012 18478 5024
rect 18601 5015 18659 5021
rect 18601 5012 18613 5015
rect 18472 4984 18613 5012
rect 18472 4972 18478 4984
rect 18601 4981 18613 4984
rect 18647 4981 18659 5015
rect 18601 4975 18659 4981
rect 19705 5015 19763 5021
rect 19705 4981 19717 5015
rect 19751 5012 19763 5015
rect 20346 5012 20352 5024
rect 19751 4984 20352 5012
rect 19751 4981 19763 4984
rect 19705 4975 19763 4981
rect 20346 4972 20352 4984
rect 20404 4972 20410 5024
rect 20441 5015 20499 5021
rect 20441 4981 20453 5015
rect 20487 5012 20499 5015
rect 20806 5012 20812 5024
rect 20487 4984 20812 5012
rect 20487 4981 20499 4984
rect 20441 4975 20499 4981
rect 20806 4972 20812 4984
rect 20864 4972 20870 5024
rect 20990 4972 20996 5024
rect 21048 5012 21054 5024
rect 21085 5015 21143 5021
rect 21085 5012 21097 5015
rect 21048 4984 21097 5012
rect 21048 4972 21054 4984
rect 21085 4981 21097 4984
rect 21131 4981 21143 5015
rect 21818 5012 21824 5024
rect 21779 4984 21824 5012
rect 21085 4975 21143 4981
rect 21818 4972 21824 4984
rect 21876 4972 21882 5024
rect 22738 4972 22744 5024
rect 22796 5012 22802 5024
rect 23017 5015 23075 5021
rect 23017 5012 23029 5015
rect 22796 4984 23029 5012
rect 22796 4972 22802 4984
rect 23017 4981 23029 4984
rect 23063 4981 23075 5015
rect 23017 4975 23075 4981
rect 23753 5015 23811 5021
rect 23753 4981 23765 5015
rect 23799 5012 23811 5015
rect 24210 5012 24216 5024
rect 23799 4984 24216 5012
rect 23799 4981 23811 4984
rect 23753 4975 23811 4981
rect 24210 4972 24216 4984
rect 24268 4972 24274 5024
rect 24569 4972 24575 5024
rect 24627 5012 24633 5024
rect 24627 4984 24672 5012
rect 24627 4972 24633 4984
rect 26878 4972 26884 5024
rect 26936 5012 26942 5024
rect 27157 5015 27215 5021
rect 27157 5012 27169 5015
rect 26936 4984 27169 5012
rect 26936 4972 26942 4984
rect 27157 4981 27169 4984
rect 27203 4981 27215 5015
rect 27157 4975 27215 4981
rect 1104 4922 28060 4944
rect 1104 4870 5442 4922
rect 5494 4870 5506 4922
rect 5558 4870 5570 4922
rect 5622 4870 5634 4922
rect 5686 4870 5698 4922
rect 5750 4870 14428 4922
rect 14480 4870 14492 4922
rect 14544 4870 14556 4922
rect 14608 4870 14620 4922
rect 14672 4870 14684 4922
rect 14736 4870 23413 4922
rect 23465 4870 23477 4922
rect 23529 4870 23541 4922
rect 23593 4870 23605 4922
rect 23657 4870 23669 4922
rect 23721 4870 28060 4922
rect 1104 4848 28060 4870
rect 3786 4808 3792 4820
rect 3747 4780 3792 4808
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 4246 4768 4252 4820
rect 4304 4768 4310 4820
rect 4890 4768 4896 4820
rect 4948 4808 4954 4820
rect 7745 4811 7803 4817
rect 7745 4808 7757 4811
rect 4948 4780 7757 4808
rect 4948 4768 4954 4780
rect 7745 4777 7757 4780
rect 7791 4777 7803 4811
rect 7745 4771 7803 4777
rect 8018 4768 8024 4820
rect 8076 4808 8082 4820
rect 8205 4811 8263 4817
rect 8205 4808 8217 4811
rect 8076 4780 8217 4808
rect 8076 4768 8082 4780
rect 8205 4777 8217 4780
rect 8251 4777 8263 4811
rect 9582 4808 9588 4820
rect 9543 4780 9588 4808
rect 8205 4771 8263 4777
rect 9582 4768 9588 4780
rect 9640 4768 9646 4820
rect 11514 4768 11520 4820
rect 11572 4808 11578 4820
rect 13541 4811 13599 4817
rect 13541 4808 13553 4811
rect 11572 4780 13553 4808
rect 11572 4768 11578 4780
rect 13541 4777 13553 4780
rect 13587 4777 13599 4811
rect 17126 4808 17132 4820
rect 17087 4780 17132 4808
rect 13541 4771 13599 4777
rect 17126 4768 17132 4780
rect 17184 4768 17190 4820
rect 17586 4768 17592 4820
rect 17644 4808 17650 4820
rect 17644 4780 20300 4808
rect 17644 4768 17650 4780
rect 4264 4740 4292 4768
rect 3988 4712 4292 4740
rect 1394 4604 1400 4616
rect 1307 4576 1400 4604
rect 1394 4564 1400 4576
rect 1452 4604 1458 4616
rect 2682 4604 2688 4616
rect 1452 4576 2688 4604
rect 1452 4564 1458 4576
rect 2682 4564 2688 4576
rect 2740 4564 2746 4616
rect 3988 4613 4016 4712
rect 4338 4700 4344 4752
rect 4396 4700 4402 4752
rect 6270 4700 6276 4752
rect 6328 4740 6334 4752
rect 6917 4743 6975 4749
rect 6917 4740 6929 4743
rect 6328 4712 6929 4740
rect 6328 4700 6334 4712
rect 6917 4709 6929 4712
rect 6963 4709 6975 4743
rect 6917 4703 6975 4709
rect 8294 4700 8300 4752
rect 8352 4740 8358 4752
rect 8478 4740 8484 4752
rect 8352 4712 8484 4740
rect 8352 4700 8358 4712
rect 8478 4700 8484 4712
rect 8536 4700 8542 4752
rect 10459 4743 10517 4749
rect 10459 4709 10471 4743
rect 10505 4740 10517 4743
rect 10594 4740 10600 4752
rect 10505 4712 10600 4740
rect 10505 4709 10517 4712
rect 10459 4703 10517 4709
rect 10594 4700 10600 4712
rect 10652 4740 10658 4752
rect 11882 4740 11888 4752
rect 10652 4712 11888 4740
rect 10652 4700 10658 4712
rect 11882 4700 11888 4712
rect 11940 4700 11946 4752
rect 20272 4740 20300 4780
rect 20346 4768 20352 4820
rect 20404 4808 20410 4820
rect 20404 4780 24256 4808
rect 20404 4768 20410 4780
rect 20530 4740 20536 4752
rect 20272 4712 20536 4740
rect 20530 4700 20536 4712
rect 20588 4700 20594 4752
rect 22094 4700 22100 4752
rect 22152 4740 22158 4752
rect 22152 4712 22232 4740
rect 22152 4700 22158 4712
rect 4249 4675 4307 4681
rect 4249 4641 4261 4675
rect 4295 4672 4307 4675
rect 4356 4672 4384 4700
rect 4295 4644 4384 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 6730 4632 6736 4684
rect 6788 4672 6794 4684
rect 7006 4672 7012 4684
rect 6788 4644 7012 4672
rect 6788 4632 6794 4644
rect 7006 4632 7012 4644
rect 7064 4632 7070 4684
rect 7466 4632 7472 4684
rect 7524 4672 7530 4684
rect 7837 4675 7895 4681
rect 7837 4672 7849 4675
rect 7524 4644 7849 4672
rect 7524 4632 7530 4644
rect 7837 4641 7849 4644
rect 7883 4641 7895 4675
rect 11974 4672 11980 4684
rect 7837 4635 7895 4641
rect 7944 4644 11980 4672
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4604 4399 4607
rect 4706 4604 4712 4616
rect 4387 4576 4712 4604
rect 4387 4573 4399 4576
rect 4341 4567 4399 4573
rect 1670 4545 1676 4548
rect 1664 4499 1676 4545
rect 1728 4536 1734 4548
rect 4080 4536 4108 4567
rect 4706 4564 4712 4576
rect 4764 4564 4770 4616
rect 5074 4604 5080 4616
rect 5035 4576 5080 4604
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 6546 4564 6552 4616
rect 6604 4604 6610 4616
rect 7101 4607 7159 4613
rect 7101 4604 7113 4607
rect 6604 4576 7113 4604
rect 6604 4564 6610 4576
rect 7101 4573 7113 4576
rect 7147 4573 7159 4607
rect 7101 4567 7159 4573
rect 7745 4607 7803 4613
rect 7745 4573 7757 4607
rect 7791 4604 7803 4607
rect 7944 4604 7972 4644
rect 11974 4632 11980 4644
rect 12032 4632 12038 4684
rect 16390 4672 16396 4684
rect 14752 4644 16396 4672
rect 7791 4576 7972 4604
rect 8021 4607 8079 4613
rect 7791 4573 7803 4576
rect 7745 4567 7803 4573
rect 8021 4573 8033 4607
rect 8067 4573 8079 4607
rect 8021 4567 8079 4573
rect 4246 4536 4252 4548
rect 1728 4508 1764 4536
rect 2792 4508 4252 4536
rect 1670 4496 1676 4499
rect 1728 4496 1734 4508
rect 2792 4477 2820 4508
rect 4246 4496 4252 4508
rect 4304 4496 4310 4548
rect 5350 4545 5356 4548
rect 5344 4499 5356 4545
rect 5408 4536 5414 4548
rect 8036 4536 8064 4567
rect 9214 4564 9220 4616
rect 9272 4604 9278 4616
rect 9309 4607 9367 4613
rect 9309 4604 9321 4607
rect 9272 4576 9321 4604
rect 9272 4564 9278 4576
rect 9309 4573 9321 4576
rect 9355 4573 9367 4607
rect 9490 4604 9496 4616
rect 9451 4576 9496 4604
rect 9309 4567 9367 4573
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 9585 4607 9643 4613
rect 9585 4573 9597 4607
rect 9631 4604 9643 4607
rect 9858 4604 9864 4616
rect 9631 4576 9864 4604
rect 9631 4573 9643 4576
rect 9585 4567 9643 4573
rect 9858 4564 9864 4576
rect 9916 4564 9922 4616
rect 10226 4604 10232 4616
rect 10187 4576 10232 4604
rect 10226 4564 10232 4576
rect 10284 4564 10290 4616
rect 11698 4604 11704 4616
rect 11659 4576 11704 4604
rect 11698 4564 11704 4576
rect 11756 4564 11762 4616
rect 12161 4607 12219 4613
rect 12161 4573 12173 4607
rect 12207 4604 12219 4607
rect 12207 4576 12572 4604
rect 12207 4573 12219 4576
rect 12161 4567 12219 4573
rect 12544 4548 12572 4576
rect 12802 4564 12808 4616
rect 12860 4604 12866 4616
rect 14090 4604 14096 4616
rect 12860 4576 14096 4604
rect 12860 4564 12866 4576
rect 14090 4564 14096 4576
rect 14148 4564 14154 4616
rect 14752 4613 14780 4644
rect 16390 4632 16396 4644
rect 16448 4632 16454 4684
rect 17310 4632 17316 4684
rect 17368 4672 17374 4684
rect 19245 4675 19303 4681
rect 19245 4672 19257 4675
rect 17368 4644 19257 4672
rect 17368 4632 17374 4644
rect 19245 4641 19257 4644
rect 19291 4641 19303 4675
rect 19245 4635 19303 4641
rect 22204 4672 22232 4712
rect 22830 4700 22836 4752
rect 22888 4740 22894 4752
rect 22888 4712 23244 4740
rect 22888 4700 22894 4712
rect 22278 4672 22284 4684
rect 22204 4644 22284 4672
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 14737 4607 14795 4613
rect 14737 4573 14749 4607
rect 14783 4573 14795 4607
rect 15470 4604 15476 4616
rect 15431 4576 15476 4604
rect 14737 4567 14795 4573
rect 5408 4508 5444 4536
rect 8036 4508 9812 4536
rect 5350 4496 5356 4499
rect 5408 4496 5414 4508
rect 2777 4471 2835 4477
rect 2777 4437 2789 4471
rect 2823 4437 2835 4471
rect 2777 4431 2835 4437
rect 6457 4471 6515 4477
rect 6457 4437 6469 4471
rect 6503 4468 6515 4471
rect 6730 4468 6736 4480
rect 6503 4440 6736 4468
rect 6503 4437 6515 4440
rect 6457 4431 6515 4437
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 9784 4477 9812 4508
rect 10778 4496 10784 4548
rect 10836 4536 10842 4548
rect 12406 4539 12464 4545
rect 12406 4536 12418 4539
rect 10836 4508 12418 4536
rect 10836 4496 10842 4508
rect 12406 4505 12418 4508
rect 12452 4505 12464 4539
rect 12406 4499 12464 4505
rect 12526 4496 12532 4548
rect 12584 4496 12590 4548
rect 12710 4496 12716 4548
rect 12768 4536 12774 4548
rect 13170 4536 13176 4548
rect 12768 4508 13176 4536
rect 12768 4496 12774 4508
rect 13170 4496 13176 4508
rect 13228 4496 13234 4548
rect 14292 4536 14320 4567
rect 15470 4564 15476 4576
rect 15528 4564 15534 4616
rect 16206 4564 16212 4616
rect 16264 4604 16270 4616
rect 16761 4607 16819 4613
rect 16761 4604 16773 4607
rect 16264 4576 16773 4604
rect 16264 4564 16270 4576
rect 16761 4573 16773 4576
rect 16807 4573 16819 4607
rect 16761 4567 16819 4573
rect 17589 4607 17647 4613
rect 17589 4573 17601 4607
rect 17635 4573 17647 4607
rect 17589 4567 17647 4573
rect 18325 4607 18383 4613
rect 18325 4573 18337 4607
rect 18371 4604 18383 4607
rect 20530 4604 20536 4616
rect 18371 4576 20536 4604
rect 18371 4573 18383 4576
rect 18325 4567 18383 4573
rect 15286 4536 15292 4548
rect 14292 4508 15292 4536
rect 15286 4496 15292 4508
rect 15344 4496 15350 4548
rect 16666 4496 16672 4548
rect 16724 4536 16730 4548
rect 16945 4539 17003 4545
rect 16945 4536 16957 4539
rect 16724 4508 16957 4536
rect 16724 4496 16730 4508
rect 16945 4505 16957 4508
rect 16991 4505 17003 4539
rect 17604 4536 17632 4567
rect 20530 4564 20536 4576
rect 20588 4564 20594 4616
rect 21085 4607 21143 4613
rect 21085 4573 21097 4607
rect 21131 4604 21143 4607
rect 22204 4604 22232 4644
rect 22278 4632 22284 4644
rect 22336 4632 22342 4684
rect 23014 4604 23020 4616
rect 21131 4576 22232 4604
rect 22296 4576 23020 4604
rect 21131 4573 21143 4576
rect 21085 4567 21143 4573
rect 19058 4536 19064 4548
rect 17604 4508 19064 4536
rect 16945 4499 17003 4505
rect 19058 4496 19064 4508
rect 19116 4496 19122 4548
rect 19512 4539 19570 4545
rect 19512 4505 19524 4539
rect 19558 4536 19570 4539
rect 20254 4536 20260 4548
rect 19558 4508 20260 4536
rect 19558 4505 19570 4508
rect 19512 4499 19570 4505
rect 20254 4496 20260 4508
rect 20312 4496 20318 4548
rect 21352 4539 21410 4545
rect 21352 4505 21364 4539
rect 21398 4536 21410 4539
rect 21818 4536 21824 4548
rect 21398 4508 21824 4536
rect 21398 4505 21410 4508
rect 21352 4499 21410 4505
rect 21818 4496 21824 4508
rect 21876 4496 21882 4548
rect 9769 4471 9827 4477
rect 9769 4437 9781 4471
rect 9815 4437 9827 4471
rect 9769 4431 9827 4437
rect 11517 4471 11575 4477
rect 11517 4437 11529 4471
rect 11563 4468 11575 4471
rect 13262 4468 13268 4480
rect 11563 4440 13268 4468
rect 11563 4437 11575 4440
rect 11517 4431 11575 4437
rect 13262 4428 13268 4440
rect 13320 4428 13326 4480
rect 13814 4428 13820 4480
rect 13872 4468 13878 4480
rect 14093 4471 14151 4477
rect 14093 4468 14105 4471
rect 13872 4440 14105 4468
rect 13872 4428 13878 4440
rect 14093 4437 14105 4440
rect 14139 4437 14151 4471
rect 14093 4431 14151 4437
rect 14826 4428 14832 4480
rect 14884 4468 14890 4480
rect 14921 4471 14979 4477
rect 14921 4468 14933 4471
rect 14884 4440 14933 4468
rect 14884 4428 14890 4440
rect 14921 4437 14933 4440
rect 14967 4437 14979 4471
rect 14921 4431 14979 4437
rect 15194 4428 15200 4480
rect 15252 4468 15258 4480
rect 15657 4471 15715 4477
rect 15657 4468 15669 4471
rect 15252 4440 15669 4468
rect 15252 4428 15258 4440
rect 15657 4437 15669 4440
rect 15703 4437 15715 4471
rect 15657 4431 15715 4437
rect 16574 4428 16580 4480
rect 16632 4468 16638 4480
rect 17773 4471 17831 4477
rect 17773 4468 17785 4471
rect 16632 4440 17785 4468
rect 16632 4428 16638 4440
rect 17773 4437 17785 4440
rect 17819 4437 17831 4471
rect 17773 4431 17831 4437
rect 17954 4428 17960 4480
rect 18012 4468 18018 4480
rect 18509 4471 18567 4477
rect 18509 4468 18521 4471
rect 18012 4440 18521 4468
rect 18012 4428 18018 4440
rect 18509 4437 18521 4440
rect 18555 4437 18567 4471
rect 20622 4468 20628 4480
rect 20583 4440 20628 4468
rect 18509 4431 18567 4437
rect 20622 4428 20628 4440
rect 20680 4428 20686 4480
rect 21542 4428 21548 4480
rect 21600 4468 21606 4480
rect 22296 4468 22324 4576
rect 23014 4564 23020 4576
rect 23072 4564 23078 4616
rect 23109 4607 23167 4613
rect 23109 4573 23121 4607
rect 23155 4604 23167 4607
rect 23216 4604 23244 4712
rect 23290 4700 23296 4752
rect 23348 4700 23354 4752
rect 23308 4672 23336 4700
rect 24228 4672 24256 4780
rect 24302 4768 24308 4820
rect 24360 4808 24366 4820
rect 26142 4808 26148 4820
rect 24360 4780 26148 4808
rect 24360 4768 24366 4780
rect 26142 4768 26148 4780
rect 26200 4768 26206 4820
rect 26878 4808 26884 4820
rect 26839 4780 26884 4808
rect 26878 4768 26884 4780
rect 26936 4768 26942 4820
rect 25774 4700 25780 4752
rect 25832 4740 25838 4752
rect 27065 4743 27123 4749
rect 27065 4740 27077 4743
rect 25832 4712 27077 4740
rect 25832 4700 25838 4712
rect 27065 4709 27077 4712
rect 27111 4709 27123 4743
rect 27065 4703 27123 4709
rect 23308 4644 24180 4672
rect 24228 4644 24716 4672
rect 23382 4604 23388 4616
rect 23155 4576 23244 4604
rect 23343 4576 23388 4604
rect 23155 4573 23167 4576
rect 23109 4567 23167 4573
rect 23382 4564 23388 4576
rect 23440 4564 23446 4616
rect 24152 4604 24180 4644
rect 24302 4604 24308 4616
rect 24152 4576 24308 4604
rect 24302 4564 24308 4576
rect 24360 4564 24366 4616
rect 24581 4607 24639 4613
rect 24581 4573 24593 4607
rect 24627 4573 24639 4607
rect 24688 4604 24716 4644
rect 27154 4604 27160 4616
rect 24688 4576 27160 4604
rect 24581 4567 24639 4573
rect 22554 4496 22560 4548
rect 22612 4536 22618 4548
rect 24596 4536 24624 4567
rect 27154 4564 27160 4576
rect 27212 4564 27218 4616
rect 24854 4545 24860 4548
rect 22612 4508 24624 4536
rect 22612 4496 22618 4508
rect 24848 4499 24860 4545
rect 24912 4536 24918 4548
rect 26694 4536 26700 4548
rect 24912 4508 24948 4536
rect 26655 4508 26700 4536
rect 24854 4496 24860 4499
rect 24912 4496 24918 4508
rect 26694 4496 26700 4508
rect 26752 4496 26758 4548
rect 26970 4545 26976 4548
rect 26913 4539 26976 4545
rect 26913 4505 26925 4539
rect 26959 4505 26976 4539
rect 26913 4499 26976 4505
rect 26970 4496 26976 4499
rect 27028 4496 27034 4548
rect 22462 4468 22468 4480
rect 21600 4440 22324 4468
rect 22423 4440 22468 4468
rect 21600 4428 21606 4440
rect 22462 4428 22468 4440
rect 22520 4428 22526 4480
rect 22922 4468 22928 4480
rect 22883 4440 22928 4468
rect 22922 4428 22928 4440
rect 22980 4428 22986 4480
rect 23293 4471 23351 4477
rect 23293 4437 23305 4471
rect 23339 4468 23351 4471
rect 23474 4468 23480 4480
rect 23339 4440 23480 4468
rect 23339 4437 23351 4440
rect 23293 4431 23351 4437
rect 23474 4428 23480 4440
rect 23532 4428 23538 4480
rect 24394 4428 24400 4480
rect 24452 4468 24458 4480
rect 25961 4471 26019 4477
rect 25961 4468 25973 4471
rect 24452 4440 25973 4468
rect 24452 4428 24458 4440
rect 25961 4437 25973 4440
rect 26007 4437 26019 4471
rect 25961 4431 26019 4437
rect 1104 4378 28060 4400
rect 1104 4326 9935 4378
rect 9987 4326 9999 4378
rect 10051 4326 10063 4378
rect 10115 4326 10127 4378
rect 10179 4326 10191 4378
rect 10243 4326 18920 4378
rect 18972 4326 18984 4378
rect 19036 4326 19048 4378
rect 19100 4326 19112 4378
rect 19164 4326 19176 4378
rect 19228 4326 28060 4378
rect 1104 4304 28060 4326
rect 1670 4264 1676 4276
rect 1631 4236 1676 4264
rect 1670 4224 1676 4236
rect 1728 4224 1734 4276
rect 3418 4224 3424 4276
rect 3476 4264 3482 4276
rect 4338 4264 4344 4276
rect 3476 4236 4344 4264
rect 3476 4224 3482 4236
rect 4338 4224 4344 4236
rect 4396 4224 4402 4276
rect 4890 4264 4896 4276
rect 4851 4236 4896 4264
rect 4890 4224 4896 4236
rect 4948 4224 4954 4276
rect 5350 4264 5356 4276
rect 5311 4236 5356 4264
rect 5350 4224 5356 4236
rect 5408 4224 5414 4276
rect 7742 4264 7748 4276
rect 7576 4236 7748 4264
rect 2958 4156 2964 4208
rect 3016 4196 3022 4208
rect 3016 4168 3096 4196
rect 3016 4156 3022 4168
rect 842 4088 848 4140
rect 900 4128 906 4140
rect 1486 4128 1492 4140
rect 900 4100 1492 4128
rect 900 4088 906 4100
rect 1486 4088 1492 4100
rect 1544 4088 1550 4140
rect 1854 4128 1860 4140
rect 1815 4100 1860 4128
rect 1854 4088 1860 4100
rect 1912 4088 1918 4140
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4128 2651 4131
rect 2682 4128 2688 4140
rect 2639 4100 2688 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 2682 4088 2688 4100
rect 2740 4088 2746 4140
rect 2866 4137 2872 4140
rect 2860 4091 2872 4137
rect 2924 4128 2930 4140
rect 3068 4128 3096 4168
rect 4246 4156 4252 4208
rect 4304 4196 4310 4208
rect 4433 4199 4491 4205
rect 4433 4196 4445 4199
rect 4304 4168 4445 4196
rect 4304 4156 4310 4168
rect 4433 4165 4445 4168
rect 4479 4165 4491 4199
rect 4433 4159 4491 4165
rect 4540 4168 4844 4196
rect 2924 4100 2960 4128
rect 3068 4100 3648 4128
rect 2866 4088 2872 4091
rect 2924 4088 2930 4100
rect 3620 4060 3648 4100
rect 3970 4088 3976 4140
rect 4028 4128 4034 4140
rect 4540 4128 4568 4168
rect 4706 4128 4712 4140
rect 4028 4100 4568 4128
rect 4667 4100 4712 4128
rect 4028 4088 4034 4100
rect 4706 4088 4712 4100
rect 4764 4088 4770 4140
rect 4430 4060 4436 4072
rect 3620 4032 4436 4060
rect 4430 4020 4436 4032
rect 4488 4020 4494 4072
rect 4614 4060 4620 4072
rect 4575 4032 4620 4060
rect 4614 4020 4620 4032
rect 4672 4020 4678 4072
rect 4816 4060 4844 4168
rect 6546 4156 6552 4208
rect 6604 4196 6610 4208
rect 6604 4168 6960 4196
rect 6604 4156 6610 4168
rect 4982 4088 4988 4140
rect 5040 4128 5046 4140
rect 5350 4128 5356 4140
rect 5040 4100 5356 4128
rect 5040 4088 5046 4100
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 5537 4131 5595 4137
rect 5537 4097 5549 4131
rect 5583 4128 5595 4131
rect 5810 4128 5816 4140
rect 5583 4100 5816 4128
rect 5583 4097 5595 4100
rect 5537 4091 5595 4097
rect 5810 4088 5816 4100
rect 5868 4088 5874 4140
rect 6454 4128 6460 4140
rect 6415 4100 6460 4128
rect 6454 4088 6460 4100
rect 6512 4088 6518 4140
rect 6638 4128 6644 4140
rect 6599 4100 6644 4128
rect 6638 4088 6644 4100
rect 6696 4088 6702 4140
rect 6730 4088 6736 4140
rect 6788 4128 6794 4140
rect 6932 4128 6960 4168
rect 7576 4137 7604 4236
rect 7742 4224 7748 4236
rect 7800 4224 7806 4276
rect 7837 4267 7895 4273
rect 7837 4233 7849 4267
rect 7883 4264 7895 4267
rect 8018 4264 8024 4276
rect 7883 4236 8024 4264
rect 7883 4233 7895 4236
rect 7837 4227 7895 4233
rect 8018 4224 8024 4236
rect 8076 4224 8082 4276
rect 8202 4224 8208 4276
rect 8260 4264 8266 4276
rect 8260 4236 8432 4264
rect 8260 4224 8266 4236
rect 7009 4131 7067 4137
rect 7009 4128 7021 4131
rect 6788 4100 6833 4128
rect 6932 4100 7021 4128
rect 6788 4088 6794 4100
rect 7009 4097 7021 4100
rect 7055 4097 7067 4131
rect 7009 4091 7067 4097
rect 7561 4131 7619 4137
rect 7561 4097 7573 4131
rect 7607 4097 7619 4131
rect 7561 4091 7619 4097
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4128 7711 4131
rect 7742 4128 7748 4140
rect 7699 4100 7748 4128
rect 7699 4097 7711 4100
rect 7653 4091 7711 4097
rect 5902 4060 5908 4072
rect 4816 4032 5908 4060
rect 5902 4020 5908 4032
rect 5960 4020 5966 4072
rect 6178 4020 6184 4072
rect 6236 4060 6242 4072
rect 6546 4060 6552 4072
rect 6236 4032 6552 4060
rect 6236 4020 6242 4032
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 6914 4060 6920 4072
rect 6875 4032 6920 4060
rect 6914 4020 6920 4032
rect 6972 4020 6978 4072
rect 7576 4060 7604 4091
rect 7742 4088 7748 4100
rect 7800 4088 7806 4140
rect 7834 4088 7840 4140
rect 7892 4128 7898 4140
rect 8202 4128 8208 4140
rect 7892 4100 8208 4128
rect 7892 4088 7898 4100
rect 8202 4088 8208 4100
rect 8260 4128 8266 4140
rect 8297 4131 8355 4137
rect 8297 4128 8309 4131
rect 8260 4100 8309 4128
rect 8260 4088 8266 4100
rect 8297 4097 8309 4100
rect 8343 4097 8355 4131
rect 8404 4128 8432 4236
rect 10502 4224 10508 4276
rect 10560 4264 10566 4276
rect 10870 4264 10876 4276
rect 10560 4236 10876 4264
rect 10560 4224 10566 4236
rect 10870 4224 10876 4236
rect 10928 4224 10934 4276
rect 11698 4224 11704 4276
rect 11756 4264 11762 4276
rect 13170 4264 13176 4276
rect 11756 4236 13176 4264
rect 11756 4224 11762 4236
rect 13170 4224 13176 4236
rect 13228 4224 13234 4276
rect 18708 4236 21128 4264
rect 10686 4156 10692 4208
rect 10744 4196 10750 4208
rect 12897 4199 12955 4205
rect 12897 4196 12909 4199
rect 10744 4168 12909 4196
rect 10744 4156 10750 4168
rect 12897 4165 12909 4168
rect 12943 4165 12955 4199
rect 12897 4159 12955 4165
rect 15749 4199 15807 4205
rect 15749 4165 15761 4199
rect 15795 4196 15807 4199
rect 17586 4196 17592 4208
rect 15795 4168 17592 4196
rect 15795 4165 15807 4168
rect 15749 4159 15807 4165
rect 17586 4156 17592 4168
rect 17644 4156 17650 4208
rect 18708 4205 18736 4236
rect 18693 4199 18751 4205
rect 18693 4165 18705 4199
rect 18739 4165 18751 4199
rect 18693 4159 18751 4165
rect 19518 4156 19524 4208
rect 19576 4196 19582 4208
rect 19576 4168 20668 4196
rect 19576 4156 19582 4168
rect 8553 4131 8611 4137
rect 8553 4128 8565 4131
rect 8404 4100 8565 4128
rect 8297 4091 8355 4097
rect 8553 4097 8565 4100
rect 8599 4097 8611 4131
rect 8553 4091 8611 4097
rect 9122 4088 9128 4140
rect 9180 4128 9186 4140
rect 10778 4128 10784 4140
rect 9180 4100 10784 4128
rect 9180 4088 9186 4100
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 11514 4128 11520 4140
rect 11475 4100 11520 4128
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 11974 4137 11980 4140
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4097 11759 4131
rect 11701 4091 11759 4097
rect 11789 4131 11847 4137
rect 11789 4097 11801 4131
rect 11835 4097 11847 4131
rect 11789 4091 11847 4097
rect 11931 4131 11980 4137
rect 11931 4097 11943 4131
rect 11977 4097 11980 4131
rect 11931 4091 11980 4097
rect 7576 4032 7880 4060
rect 7852 4004 7880 4032
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 9950 4060 9956 4072
rect 9456 4032 9956 4060
rect 9456 4020 9462 4032
rect 9950 4020 9956 4032
rect 10008 4020 10014 4072
rect 10137 4063 10195 4069
rect 10137 4029 10149 4063
rect 10183 4029 10195 4063
rect 10137 4023 10195 4029
rect 10413 4063 10471 4069
rect 10413 4029 10425 4063
rect 10459 4060 10471 4063
rect 10870 4060 10876 4072
rect 10459 4032 10876 4060
rect 10459 4029 10471 4032
rect 10413 4023 10471 4029
rect 4246 3952 4252 4004
rect 4304 3992 4310 4004
rect 4798 3992 4804 4004
rect 4304 3964 4804 3992
rect 4304 3952 4310 3964
rect 4798 3952 4804 3964
rect 4856 3952 4862 4004
rect 5258 3952 5264 4004
rect 5316 3992 5322 4004
rect 6638 3992 6644 4004
rect 5316 3964 6644 3992
rect 5316 3952 5322 3964
rect 6638 3952 6644 3964
rect 6696 3952 6702 4004
rect 7190 3952 7196 4004
rect 7248 3992 7254 4004
rect 7248 3964 7696 3992
rect 7248 3952 7254 3964
rect 2866 3884 2872 3936
rect 2924 3924 2930 3936
rect 3326 3924 3332 3936
rect 2924 3896 3332 3924
rect 2924 3884 2930 3896
rect 3326 3884 3332 3896
rect 3384 3884 3390 3936
rect 3973 3927 4031 3933
rect 3973 3893 3985 3927
rect 4019 3924 4031 3927
rect 4062 3924 4068 3936
rect 4019 3896 4068 3924
rect 4019 3893 4031 3896
rect 3973 3887 4031 3893
rect 4062 3884 4068 3896
rect 4120 3924 4126 3936
rect 4433 3927 4491 3933
rect 4433 3924 4445 3927
rect 4120 3896 4445 3924
rect 4120 3884 4126 3896
rect 4433 3893 4445 3896
rect 4479 3893 4491 3927
rect 4433 3887 4491 3893
rect 6362 3884 6368 3936
rect 6420 3924 6426 3936
rect 6822 3924 6828 3936
rect 6420 3896 6828 3924
rect 6420 3884 6426 3896
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 7558 3924 7564 3936
rect 6972 3896 7564 3924
rect 6972 3884 6978 3896
rect 7558 3884 7564 3896
rect 7616 3884 7622 3936
rect 7668 3924 7696 3964
rect 7834 3952 7840 4004
rect 7892 3952 7898 4004
rect 9490 3952 9496 4004
rect 9548 3992 9554 4004
rect 9677 3995 9735 4001
rect 9677 3992 9689 3995
rect 9548 3964 9689 3992
rect 9548 3952 9554 3964
rect 9677 3961 9689 3964
rect 9723 3961 9735 3995
rect 9677 3955 9735 3961
rect 9214 3924 9220 3936
rect 7668 3896 9220 3924
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 10152 3924 10180 4023
rect 10870 4020 10876 4032
rect 10928 4060 10934 4072
rect 11716 4060 11744 4091
rect 10928 4032 11744 4060
rect 10928 4020 10934 4032
rect 10318 3952 10324 4004
rect 10376 3992 10382 4004
rect 10686 3992 10692 4004
rect 10376 3964 10692 3992
rect 10376 3952 10382 3964
rect 10686 3952 10692 3964
rect 10744 3952 10750 4004
rect 11238 3952 11244 4004
rect 11296 3992 11302 4004
rect 11698 3992 11704 4004
rect 11296 3964 11704 3992
rect 11296 3952 11302 3964
rect 11698 3952 11704 3964
rect 11756 3952 11762 4004
rect 10410 3924 10416 3936
rect 10152 3896 10416 3924
rect 10410 3884 10416 3896
rect 10468 3884 10474 3936
rect 10962 3884 10968 3936
rect 11020 3924 11026 3936
rect 11799 3924 11827 4091
rect 11974 4088 11980 4091
rect 12032 4088 12038 4140
rect 12713 4131 12771 4137
rect 12713 4128 12725 4131
rect 12084 4100 12725 4128
rect 12084 4001 12112 4100
rect 12713 4097 12725 4100
rect 12759 4097 12771 4131
rect 12713 4091 12771 4097
rect 13357 4131 13415 4137
rect 13357 4097 13369 4131
rect 13403 4128 13415 4131
rect 13814 4128 13820 4140
rect 13403 4100 13820 4128
rect 13403 4097 13415 4100
rect 13357 4091 13415 4097
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 14093 4131 14151 4137
rect 14093 4097 14105 4131
rect 14139 4097 14151 4131
rect 14093 4091 14151 4097
rect 14829 4131 14887 4137
rect 14829 4097 14841 4131
rect 14875 4128 14887 4131
rect 14918 4128 14924 4140
rect 14875 4100 14924 4128
rect 14875 4097 14887 4100
rect 14829 4091 14887 4097
rect 12529 4063 12587 4069
rect 12529 4029 12541 4063
rect 12575 4029 12587 4063
rect 12529 4023 12587 4029
rect 12069 3995 12127 4001
rect 12069 3961 12081 3995
rect 12115 3961 12127 3995
rect 12069 3955 12127 3961
rect 12434 3952 12440 4004
rect 12492 3992 12498 4004
rect 12544 3992 12572 4023
rect 13262 4020 13268 4072
rect 13320 4060 13326 4072
rect 14108 4060 14136 4091
rect 14918 4088 14924 4100
rect 14976 4088 14982 4140
rect 16669 4131 16727 4137
rect 16669 4097 16681 4131
rect 16715 4128 16727 4131
rect 16758 4128 16764 4140
rect 16715 4100 16764 4128
rect 16715 4097 16727 4100
rect 16669 4091 16727 4097
rect 16758 4088 16764 4100
rect 16816 4088 16822 4140
rect 17773 4131 17831 4137
rect 17773 4097 17785 4131
rect 17819 4128 17831 4131
rect 18138 4128 18144 4140
rect 17819 4100 18144 4128
rect 17819 4097 17831 4100
rect 17773 4091 17831 4097
rect 18138 4088 18144 4100
rect 18196 4088 18202 4140
rect 19334 4128 19340 4140
rect 18248 4100 19340 4128
rect 13320 4032 14136 4060
rect 13320 4020 13326 4032
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 18046 4060 18052 4072
rect 16264 4032 18052 4060
rect 16264 4020 16270 4032
rect 18046 4020 18052 4032
rect 18104 4020 18110 4072
rect 18248 4069 18276 4100
rect 19334 4088 19340 4100
rect 19392 4088 19398 4140
rect 19613 4131 19671 4137
rect 19613 4097 19625 4131
rect 19659 4128 19671 4131
rect 20438 4128 20444 4140
rect 19659 4100 20444 4128
rect 19659 4097 19671 4100
rect 19613 4091 19671 4097
rect 20438 4088 20444 4100
rect 20496 4088 20502 4140
rect 20533 4131 20591 4137
rect 20533 4097 20545 4131
rect 20579 4097 20591 4131
rect 20640 4128 20668 4168
rect 20993 4131 21051 4137
rect 20993 4128 21005 4131
rect 20640 4100 21005 4128
rect 20533 4091 20591 4097
rect 20993 4097 21005 4100
rect 21039 4097 21051 4131
rect 21100 4128 21128 4236
rect 23474 4224 23480 4276
rect 23532 4264 23538 4276
rect 23750 4264 23756 4276
rect 23532 4236 23756 4264
rect 23532 4224 23538 4236
rect 23750 4224 23756 4236
rect 23808 4264 23814 4276
rect 23845 4267 23903 4273
rect 23845 4264 23857 4267
rect 23808 4236 23857 4264
rect 23808 4224 23814 4236
rect 23845 4233 23857 4236
rect 23891 4233 23903 4267
rect 23845 4227 23903 4233
rect 24394 4224 24400 4276
rect 24452 4264 24458 4276
rect 24765 4267 24823 4273
rect 24765 4264 24777 4267
rect 24452 4236 24777 4264
rect 24452 4224 24458 4236
rect 24765 4233 24777 4236
rect 24811 4233 24823 4267
rect 24765 4227 24823 4233
rect 26142 4224 26148 4276
rect 26200 4264 26206 4276
rect 26329 4267 26387 4273
rect 26329 4264 26341 4267
rect 26200 4236 26341 4264
rect 26200 4224 26206 4236
rect 26329 4233 26341 4236
rect 26375 4233 26387 4267
rect 26329 4227 26387 4233
rect 26878 4224 26884 4276
rect 26936 4264 26942 4276
rect 27173 4267 27231 4273
rect 27173 4264 27185 4267
rect 26936 4236 27185 4264
rect 26936 4224 26942 4236
rect 27173 4233 27185 4236
rect 27219 4233 27231 4267
rect 27173 4227 27231 4233
rect 22094 4156 22100 4208
rect 22152 4156 22158 4208
rect 22732 4199 22790 4205
rect 22732 4165 22744 4199
rect 22778 4196 22790 4199
rect 22922 4196 22928 4208
rect 22778 4168 22928 4196
rect 22778 4165 22790 4168
rect 22732 4159 22790 4165
rect 22922 4156 22928 4168
rect 22980 4156 22986 4208
rect 26234 4196 26240 4208
rect 26195 4168 26240 4196
rect 26234 4156 26240 4168
rect 26292 4156 26298 4208
rect 26786 4156 26792 4208
rect 26844 4196 26850 4208
rect 26973 4199 27031 4205
rect 26973 4196 26985 4199
rect 26844 4168 26985 4196
rect 26844 4156 26850 4168
rect 26973 4165 26985 4168
rect 27019 4165 27031 4199
rect 26973 4159 27031 4165
rect 21726 4128 21732 4140
rect 21100 4100 21732 4128
rect 20993 4091 21051 4097
rect 18233 4063 18291 4069
rect 18233 4029 18245 4063
rect 18279 4029 18291 4063
rect 18233 4023 18291 4029
rect 19153 4063 19211 4069
rect 19153 4029 19165 4063
rect 19199 4060 19211 4063
rect 19426 4060 19432 4072
rect 19199 4032 19432 4060
rect 19199 4029 19211 4032
rect 19153 4023 19211 4029
rect 19426 4020 19432 4032
rect 19484 4020 19490 4072
rect 19518 4020 19524 4072
rect 19576 4060 19582 4072
rect 20548 4060 20576 4091
rect 21726 4088 21732 4100
rect 21784 4088 21790 4140
rect 22005 4131 22063 4137
rect 22005 4097 22017 4131
rect 22051 4097 22063 4131
rect 22112 4128 22140 4156
rect 22370 4128 22376 4140
rect 22112 4100 22376 4128
rect 22005 4091 22063 4097
rect 22020 4060 22048 4091
rect 22370 4088 22376 4100
rect 22428 4088 22434 4140
rect 22554 4128 22560 4140
rect 22480 4100 22560 4128
rect 19576 4032 20576 4060
rect 20640 4032 22048 4060
rect 19576 4020 19582 4032
rect 13354 3992 13360 4004
rect 12492 3964 13360 3992
rect 12492 3952 12498 3964
rect 13354 3952 13360 3964
rect 13412 3952 13418 4004
rect 14090 3952 14096 4004
rect 14148 3992 14154 4004
rect 15013 3995 15071 4001
rect 15013 3992 15025 3995
rect 14148 3964 15025 3992
rect 14148 3952 14154 3964
rect 15013 3961 15025 3964
rect 15059 3961 15071 3995
rect 15013 3955 15071 3961
rect 15746 3952 15752 4004
rect 15804 3992 15810 4004
rect 16853 3995 16911 4001
rect 16853 3992 16865 3995
rect 15804 3964 16865 3992
rect 15804 3952 15810 3964
rect 16853 3961 16865 3964
rect 16899 3961 16911 3995
rect 16853 3955 16911 3961
rect 18141 3995 18199 4001
rect 18141 3961 18153 3995
rect 18187 3992 18199 3995
rect 18598 3992 18604 4004
rect 18187 3964 18604 3992
rect 18187 3961 18199 3964
rect 18141 3955 18199 3961
rect 18598 3952 18604 3964
rect 18656 3992 18662 4004
rect 18969 3995 19027 4001
rect 18969 3992 18981 3995
rect 18656 3964 18981 3992
rect 18656 3952 18662 3964
rect 18969 3961 18981 3964
rect 19015 3961 19027 3995
rect 20349 3995 20407 4001
rect 20349 3992 20361 3995
rect 18969 3955 19027 3961
rect 19076 3964 20361 3992
rect 11020 3896 11827 3924
rect 11020 3884 11026 3896
rect 12986 3884 12992 3936
rect 13044 3924 13050 3936
rect 13541 3927 13599 3933
rect 13541 3924 13553 3927
rect 13044 3896 13553 3924
rect 13044 3884 13050 3896
rect 13541 3893 13553 3896
rect 13587 3893 13599 3927
rect 13541 3887 13599 3893
rect 13630 3884 13636 3936
rect 13688 3924 13694 3936
rect 14277 3927 14335 3933
rect 14277 3924 14289 3927
rect 13688 3896 14289 3924
rect 13688 3884 13694 3896
rect 14277 3893 14289 3896
rect 14323 3893 14335 3927
rect 14277 3887 14335 3893
rect 15841 3927 15899 3933
rect 15841 3893 15853 3927
rect 15887 3924 15899 3927
rect 16206 3924 16212 3936
rect 15887 3896 16212 3924
rect 15887 3893 15899 3896
rect 15841 3887 15899 3893
rect 16206 3884 16212 3896
rect 16264 3884 16270 3936
rect 16390 3884 16396 3936
rect 16448 3924 16454 3936
rect 19076 3924 19104 3964
rect 20349 3961 20361 3964
rect 20395 3961 20407 3995
rect 20349 3955 20407 3961
rect 20438 3952 20444 4004
rect 20496 3992 20502 4004
rect 20640 3992 20668 4032
rect 22094 4020 22100 4072
rect 22152 4060 22158 4072
rect 22278 4060 22284 4072
rect 22152 4032 22284 4060
rect 22152 4020 22158 4032
rect 22278 4020 22284 4032
rect 22336 4060 22342 4072
rect 22480 4069 22508 4100
rect 22554 4088 22560 4100
rect 22612 4088 22618 4140
rect 23014 4088 23020 4140
rect 23072 4128 23078 4140
rect 24578 4128 24584 4140
rect 23072 4100 24584 4128
rect 23072 4088 23078 4100
rect 24578 4088 24584 4100
rect 24636 4088 24642 4140
rect 24762 4088 24768 4140
rect 24820 4128 24826 4140
rect 24857 4131 24915 4137
rect 24857 4128 24869 4131
rect 24820 4100 24869 4128
rect 24820 4088 24826 4100
rect 24857 4097 24869 4100
rect 24903 4097 24915 4131
rect 24857 4091 24915 4097
rect 25317 4131 25375 4137
rect 25317 4097 25329 4131
rect 25363 4128 25375 4131
rect 26326 4128 26332 4140
rect 25363 4100 26332 4128
rect 25363 4097 25375 4100
rect 25317 4091 25375 4097
rect 26326 4088 26332 4100
rect 26384 4088 26390 4140
rect 22465 4063 22523 4069
rect 22465 4060 22477 4063
rect 22336 4032 22477 4060
rect 22336 4020 22342 4032
rect 22465 4029 22477 4032
rect 22511 4029 22523 4063
rect 22465 4023 22523 4029
rect 23750 4020 23756 4072
rect 23808 4060 23814 4072
rect 23808 4032 25544 4060
rect 23808 4020 23814 4032
rect 20496 3964 20668 3992
rect 21177 3995 21235 4001
rect 20496 3952 20502 3964
rect 21177 3961 21189 3995
rect 21223 3992 21235 3995
rect 24397 3995 24455 4001
rect 21223 3964 22094 3992
rect 21223 3961 21235 3964
rect 21177 3955 21235 3961
rect 16448 3896 19104 3924
rect 19797 3927 19855 3933
rect 16448 3884 16454 3896
rect 19797 3893 19809 3927
rect 19843 3924 19855 3927
rect 20254 3924 20260 3936
rect 19843 3896 20260 3924
rect 19843 3893 19855 3896
rect 19797 3887 19855 3893
rect 20254 3884 20260 3896
rect 20312 3884 20318 3936
rect 20530 3884 20536 3936
rect 20588 3924 20594 3936
rect 21821 3927 21879 3933
rect 21821 3924 21833 3927
rect 20588 3896 21833 3924
rect 20588 3884 20594 3896
rect 21821 3893 21833 3896
rect 21867 3893 21879 3927
rect 22066 3924 22094 3964
rect 24397 3961 24409 3995
rect 24443 3992 24455 3995
rect 24854 3992 24860 4004
rect 24443 3964 24860 3992
rect 24443 3961 24455 3964
rect 24397 3955 24455 3961
rect 24854 3952 24860 3964
rect 24912 3952 24918 4004
rect 25516 4001 25544 4032
rect 25501 3995 25559 4001
rect 25501 3961 25513 3995
rect 25547 3961 25559 3995
rect 25501 3955 25559 3961
rect 27341 3995 27399 4001
rect 27341 3961 27353 3995
rect 27387 3992 27399 3995
rect 27522 3992 27528 4004
rect 27387 3964 27528 3992
rect 27387 3961 27399 3964
rect 27341 3955 27399 3961
rect 27522 3952 27528 3964
rect 27580 3952 27586 4004
rect 25406 3924 25412 3936
rect 22066 3896 25412 3924
rect 21821 3887 21879 3893
rect 25406 3884 25412 3896
rect 25464 3884 25470 3936
rect 25866 3884 25872 3936
rect 25924 3924 25930 3936
rect 27157 3927 27215 3933
rect 27157 3924 27169 3927
rect 25924 3896 27169 3924
rect 25924 3884 25930 3896
rect 27157 3893 27169 3896
rect 27203 3893 27215 3927
rect 27157 3887 27215 3893
rect 1104 3834 28060 3856
rect 1104 3782 5442 3834
rect 5494 3782 5506 3834
rect 5558 3782 5570 3834
rect 5622 3782 5634 3834
rect 5686 3782 5698 3834
rect 5750 3782 14428 3834
rect 14480 3782 14492 3834
rect 14544 3782 14556 3834
rect 14608 3782 14620 3834
rect 14672 3782 14684 3834
rect 14736 3782 23413 3834
rect 23465 3782 23477 3834
rect 23529 3782 23541 3834
rect 23593 3782 23605 3834
rect 23657 3782 23669 3834
rect 23721 3782 28060 3834
rect 1104 3760 28060 3782
rect 2409 3723 2467 3729
rect 2409 3689 2421 3723
rect 2455 3720 2467 3723
rect 2958 3720 2964 3732
rect 2455 3692 2964 3720
rect 2455 3689 2467 3692
rect 2409 3683 2467 3689
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3234 3680 3240 3732
rect 3292 3720 3298 3732
rect 4338 3720 4344 3732
rect 3292 3692 4344 3720
rect 3292 3680 3298 3692
rect 4338 3680 4344 3692
rect 4396 3680 4402 3732
rect 4430 3680 4436 3732
rect 4488 3720 4494 3732
rect 6914 3720 6920 3732
rect 4488 3692 6920 3720
rect 4488 3680 4494 3692
rect 6914 3680 6920 3692
rect 6972 3680 6978 3732
rect 7282 3720 7288 3732
rect 7243 3692 7288 3720
rect 7282 3680 7288 3692
rect 7340 3680 7346 3732
rect 7466 3720 7472 3732
rect 7427 3692 7472 3720
rect 7466 3680 7472 3692
rect 7524 3680 7530 3732
rect 7742 3680 7748 3732
rect 7800 3720 7806 3732
rect 10137 3723 10195 3729
rect 10137 3720 10149 3723
rect 7800 3692 10149 3720
rect 7800 3680 7806 3692
rect 10137 3689 10149 3692
rect 10183 3689 10195 3723
rect 10962 3720 10968 3732
rect 10137 3683 10195 3689
rect 10244 3692 10968 3720
rect 3053 3655 3111 3661
rect 3053 3621 3065 3655
rect 3099 3652 3111 3655
rect 8478 3652 8484 3664
rect 3099 3624 8484 3652
rect 3099 3621 3111 3624
rect 3053 3615 3111 3621
rect 8478 3612 8484 3624
rect 8536 3612 8542 3664
rect 8754 3612 8760 3664
rect 8812 3652 8818 3664
rect 8812 3624 9904 3652
rect 8812 3612 8818 3624
rect 1210 3544 1216 3596
rect 1268 3584 1274 3596
rect 2958 3584 2964 3596
rect 1268 3556 2964 3584
rect 1268 3544 1274 3556
rect 2958 3544 2964 3556
rect 3016 3544 3022 3596
rect 4798 3584 4804 3596
rect 3160 3556 3832 3584
rect 1949 3519 2007 3525
rect 1949 3485 1961 3519
rect 1995 3485 2007 3519
rect 1949 3479 2007 3485
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3516 2651 3519
rect 2774 3516 2780 3528
rect 2639 3488 2780 3516
rect 2639 3485 2651 3488
rect 2593 3479 2651 3485
rect 1964 3448 1992 3479
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 3160 3448 3188 3556
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3485 3295 3519
rect 3237 3479 3295 3485
rect 1964 3420 3188 3448
rect 3252 3448 3280 3479
rect 3694 3448 3700 3460
rect 3252 3420 3700 3448
rect 3694 3408 3700 3420
rect 3752 3408 3758 3460
rect 3804 3448 3832 3556
rect 4724 3556 4804 3584
rect 4246 3516 4252 3528
rect 4207 3488 4252 3516
rect 4246 3476 4252 3488
rect 4304 3476 4310 3528
rect 4724 3525 4752 3556
rect 4798 3544 4804 3556
rect 4856 3544 4862 3596
rect 5534 3584 5540 3596
rect 5447 3556 5540 3584
rect 5534 3544 5540 3556
rect 5592 3584 5598 3596
rect 7834 3584 7840 3596
rect 5592 3556 7840 3584
rect 5592 3544 5598 3556
rect 7834 3544 7840 3556
rect 7892 3584 7898 3596
rect 7929 3587 7987 3593
rect 7929 3584 7941 3587
rect 7892 3556 7941 3584
rect 7892 3544 7898 3556
rect 7929 3553 7941 3556
rect 7975 3553 7987 3587
rect 7929 3547 7987 3553
rect 8018 3544 8024 3596
rect 8076 3584 8082 3596
rect 8076 3556 9168 3584
rect 8076 3544 8082 3556
rect 4709 3519 4767 3525
rect 4709 3485 4721 3519
rect 4755 3485 4767 3519
rect 4709 3479 4767 3485
rect 4890 3476 4896 3528
rect 4948 3518 4954 3528
rect 5721 3519 5779 3525
rect 4948 3490 4991 3518
rect 4948 3476 4954 3490
rect 5721 3485 5733 3519
rect 5767 3516 5779 3519
rect 5810 3516 5816 3528
rect 5767 3488 5816 3516
rect 5767 3485 5779 3488
rect 5721 3479 5779 3485
rect 5810 3476 5816 3488
rect 5868 3476 5874 3528
rect 6549 3519 6607 3525
rect 6549 3485 6561 3519
rect 6595 3516 6607 3519
rect 6914 3516 6920 3528
rect 6595 3488 6920 3516
rect 6595 3485 6607 3488
rect 6549 3479 6607 3485
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 7193 3519 7251 3525
rect 7193 3485 7205 3519
rect 7239 3485 7251 3519
rect 7193 3479 7251 3485
rect 5077 3451 5135 3457
rect 5077 3448 5089 3451
rect 3804 3420 4844 3448
rect 1762 3380 1768 3392
rect 1723 3352 1768 3380
rect 1762 3340 1768 3352
rect 1820 3340 1826 3392
rect 2498 3340 2504 3392
rect 2556 3380 2562 3392
rect 2866 3380 2872 3392
rect 2556 3352 2872 3380
rect 2556 3340 2562 3352
rect 2866 3340 2872 3352
rect 2924 3340 2930 3392
rect 2958 3340 2964 3392
rect 3016 3380 3022 3392
rect 3418 3380 3424 3392
rect 3016 3352 3424 3380
rect 3016 3340 3022 3352
rect 3418 3340 3424 3352
rect 3476 3340 3482 3392
rect 3970 3340 3976 3392
rect 4028 3380 4034 3392
rect 4065 3383 4123 3389
rect 4065 3380 4077 3383
rect 4028 3352 4077 3380
rect 4028 3340 4034 3352
rect 4065 3349 4077 3352
rect 4111 3349 4123 3383
rect 4816 3380 4844 3420
rect 5000 3420 5089 3448
rect 5000 3380 5028 3420
rect 5077 3417 5089 3420
rect 5123 3417 5135 3451
rect 5077 3411 5135 3417
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 5316 3420 6592 3448
rect 5316 3408 5322 3420
rect 5902 3380 5908 3392
rect 4816 3352 5028 3380
rect 5863 3352 5908 3380
rect 4065 3343 4123 3349
rect 5902 3340 5908 3352
rect 5960 3340 5966 3392
rect 6365 3383 6423 3389
rect 6365 3349 6377 3383
rect 6411 3380 6423 3383
rect 6454 3380 6460 3392
rect 6411 3352 6460 3380
rect 6411 3349 6423 3352
rect 6365 3343 6423 3349
rect 6454 3340 6460 3352
rect 6512 3340 6518 3392
rect 6564 3380 6592 3420
rect 6730 3408 6736 3460
rect 6788 3448 6794 3460
rect 7009 3451 7067 3457
rect 7009 3448 7021 3451
rect 6788 3420 7021 3448
rect 6788 3408 6794 3420
rect 7009 3417 7021 3420
rect 7055 3417 7067 3451
rect 7208 3448 7236 3479
rect 7282 3476 7288 3528
rect 7340 3516 7346 3528
rect 9140 3525 9168 3556
rect 8113 3519 8171 3525
rect 7340 3488 7385 3516
rect 7340 3476 7346 3488
rect 8113 3485 8125 3519
rect 8159 3485 8171 3519
rect 8113 3479 8171 3485
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 7558 3448 7564 3460
rect 7208 3420 7564 3448
rect 7009 3411 7067 3417
rect 7558 3408 7564 3420
rect 7616 3408 7622 3460
rect 8128 3448 8156 3479
rect 9490 3476 9496 3528
rect 9548 3516 9554 3528
rect 9876 3525 9904 3624
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 10244 3652 10272 3692
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 11422 3680 11428 3732
rect 11480 3720 11486 3732
rect 15473 3723 15531 3729
rect 15473 3720 15485 3723
rect 11480 3692 15485 3720
rect 11480 3680 11486 3692
rect 15473 3689 15485 3692
rect 15519 3689 15531 3723
rect 15473 3683 15531 3689
rect 16114 3680 16120 3732
rect 16172 3720 16178 3732
rect 16485 3723 16543 3729
rect 16485 3720 16497 3723
rect 16172 3692 16497 3720
rect 16172 3680 16178 3692
rect 16485 3689 16497 3692
rect 16531 3689 16543 3723
rect 16485 3683 16543 3689
rect 17313 3723 17371 3729
rect 17313 3689 17325 3723
rect 17359 3720 17371 3723
rect 17494 3720 17500 3732
rect 17359 3692 17500 3720
rect 17359 3689 17371 3692
rect 17313 3683 17371 3689
rect 17494 3680 17500 3692
rect 17552 3680 17558 3732
rect 18601 3723 18659 3729
rect 18601 3689 18613 3723
rect 18647 3720 18659 3723
rect 20898 3720 20904 3732
rect 18647 3692 20904 3720
rect 18647 3689 18659 3692
rect 18601 3683 18659 3689
rect 20898 3680 20904 3692
rect 20956 3680 20962 3732
rect 21082 3720 21088 3732
rect 21043 3692 21088 3720
rect 21082 3680 21088 3692
rect 21140 3680 21146 3732
rect 21266 3720 21272 3732
rect 21227 3692 21272 3720
rect 21266 3680 21272 3692
rect 21324 3680 21330 3732
rect 23106 3720 23112 3732
rect 21376 3692 23112 3720
rect 10008 3624 10272 3652
rect 11977 3655 12035 3661
rect 10008 3612 10014 3624
rect 11977 3621 11989 3655
rect 12023 3652 12035 3655
rect 12802 3652 12808 3664
rect 12023 3624 12434 3652
rect 12763 3624 12808 3652
rect 12023 3621 12035 3624
rect 11977 3615 12035 3621
rect 11606 3544 11612 3596
rect 11664 3544 11670 3596
rect 12406 3584 12434 3624
rect 12802 3612 12808 3624
rect 12860 3612 12866 3664
rect 15102 3612 15108 3664
rect 15160 3652 15166 3664
rect 17034 3652 17040 3664
rect 15160 3624 17040 3652
rect 15160 3612 15166 3624
rect 17034 3612 17040 3624
rect 17092 3612 17098 3664
rect 17126 3612 17132 3664
rect 17184 3652 17190 3664
rect 17954 3652 17960 3664
rect 17184 3624 17960 3652
rect 17184 3612 17190 3624
rect 17954 3612 17960 3624
rect 18012 3612 18018 3664
rect 20441 3655 20499 3661
rect 19260 3624 20116 3652
rect 16117 3587 16175 3593
rect 12406 3556 12664 3584
rect 9585 3519 9643 3525
rect 9585 3516 9597 3519
rect 9548 3488 9597 3516
rect 9548 3476 9554 3488
rect 9585 3485 9597 3488
rect 9631 3485 9643 3519
rect 9585 3479 9643 3485
rect 9861 3519 9919 3525
rect 9861 3485 9873 3519
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 9953 3519 10011 3525
rect 9953 3485 9965 3519
rect 9999 3516 10011 3519
rect 10594 3516 10600 3528
rect 9999 3488 10600 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 10594 3476 10600 3488
rect 10652 3476 10658 3528
rect 10965 3519 11023 3525
rect 10965 3485 10977 3519
rect 11011 3516 11023 3519
rect 11330 3516 11336 3528
rect 11011 3488 11336 3516
rect 11011 3485 11023 3488
rect 10965 3479 11023 3485
rect 11330 3476 11336 3488
rect 11388 3476 11394 3528
rect 11422 3476 11428 3528
rect 11480 3516 11486 3528
rect 11624 3516 11652 3544
rect 11701 3519 11759 3525
rect 11701 3516 11713 3519
rect 11480 3488 11525 3516
rect 11624 3488 11713 3516
rect 11480 3476 11486 3488
rect 11701 3485 11713 3488
rect 11747 3485 11759 3519
rect 11701 3479 11759 3485
rect 11793 3519 11851 3525
rect 11793 3485 11805 3519
rect 11839 3516 11851 3519
rect 11882 3516 11888 3528
rect 11839 3488 11888 3516
rect 11839 3485 11851 3488
rect 11793 3479 11851 3485
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 12434 3476 12440 3528
rect 12492 3516 12498 3528
rect 12636 3525 12664 3556
rect 16117 3553 16129 3587
rect 16163 3584 16175 3587
rect 16945 3587 17003 3593
rect 16945 3584 16957 3587
rect 16163 3556 16957 3584
rect 16163 3553 16175 3556
rect 16117 3547 16175 3553
rect 16945 3553 16957 3556
rect 16991 3584 17003 3587
rect 18138 3584 18144 3596
rect 16991 3556 18144 3584
rect 16991 3553 17003 3556
rect 16945 3547 17003 3553
rect 18138 3544 18144 3556
rect 18196 3544 18202 3596
rect 18233 3587 18291 3593
rect 18233 3553 18245 3587
rect 18279 3584 18291 3587
rect 18598 3584 18604 3596
rect 18279 3556 18604 3584
rect 18279 3553 18291 3556
rect 18233 3547 18291 3553
rect 18598 3544 18604 3556
rect 18656 3584 18662 3596
rect 19260 3584 19288 3624
rect 20088 3593 20116 3624
rect 20441 3621 20453 3655
rect 20487 3652 20499 3655
rect 21376 3652 21404 3692
rect 23106 3680 23112 3692
rect 23164 3680 23170 3732
rect 25866 3680 25872 3732
rect 25924 3720 25930 3732
rect 26142 3720 26148 3732
rect 25924 3692 26148 3720
rect 25924 3680 25930 3692
rect 26142 3680 26148 3692
rect 26200 3720 26206 3732
rect 26973 3723 27031 3729
rect 26973 3720 26985 3723
rect 26200 3692 26985 3720
rect 26200 3680 26206 3692
rect 26973 3689 26985 3692
rect 27019 3689 27031 3723
rect 26973 3683 27031 3689
rect 20487 3624 21404 3652
rect 20487 3621 20499 3624
rect 20441 3615 20499 3621
rect 21450 3612 21456 3664
rect 21508 3652 21514 3664
rect 25317 3655 25375 3661
rect 25317 3652 25329 3655
rect 21508 3624 25329 3652
rect 21508 3612 21514 3624
rect 25317 3621 25329 3624
rect 25363 3621 25375 3655
rect 25317 3615 25375 3621
rect 25590 3612 25596 3664
rect 25648 3652 25654 3664
rect 26329 3655 26387 3661
rect 26329 3652 26341 3655
rect 25648 3624 26341 3652
rect 25648 3612 25654 3624
rect 26329 3621 26341 3624
rect 26375 3621 26387 3655
rect 26329 3615 26387 3621
rect 26602 3612 26608 3664
rect 26660 3652 26666 3664
rect 27157 3655 27215 3661
rect 27157 3652 27169 3655
rect 26660 3624 27169 3652
rect 26660 3612 26666 3624
rect 27157 3621 27169 3624
rect 27203 3621 27215 3655
rect 27157 3615 27215 3621
rect 18656 3556 19288 3584
rect 18656 3544 18662 3556
rect 12621 3519 12679 3525
rect 12492 3488 12537 3516
rect 12492 3476 12498 3488
rect 12621 3485 12633 3519
rect 12667 3485 12679 3519
rect 13262 3516 13268 3528
rect 13223 3488 13268 3516
rect 12621 3479 12679 3485
rect 13262 3476 13268 3488
rect 13320 3476 13326 3528
rect 14093 3519 14151 3525
rect 14093 3485 14105 3519
rect 14139 3516 14151 3519
rect 14182 3516 14188 3528
rect 14139 3488 14188 3516
rect 14139 3485 14151 3488
rect 14093 3479 14151 3485
rect 14182 3476 14188 3488
rect 14240 3476 14246 3528
rect 14366 3525 14372 3528
rect 14360 3479 14372 3525
rect 14424 3516 14430 3528
rect 16301 3519 16359 3525
rect 14424 3488 14460 3516
rect 14366 3476 14372 3479
rect 14424 3476 14430 3488
rect 16301 3485 16313 3519
rect 16347 3516 16359 3519
rect 16482 3516 16488 3528
rect 16347 3488 16488 3516
rect 16347 3485 16359 3488
rect 16301 3479 16359 3485
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 17129 3519 17187 3525
rect 17129 3485 17141 3519
rect 17175 3516 17187 3519
rect 17402 3516 17408 3528
rect 17175 3488 17408 3516
rect 17175 3485 17187 3488
rect 17129 3479 17187 3485
rect 17402 3476 17408 3488
rect 17460 3476 17466 3528
rect 18417 3519 18475 3525
rect 18417 3485 18429 3519
rect 18463 3516 18475 3519
rect 18690 3516 18696 3528
rect 18463 3488 18696 3516
rect 18463 3485 18475 3488
rect 18417 3479 18475 3485
rect 18690 3476 18696 3488
rect 18748 3476 18754 3528
rect 19260 3525 19288 3556
rect 19613 3587 19671 3593
rect 19613 3553 19625 3587
rect 19659 3584 19671 3587
rect 20073 3587 20131 3593
rect 19659 3556 19840 3584
rect 19659 3553 19671 3556
rect 19613 3547 19671 3553
rect 19245 3519 19303 3525
rect 19245 3485 19257 3519
rect 19291 3485 19303 3519
rect 19245 3479 19303 3485
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 19484 3488 19529 3516
rect 19484 3476 19490 3488
rect 9674 3448 9680 3460
rect 8128 3420 9680 3448
rect 9674 3408 9680 3420
rect 9732 3408 9738 3460
rect 9769 3451 9827 3457
rect 9769 3417 9781 3451
rect 9815 3448 9827 3451
rect 10870 3448 10876 3460
rect 9815 3420 10876 3448
rect 9815 3417 9827 3420
rect 9769 3411 9827 3417
rect 10870 3408 10876 3420
rect 10928 3448 10934 3460
rect 11609 3451 11667 3457
rect 11609 3448 11621 3451
rect 10928 3420 11621 3448
rect 10928 3408 10934 3420
rect 11609 3417 11621 3420
rect 11655 3417 11667 3451
rect 11609 3411 11667 3417
rect 11974 3408 11980 3460
rect 12032 3448 12038 3460
rect 12032 3420 13492 3448
rect 12032 3408 12038 3420
rect 8297 3383 8355 3389
rect 8297 3380 8309 3383
rect 6564 3352 8309 3380
rect 8297 3349 8309 3352
rect 8343 3349 8355 3383
rect 8297 3343 8355 3349
rect 8386 3340 8392 3392
rect 8444 3380 8450 3392
rect 8941 3383 8999 3389
rect 8941 3380 8953 3383
rect 8444 3352 8953 3380
rect 8444 3340 8450 3352
rect 8941 3349 8953 3352
rect 8987 3349 8999 3383
rect 8941 3343 8999 3349
rect 10781 3383 10839 3389
rect 10781 3349 10793 3383
rect 10827 3380 10839 3383
rect 11882 3380 11888 3392
rect 10827 3352 11888 3380
rect 10827 3349 10839 3352
rect 10781 3343 10839 3349
rect 11882 3340 11888 3352
rect 11940 3340 11946 3392
rect 13464 3389 13492 3420
rect 15010 3408 15016 3460
rect 15068 3448 15074 3460
rect 19334 3448 19340 3460
rect 15068 3420 19340 3448
rect 15068 3408 15074 3420
rect 19334 3408 19340 3420
rect 19392 3408 19398 3460
rect 19812 3448 19840 3556
rect 20073 3553 20085 3587
rect 20119 3553 20131 3587
rect 20073 3547 20131 3553
rect 20840 3556 25544 3584
rect 20254 3516 20260 3528
rect 20215 3488 20260 3516
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 20840 3448 20868 3556
rect 21726 3516 21732 3528
rect 21687 3488 21732 3516
rect 21726 3476 21732 3488
rect 21784 3476 21790 3528
rect 22005 3519 22063 3525
rect 22005 3485 22017 3519
rect 22051 3516 22063 3519
rect 22051 3488 23060 3516
rect 22051 3485 22063 3488
rect 22005 3479 22063 3485
rect 19812 3420 20868 3448
rect 20901 3451 20959 3457
rect 20901 3417 20913 3451
rect 20947 3448 20959 3451
rect 22462 3448 22468 3460
rect 20947 3420 22468 3448
rect 20947 3417 20959 3420
rect 20901 3411 20959 3417
rect 22462 3408 22468 3420
rect 22520 3408 22526 3460
rect 23032 3448 23060 3488
rect 23106 3476 23112 3528
rect 23164 3516 23170 3528
rect 23201 3519 23259 3525
rect 23201 3516 23213 3519
rect 23164 3488 23213 3516
rect 23164 3476 23170 3488
rect 23201 3485 23213 3488
rect 23247 3485 23259 3519
rect 23201 3479 23259 3485
rect 23290 3476 23296 3528
rect 23348 3516 23354 3528
rect 23477 3519 23535 3525
rect 23477 3516 23489 3519
rect 23348 3488 23489 3516
rect 23348 3476 23354 3488
rect 23477 3485 23489 3488
rect 23523 3485 23535 3519
rect 24578 3516 24584 3528
rect 24539 3488 24584 3516
rect 23477 3479 23535 3485
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 24762 3476 24768 3528
rect 24820 3516 24826 3528
rect 25516 3525 25544 3556
rect 24857 3519 24915 3525
rect 24857 3516 24869 3519
rect 24820 3488 24869 3516
rect 24820 3476 24826 3488
rect 24857 3485 24869 3488
rect 24903 3485 24915 3519
rect 24857 3479 24915 3485
rect 25501 3519 25559 3525
rect 25501 3485 25513 3519
rect 25547 3485 25559 3519
rect 25501 3479 25559 3485
rect 23308 3448 23336 3476
rect 24872 3448 24900 3479
rect 27154 3476 27160 3528
rect 27212 3516 27218 3528
rect 28718 3516 28724 3528
rect 27212 3488 28724 3516
rect 27212 3476 27218 3488
rect 28718 3476 28724 3488
rect 28776 3476 28782 3528
rect 25958 3448 25964 3460
rect 23032 3420 24900 3448
rect 25919 3420 25964 3448
rect 25958 3408 25964 3420
rect 26016 3408 26022 3460
rect 26418 3408 26424 3460
rect 26476 3448 26482 3460
rect 26789 3451 26847 3457
rect 26789 3448 26801 3451
rect 26476 3420 26801 3448
rect 26476 3408 26482 3420
rect 26789 3417 26801 3420
rect 26835 3417 26847 3451
rect 26789 3411 26847 3417
rect 13449 3383 13507 3389
rect 13449 3349 13461 3383
rect 13495 3349 13507 3383
rect 13449 3343 13507 3349
rect 13538 3340 13544 3392
rect 13596 3380 13602 3392
rect 15838 3380 15844 3392
rect 13596 3352 15844 3380
rect 13596 3340 13602 3352
rect 15838 3340 15844 3352
rect 15896 3340 15902 3392
rect 16482 3340 16488 3392
rect 16540 3380 16546 3392
rect 17954 3380 17960 3392
rect 16540 3352 17960 3380
rect 16540 3340 16546 3352
rect 17954 3340 17960 3352
rect 18012 3340 18018 3392
rect 18782 3340 18788 3392
rect 18840 3380 18846 3392
rect 20254 3380 20260 3392
rect 18840 3352 20260 3380
rect 18840 3340 18846 3352
rect 20254 3340 20260 3352
rect 20312 3340 20318 3392
rect 20990 3340 20996 3392
rect 21048 3380 21054 3392
rect 21101 3383 21159 3389
rect 21101 3380 21113 3383
rect 21048 3352 21113 3380
rect 21048 3340 21054 3352
rect 21101 3349 21113 3352
rect 21147 3349 21159 3383
rect 21101 3343 21159 3349
rect 22370 3340 22376 3392
rect 22428 3380 22434 3392
rect 23017 3383 23075 3389
rect 23017 3380 23029 3383
rect 22428 3352 23029 3380
rect 22428 3340 22434 3352
rect 23017 3349 23029 3352
rect 23063 3349 23075 3383
rect 23017 3343 23075 3349
rect 23290 3340 23296 3392
rect 23348 3380 23354 3392
rect 23385 3383 23443 3389
rect 23385 3380 23397 3383
rect 23348 3352 23397 3380
rect 23348 3340 23354 3352
rect 23385 3349 23397 3352
rect 23431 3349 23443 3383
rect 24394 3380 24400 3392
rect 24355 3352 24400 3380
rect 23385 3343 23443 3349
rect 24394 3340 24400 3352
rect 24452 3340 24458 3392
rect 24762 3380 24768 3392
rect 24723 3352 24768 3380
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 25314 3340 25320 3392
rect 25372 3380 25378 3392
rect 26161 3383 26219 3389
rect 26161 3380 26173 3383
rect 25372 3352 26173 3380
rect 25372 3340 25378 3352
rect 26161 3349 26173 3352
rect 26207 3380 26219 3383
rect 26878 3380 26884 3392
rect 26207 3352 26884 3380
rect 26207 3349 26219 3352
rect 26161 3343 26219 3349
rect 26878 3340 26884 3352
rect 26936 3380 26942 3392
rect 26989 3383 27047 3389
rect 26989 3380 27001 3383
rect 26936 3352 27001 3380
rect 26936 3340 26942 3352
rect 26989 3349 27001 3352
rect 27035 3349 27047 3383
rect 26989 3343 27047 3349
rect 1104 3290 28060 3312
rect 1104 3238 9935 3290
rect 9987 3238 9999 3290
rect 10051 3238 10063 3290
rect 10115 3238 10127 3290
rect 10179 3238 10191 3290
rect 10243 3238 18920 3290
rect 18972 3238 18984 3290
rect 19036 3238 19048 3290
rect 19100 3238 19112 3290
rect 19164 3238 19176 3290
rect 19228 3238 28060 3290
rect 1104 3216 28060 3238
rect 4798 3136 4804 3188
rect 4856 3176 4862 3188
rect 5534 3176 5540 3188
rect 4856 3148 5540 3176
rect 4856 3136 4862 3148
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 6178 3136 6184 3188
rect 6236 3176 6242 3188
rect 6236 3148 6776 3176
rect 6236 3136 6242 3148
rect 2682 3108 2688 3120
rect 1504 3080 2688 3108
rect 1504 3049 1532 3080
rect 2682 3068 2688 3080
rect 2740 3108 2746 3120
rect 5074 3108 5080 3120
rect 2740 3080 5080 3108
rect 2740 3068 2746 3080
rect 1762 3049 1768 3052
rect 1489 3043 1547 3049
rect 1489 3009 1501 3043
rect 1535 3009 1547 3043
rect 1756 3040 1768 3049
rect 1723 3012 1768 3040
rect 1489 3003 1547 3009
rect 1756 3003 1768 3012
rect 1762 3000 1768 3003
rect 1820 3000 1826 3052
rect 2314 3000 2320 3052
rect 2372 3040 2378 3052
rect 3234 3040 3240 3052
rect 2372 3012 3240 3040
rect 2372 3000 2378 3012
rect 3234 3000 3240 3012
rect 3292 3000 3298 3052
rect 3344 3049 3372 3080
rect 5074 3068 5080 3080
rect 5132 3068 5138 3120
rect 5258 3068 5264 3120
rect 5316 3108 5322 3120
rect 5353 3111 5411 3117
rect 5353 3108 5365 3111
rect 5316 3080 5365 3108
rect 5316 3068 5322 3080
rect 5353 3077 5365 3080
rect 5399 3077 5411 3111
rect 5353 3071 5411 3077
rect 5442 3068 5448 3120
rect 5500 3108 5506 3120
rect 5500 3080 5545 3108
rect 5500 3068 5506 3080
rect 3602 3049 3608 3052
rect 3329 3043 3387 3049
rect 3329 3009 3341 3043
rect 3375 3009 3387 3043
rect 3329 3003 3387 3009
rect 3596 3003 3608 3049
rect 3660 3040 3666 3052
rect 4614 3040 4620 3052
rect 3660 3012 3696 3040
rect 4347 3012 4620 3040
rect 3602 3000 3608 3003
rect 3660 3000 3666 3012
rect 2590 2864 2596 2916
rect 2648 2904 2654 2916
rect 3326 2904 3332 2916
rect 2648 2876 3332 2904
rect 2648 2864 2654 2876
rect 3326 2864 3332 2876
rect 3384 2864 3390 2916
rect 2869 2839 2927 2845
rect 2869 2805 2881 2839
rect 2915 2836 2927 2839
rect 4347 2836 4375 3012
rect 4614 3000 4620 3012
rect 4672 3040 4678 3052
rect 5169 3043 5227 3049
rect 5169 3040 5181 3043
rect 4672 3012 5181 3040
rect 4672 3000 4678 3012
rect 5169 3009 5181 3012
rect 5215 3009 5227 3043
rect 5169 3003 5227 3009
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3040 5595 3043
rect 6270 3040 6276 3052
rect 5583 3012 6276 3040
rect 5583 3009 5595 3012
rect 5537 3003 5595 3009
rect 6270 3000 6276 3012
rect 6328 3000 6334 3052
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 5074 2932 5080 2984
rect 5132 2972 5138 2984
rect 6380 2972 6408 3003
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 6621 3043 6679 3049
rect 6621 3040 6633 3043
rect 6512 3012 6633 3040
rect 6512 3000 6518 3012
rect 6621 3009 6633 3012
rect 6667 3009 6679 3043
rect 6748 3040 6776 3148
rect 6914 3136 6920 3188
rect 6972 3176 6978 3188
rect 7190 3176 7196 3188
rect 6972 3148 7196 3176
rect 6972 3136 6978 3148
rect 7190 3136 7196 3148
rect 7248 3136 7254 3188
rect 7282 3136 7288 3188
rect 7340 3176 7346 3188
rect 9585 3179 9643 3185
rect 9585 3176 9597 3179
rect 7340 3148 9597 3176
rect 7340 3136 7346 3148
rect 9585 3145 9597 3148
rect 9631 3145 9643 3179
rect 9585 3139 9643 3145
rect 7374 3068 7380 3120
rect 7432 3108 7438 3120
rect 7926 3108 7932 3120
rect 7432 3080 7932 3108
rect 7432 3068 7438 3080
rect 7926 3068 7932 3080
rect 7984 3068 7990 3120
rect 8478 3117 8484 3120
rect 8472 3108 8484 3117
rect 8439 3080 8484 3108
rect 8472 3071 8484 3080
rect 8478 3068 8484 3071
rect 8536 3068 8542 3120
rect 8202 3040 8208 3052
rect 6748 3012 7420 3040
rect 8163 3012 8208 3040
rect 6621 3003 6679 3009
rect 5132 2944 6408 2972
rect 7392 2972 7420 3012
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 9600 3040 9628 3139
rect 9674 3136 9680 3188
rect 9732 3176 9738 3188
rect 10597 3179 10655 3185
rect 10597 3176 10609 3179
rect 9732 3148 10609 3176
rect 9732 3136 9738 3148
rect 10597 3145 10609 3148
rect 10643 3145 10655 3179
rect 10597 3139 10655 3145
rect 10870 3136 10876 3188
rect 10928 3136 10934 3188
rect 12526 3176 12532 3188
rect 11532 3148 12532 3176
rect 10229 3111 10287 3117
rect 10229 3077 10241 3111
rect 10275 3108 10287 3111
rect 10502 3108 10508 3120
rect 10275 3080 10508 3108
rect 10275 3077 10287 3080
rect 10229 3071 10287 3077
rect 10502 3068 10508 3080
rect 10560 3108 10566 3120
rect 10888 3108 10916 3136
rect 10560 3080 10916 3108
rect 10560 3068 10566 3080
rect 10045 3043 10103 3049
rect 10045 3040 10057 3043
rect 8312 3012 9260 3040
rect 9600 3012 10057 3040
rect 8312 2972 8340 3012
rect 7392 2944 8340 2972
rect 9232 2972 9260 3012
rect 10045 3009 10057 3012
rect 10091 3009 10103 3043
rect 10045 3003 10103 3009
rect 10321 3043 10379 3049
rect 10321 3009 10333 3043
rect 10367 3009 10379 3043
rect 10321 3003 10379 3009
rect 10413 3043 10471 3049
rect 10413 3009 10425 3043
rect 10459 3040 10471 3043
rect 10594 3040 10600 3052
rect 10459 3012 10600 3040
rect 10459 3009 10471 3012
rect 10413 3003 10471 3009
rect 10336 2972 10364 3003
rect 10594 3000 10600 3012
rect 10652 3000 10658 3052
rect 11532 3049 11560 3148
rect 12526 3136 12532 3148
rect 12584 3136 12590 3188
rect 13262 3136 13268 3188
rect 13320 3176 13326 3188
rect 14185 3179 14243 3185
rect 14185 3176 14197 3179
rect 13320 3148 14197 3176
rect 13320 3136 13326 3148
rect 14185 3145 14197 3148
rect 14231 3145 14243 3179
rect 14185 3139 14243 3145
rect 14274 3136 14280 3188
rect 14332 3176 14338 3188
rect 15102 3176 15108 3188
rect 14332 3148 15108 3176
rect 14332 3136 14338 3148
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 15197 3179 15255 3185
rect 15197 3145 15209 3179
rect 15243 3176 15255 3179
rect 15286 3176 15292 3188
rect 15243 3148 15292 3176
rect 15243 3145 15255 3148
rect 15197 3139 15255 3145
rect 15286 3136 15292 3148
rect 15344 3136 15350 3188
rect 16942 3176 16948 3188
rect 15764 3148 16948 3176
rect 12250 3108 12256 3120
rect 11624 3080 12256 3108
rect 11517 3043 11575 3049
rect 11517 3009 11529 3043
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 9232 2944 10364 2972
rect 5132 2932 5138 2944
rect 10686 2932 10692 2984
rect 10744 2972 10750 2984
rect 11624 2972 11652 3080
rect 12250 3068 12256 3080
rect 12308 3068 12314 3120
rect 12618 3068 12624 3120
rect 12676 3108 12682 3120
rect 15470 3108 15476 3120
rect 12676 3080 15476 3108
rect 12676 3068 12682 3080
rect 15470 3068 15476 3080
rect 15528 3068 15534 3120
rect 11784 3043 11842 3049
rect 11784 3009 11796 3043
rect 11830 3040 11842 3043
rect 12066 3040 12072 3052
rect 11830 3012 12072 3040
rect 11830 3009 11842 3012
rect 11784 3003 11842 3009
rect 12066 3000 12072 3012
rect 12124 3000 12130 3052
rect 13078 3000 13084 3052
rect 13136 3040 13142 3052
rect 13541 3043 13599 3049
rect 13541 3040 13553 3043
rect 13136 3012 13553 3040
rect 13136 3000 13142 3012
rect 13541 3009 13553 3012
rect 13587 3009 13599 3043
rect 13541 3003 13599 3009
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3040 13783 3043
rect 14369 3043 14427 3049
rect 14369 3040 14381 3043
rect 13771 3012 14381 3040
rect 13771 3009 13783 3012
rect 13725 3003 13783 3009
rect 14369 3009 14381 3012
rect 14415 3009 14427 3043
rect 14369 3003 14427 3009
rect 15013 3043 15071 3049
rect 15013 3009 15025 3043
rect 15059 3040 15071 3043
rect 15764 3040 15792 3148
rect 16942 3136 16948 3148
rect 17000 3136 17006 3188
rect 18138 3136 18144 3188
rect 18196 3176 18202 3188
rect 18414 3176 18420 3188
rect 18196 3148 18420 3176
rect 18196 3136 18202 3148
rect 18414 3136 18420 3148
rect 18472 3136 18478 3188
rect 18693 3179 18751 3185
rect 18693 3145 18705 3179
rect 18739 3176 18751 3179
rect 20070 3176 20076 3188
rect 18739 3148 20076 3176
rect 18739 3145 18751 3148
rect 18693 3139 18751 3145
rect 20070 3136 20076 3148
rect 20128 3136 20134 3188
rect 20180 3148 21588 3176
rect 16666 3068 16672 3120
rect 16724 3108 16730 3120
rect 20180 3108 20208 3148
rect 20622 3108 20628 3120
rect 16724 3080 20208 3108
rect 20583 3080 20628 3108
rect 16724 3068 16730 3080
rect 20622 3068 20628 3080
rect 20680 3068 20686 3120
rect 20841 3111 20899 3117
rect 20841 3077 20853 3111
rect 20887 3108 20899 3111
rect 20990 3108 20996 3120
rect 20887 3080 20996 3108
rect 20887 3077 20899 3080
rect 20841 3071 20899 3077
rect 20990 3068 20996 3080
rect 21048 3068 21054 3120
rect 15059 3012 15792 3040
rect 15841 3043 15899 3049
rect 15059 3009 15071 3012
rect 15013 3003 15071 3009
rect 15841 3009 15853 3043
rect 15887 3040 15899 3043
rect 16482 3040 16488 3052
rect 15887 3012 16488 3040
rect 15887 3009 15899 3012
rect 15841 3003 15899 3009
rect 16482 3000 16488 3012
rect 16540 3000 16546 3052
rect 16761 3043 16819 3049
rect 16761 3009 16773 3043
rect 16807 3009 16819 3043
rect 16761 3003 16819 3009
rect 16853 3043 16911 3049
rect 16853 3009 16865 3043
rect 16899 3040 16911 3043
rect 17218 3040 17224 3052
rect 16899 3012 17224 3040
rect 16899 3009 16911 3012
rect 16853 3003 16911 3009
rect 13354 2972 13360 2984
rect 10744 2944 11652 2972
rect 13267 2944 13360 2972
rect 10744 2932 10750 2944
rect 13354 2932 13360 2944
rect 13412 2972 13418 2984
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 13412 2944 14841 2972
rect 13412 2932 13418 2944
rect 14829 2941 14841 2944
rect 14875 2972 14887 2975
rect 15657 2975 15715 2981
rect 15657 2972 15669 2975
rect 14875 2944 15669 2972
rect 14875 2941 14887 2944
rect 14829 2935 14887 2941
rect 15657 2941 15669 2944
rect 15703 2972 15715 2975
rect 15930 2972 15936 2984
rect 15703 2944 15936 2972
rect 15703 2941 15715 2944
rect 15657 2935 15715 2941
rect 15930 2932 15936 2944
rect 15988 2932 15994 2984
rect 16776 2972 16804 3003
rect 17218 3000 17224 3012
rect 17276 3000 17282 3052
rect 17681 3043 17739 3049
rect 17681 3009 17693 3043
rect 17727 3040 17739 3043
rect 18529 3043 18587 3049
rect 17727 3012 18460 3040
rect 17727 3009 17739 3012
rect 17681 3003 17739 3009
rect 17497 2975 17555 2981
rect 17497 2972 17509 2975
rect 16776 2944 17509 2972
rect 17497 2941 17509 2944
rect 17543 2972 17555 2975
rect 18138 2972 18144 2984
rect 17543 2944 18144 2972
rect 17543 2941 17555 2944
rect 17497 2935 17555 2941
rect 18138 2932 18144 2944
rect 18196 2972 18202 2984
rect 18325 2975 18383 2981
rect 18325 2972 18337 2975
rect 18196 2944 18337 2972
rect 18196 2932 18202 2944
rect 18325 2941 18337 2944
rect 18371 2941 18383 2975
rect 18432 2972 18460 3012
rect 18529 3009 18541 3043
rect 18575 3040 18587 3043
rect 18690 3040 18696 3052
rect 18575 3012 18696 3040
rect 18575 3009 18587 3012
rect 18529 3003 18587 3009
rect 18690 3000 18696 3012
rect 18748 3000 18754 3052
rect 19705 3043 19763 3049
rect 19705 3009 19717 3043
rect 19751 3040 19763 3043
rect 19978 3040 19984 3052
rect 19751 3012 19984 3040
rect 19751 3009 19763 3012
rect 19705 3003 19763 3009
rect 19978 3000 19984 3012
rect 20036 3000 20042 3052
rect 21174 3040 21180 3052
rect 20180 3012 21180 3040
rect 20180 2981 20208 3012
rect 21174 3000 21180 3012
rect 21232 3000 21238 3052
rect 20165 2975 20223 2981
rect 18432 2944 19748 2972
rect 18325 2935 18383 2941
rect 19720 2916 19748 2944
rect 20165 2941 20177 2975
rect 20211 2941 20223 2975
rect 20165 2935 20223 2941
rect 20806 2932 20812 2984
rect 20864 2972 20870 2984
rect 21450 2972 21456 2984
rect 20864 2944 21456 2972
rect 20864 2932 20870 2944
rect 21450 2932 21456 2944
rect 21508 2932 21514 2984
rect 4890 2864 4896 2916
rect 4948 2904 4954 2916
rect 5721 2907 5779 2913
rect 5721 2904 5733 2907
rect 4948 2876 5733 2904
rect 4948 2864 4954 2876
rect 5721 2873 5733 2876
rect 5767 2873 5779 2907
rect 5721 2867 5779 2873
rect 10410 2864 10416 2916
rect 10468 2904 10474 2916
rect 11238 2904 11244 2916
rect 10468 2876 11244 2904
rect 10468 2864 10474 2876
rect 11238 2864 11244 2876
rect 11296 2864 11302 2916
rect 12526 2864 12532 2916
rect 12584 2904 12590 2916
rect 15378 2904 15384 2916
rect 12584 2876 15384 2904
rect 12584 2864 12590 2876
rect 15378 2864 15384 2876
rect 15436 2864 15442 2916
rect 17037 2907 17095 2913
rect 17037 2873 17049 2907
rect 17083 2904 17095 2907
rect 19518 2904 19524 2916
rect 17083 2876 19524 2904
rect 17083 2873 17095 2876
rect 17037 2867 17095 2873
rect 19518 2864 19524 2876
rect 19576 2864 19582 2916
rect 19702 2864 19708 2916
rect 19760 2864 19766 2916
rect 20070 2904 20076 2916
rect 20031 2876 20076 2904
rect 20070 2864 20076 2876
rect 20128 2864 20134 2916
rect 20898 2904 20904 2916
rect 20811 2876 20904 2904
rect 4706 2836 4712 2848
rect 2915 2808 4375 2836
rect 4667 2808 4712 2836
rect 2915 2805 2927 2808
rect 2869 2799 2927 2805
rect 4706 2796 4712 2808
rect 4764 2796 4770 2848
rect 7006 2796 7012 2848
rect 7064 2836 7070 2848
rect 7558 2836 7564 2848
rect 7064 2808 7564 2836
rect 7064 2796 7070 2808
rect 7558 2796 7564 2808
rect 7616 2836 7622 2848
rect 7745 2839 7803 2845
rect 7745 2836 7757 2839
rect 7616 2808 7757 2836
rect 7616 2796 7622 2808
rect 7745 2805 7757 2808
rect 7791 2805 7803 2839
rect 7745 2799 7803 2805
rect 9858 2796 9864 2848
rect 9916 2836 9922 2848
rect 12897 2839 12955 2845
rect 12897 2836 12909 2839
rect 9916 2808 12909 2836
rect 9916 2796 9922 2808
rect 12897 2805 12909 2808
rect 12943 2805 12955 2839
rect 12897 2799 12955 2805
rect 13170 2796 13176 2848
rect 13228 2836 13234 2848
rect 16025 2839 16083 2845
rect 16025 2836 16037 2839
rect 13228 2808 16037 2836
rect 13228 2796 13234 2808
rect 16025 2805 16037 2808
rect 16071 2805 16083 2839
rect 16025 2799 16083 2805
rect 17865 2839 17923 2845
rect 17865 2805 17877 2839
rect 17911 2836 17923 2839
rect 20438 2836 20444 2848
rect 17911 2808 20444 2836
rect 17911 2805 17923 2808
rect 17865 2799 17923 2805
rect 20438 2796 20444 2808
rect 20496 2796 20502 2848
rect 20824 2845 20852 2876
rect 20898 2864 20904 2876
rect 20956 2904 20962 2916
rect 21082 2904 21088 2916
rect 20956 2876 21088 2904
rect 20956 2864 20962 2876
rect 21082 2864 21088 2876
rect 21140 2864 21146 2916
rect 21560 2904 21588 3148
rect 21634 3136 21640 3188
rect 21692 3176 21698 3188
rect 21692 3148 24716 3176
rect 21692 3136 21698 3148
rect 24394 3117 24400 3120
rect 24388 3108 24400 3117
rect 22112 3080 24164 3108
rect 24355 3080 24400 3108
rect 22112 3052 22140 3080
rect 22094 3000 22100 3052
rect 22152 3040 22158 3052
rect 22370 3049 22376 3052
rect 22364 3040 22376 3049
rect 22152 3012 22197 3040
rect 22331 3012 22376 3040
rect 22152 3000 22158 3012
rect 22364 3003 22376 3012
rect 22370 3000 22376 3003
rect 22428 3000 22434 3052
rect 23106 3000 23112 3052
rect 23164 3040 23170 3052
rect 23750 3040 23756 3052
rect 23164 3012 23756 3040
rect 23164 3000 23170 3012
rect 23750 3000 23756 3012
rect 23808 3000 23814 3052
rect 24136 3049 24164 3080
rect 24388 3071 24400 3080
rect 24394 3068 24400 3071
rect 24452 3068 24458 3120
rect 24121 3043 24179 3049
rect 24121 3009 24133 3043
rect 24167 3009 24179 3043
rect 24688 3040 24716 3148
rect 24762 3136 24768 3188
rect 24820 3176 24826 3188
rect 25501 3179 25559 3185
rect 25501 3176 25513 3179
rect 24820 3148 25513 3176
rect 24820 3136 24826 3148
rect 25501 3145 25513 3148
rect 25547 3176 25559 3179
rect 26171 3179 26229 3185
rect 25547 3148 26004 3176
rect 25547 3145 25559 3148
rect 25501 3139 25559 3145
rect 25976 3117 26004 3148
rect 26171 3145 26183 3179
rect 26217 3176 26229 3179
rect 26878 3176 26884 3188
rect 26217 3148 26884 3176
rect 26217 3145 26229 3148
rect 26171 3139 26229 3145
rect 26878 3136 26884 3148
rect 26936 3176 26942 3188
rect 27173 3179 27231 3185
rect 27173 3176 27185 3179
rect 26936 3148 27185 3176
rect 26936 3136 26942 3148
rect 27173 3145 27185 3148
rect 27219 3145 27231 3179
rect 27173 3139 27231 3145
rect 25961 3111 26019 3117
rect 25961 3077 25973 3111
rect 26007 3077 26019 3111
rect 25961 3071 26019 3077
rect 26973 3111 27031 3117
rect 26973 3077 26985 3111
rect 27019 3108 27031 3111
rect 27338 3108 27344 3120
rect 27019 3080 27344 3108
rect 27019 3077 27031 3080
rect 26973 3071 27031 3077
rect 27338 3068 27344 3080
rect 27396 3068 27402 3120
rect 24688 3012 27384 3040
rect 24121 3003 24179 3009
rect 26329 2907 26387 2913
rect 21560 2876 22094 2904
rect 20809 2839 20867 2845
rect 20809 2805 20821 2839
rect 20855 2805 20867 2839
rect 20809 2799 20867 2805
rect 20993 2839 21051 2845
rect 20993 2805 21005 2839
rect 21039 2836 21051 2839
rect 21358 2836 21364 2848
rect 21039 2808 21364 2836
rect 21039 2805 21051 2808
rect 20993 2799 21051 2805
rect 21358 2796 21364 2808
rect 21416 2796 21422 2848
rect 22066 2836 22094 2876
rect 26329 2873 26341 2907
rect 26375 2904 26387 2907
rect 27246 2904 27252 2916
rect 26375 2876 27252 2904
rect 26375 2873 26387 2876
rect 26329 2867 26387 2873
rect 27246 2864 27252 2876
rect 27304 2864 27310 2916
rect 27356 2913 27384 3012
rect 27341 2907 27399 2913
rect 27341 2873 27353 2907
rect 27387 2873 27399 2907
rect 27341 2867 27399 2873
rect 22278 2836 22284 2848
rect 22066 2808 22284 2836
rect 22278 2796 22284 2808
rect 22336 2796 22342 2848
rect 23290 2796 23296 2848
rect 23348 2836 23354 2848
rect 23477 2839 23535 2845
rect 23477 2836 23489 2839
rect 23348 2808 23489 2836
rect 23348 2796 23354 2808
rect 23477 2805 23489 2808
rect 23523 2805 23535 2839
rect 23477 2799 23535 2805
rect 24026 2796 24032 2848
rect 24084 2836 24090 2848
rect 25958 2836 25964 2848
rect 24084 2808 25964 2836
rect 24084 2796 24090 2808
rect 25958 2796 25964 2808
rect 26016 2796 26022 2848
rect 26142 2836 26148 2848
rect 26103 2808 26148 2836
rect 26142 2796 26148 2808
rect 26200 2836 26206 2848
rect 27157 2839 27215 2845
rect 27157 2836 27169 2839
rect 26200 2808 27169 2836
rect 26200 2796 26206 2808
rect 27157 2805 27169 2808
rect 27203 2805 27215 2839
rect 27157 2799 27215 2805
rect 1104 2746 28060 2768
rect 1104 2694 5442 2746
rect 5494 2694 5506 2746
rect 5558 2694 5570 2746
rect 5622 2694 5634 2746
rect 5686 2694 5698 2746
rect 5750 2694 14428 2746
rect 14480 2694 14492 2746
rect 14544 2694 14556 2746
rect 14608 2694 14620 2746
rect 14672 2694 14684 2746
rect 14736 2694 23413 2746
rect 23465 2694 23477 2746
rect 23529 2694 23541 2746
rect 23593 2694 23605 2746
rect 23657 2694 23669 2746
rect 23721 2694 28060 2746
rect 1104 2672 28060 2694
rect 3602 2592 3608 2644
rect 3660 2632 3666 2644
rect 3789 2635 3847 2641
rect 3789 2632 3801 2635
rect 3660 2604 3801 2632
rect 3660 2592 3666 2604
rect 3789 2601 3801 2604
rect 3835 2601 3847 2635
rect 3789 2595 3847 2601
rect 5261 2635 5319 2641
rect 5261 2601 5273 2635
rect 5307 2632 5319 2635
rect 5810 2632 5816 2644
rect 5307 2604 5816 2632
rect 5307 2601 5319 2604
rect 5261 2595 5319 2601
rect 5810 2592 5816 2604
rect 5868 2592 5874 2644
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 8113 2635 8171 2641
rect 8113 2632 8125 2635
rect 7248 2604 8125 2632
rect 7248 2592 7254 2604
rect 8113 2601 8125 2604
rect 8159 2601 8171 2635
rect 8113 2595 8171 2601
rect 8294 2592 8300 2644
rect 8352 2632 8358 2644
rect 8941 2635 8999 2641
rect 8941 2632 8953 2635
rect 8352 2604 8953 2632
rect 8352 2592 8358 2604
rect 8941 2601 8953 2604
rect 8987 2601 8999 2635
rect 8941 2595 8999 2601
rect 10962 2592 10968 2644
rect 11020 2632 11026 2644
rect 11020 2604 11192 2632
rect 11020 2592 11026 2604
rect 11164 2576 11192 2604
rect 11790 2592 11796 2644
rect 11848 2632 11854 2644
rect 12158 2632 12164 2644
rect 11848 2604 12164 2632
rect 11848 2592 11854 2604
rect 12158 2592 12164 2604
rect 12216 2592 12222 2644
rect 13262 2592 13268 2644
rect 13320 2632 13326 2644
rect 13722 2632 13728 2644
rect 13320 2604 13728 2632
rect 13320 2592 13326 2604
rect 13722 2592 13728 2604
rect 13780 2592 13786 2644
rect 14737 2635 14795 2641
rect 14737 2601 14749 2635
rect 14783 2632 14795 2635
rect 14918 2632 14924 2644
rect 14783 2604 14924 2632
rect 14783 2601 14795 2604
rect 14737 2595 14795 2601
rect 14918 2592 14924 2604
rect 14976 2592 14982 2644
rect 15378 2632 15384 2644
rect 15339 2604 15384 2632
rect 15378 2592 15384 2604
rect 15436 2592 15442 2644
rect 15930 2632 15936 2644
rect 15891 2604 15936 2632
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 20070 2632 20076 2644
rect 16684 2604 20076 2632
rect 3510 2524 3516 2576
rect 3568 2564 3574 2576
rect 4890 2564 4896 2576
rect 3568 2536 4896 2564
rect 3568 2524 3574 2536
rect 4890 2524 4896 2536
rect 4948 2524 4954 2576
rect 6362 2564 6368 2576
rect 5092 2536 6368 2564
rect 3694 2456 3700 2508
rect 3752 2496 3758 2508
rect 3752 2468 5028 2496
rect 3752 2456 3758 2468
rect 2222 2388 2228 2440
rect 2280 2428 2286 2440
rect 2685 2431 2743 2437
rect 2685 2428 2697 2431
rect 2280 2400 2697 2428
rect 2280 2388 2286 2400
rect 2685 2397 2697 2400
rect 2731 2397 2743 2431
rect 2685 2391 2743 2397
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2397 4031 2431
rect 4706 2428 4712 2440
rect 4667 2400 4712 2428
rect 3973 2391 4031 2397
rect 290 2320 296 2372
rect 348 2360 354 2372
rect 1857 2363 1915 2369
rect 1857 2360 1869 2363
rect 348 2332 1869 2360
rect 348 2320 354 2332
rect 1857 2329 1869 2332
rect 1903 2329 1915 2363
rect 1857 2323 1915 2329
rect 2130 2292 2136 2304
rect 2091 2264 2136 2292
rect 2130 2252 2136 2264
rect 2188 2252 2194 2304
rect 2222 2252 2228 2304
rect 2280 2292 2286 2304
rect 2869 2295 2927 2301
rect 2869 2292 2881 2295
rect 2280 2264 2881 2292
rect 2280 2252 2286 2264
rect 2869 2261 2881 2264
rect 2915 2261 2927 2295
rect 3988 2292 4016 2391
rect 4706 2388 4712 2400
rect 4764 2388 4770 2440
rect 5000 2437 5028 2468
rect 5092 2437 5120 2536
rect 6362 2524 6368 2536
rect 6420 2564 6426 2576
rect 7285 2567 7343 2573
rect 6420 2536 7144 2564
rect 6420 2524 6426 2536
rect 7006 2456 7012 2508
rect 7064 2456 7070 2508
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2397 5043 2431
rect 4985 2391 5043 2397
rect 5077 2431 5135 2437
rect 5077 2397 5089 2431
rect 5123 2397 5135 2431
rect 5077 2391 5135 2397
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 7024 2428 7052 2456
rect 7116 2437 7144 2536
rect 7285 2533 7297 2567
rect 7331 2533 7343 2567
rect 7285 2527 7343 2533
rect 7300 2496 7328 2527
rect 10502 2524 10508 2576
rect 10560 2524 10566 2576
rect 10689 2567 10747 2573
rect 10689 2533 10701 2567
rect 10735 2533 10747 2567
rect 10689 2527 10747 2533
rect 10520 2496 10548 2524
rect 7300 2468 7972 2496
rect 6779 2400 7052 2428
rect 7101 2431 7159 2437
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 7101 2397 7113 2431
rect 7147 2397 7159 2431
rect 7834 2428 7840 2440
rect 7795 2400 7840 2428
rect 7101 2391 7159 2397
rect 7834 2388 7840 2400
rect 7892 2388 7898 2440
rect 7944 2437 7972 2468
rect 10336 2468 10548 2496
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2428 9183 2431
rect 9171 2400 9674 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 4893 2363 4951 2369
rect 4893 2329 4905 2363
rect 4939 2360 4951 2363
rect 5258 2360 5264 2372
rect 4939 2332 5264 2360
rect 4939 2329 4951 2332
rect 4893 2323 4951 2329
rect 5258 2320 5264 2332
rect 5316 2320 5322 2372
rect 6914 2360 6920 2372
rect 6875 2332 6920 2360
rect 6914 2320 6920 2332
rect 6972 2320 6978 2372
rect 7006 2320 7012 2372
rect 7064 2360 7070 2372
rect 7064 2332 7109 2360
rect 7064 2320 7070 2332
rect 5902 2292 5908 2304
rect 3988 2264 5908 2292
rect 2869 2255 2927 2261
rect 5902 2252 5908 2264
rect 5960 2252 5966 2304
rect 9646 2292 9674 2400
rect 9858 2388 9864 2440
rect 9916 2428 9922 2440
rect 10336 2437 10364 2468
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 9916 2400 10149 2428
rect 9916 2388 9922 2400
rect 10137 2397 10149 2400
rect 10183 2397 10195 2431
rect 10137 2391 10195 2397
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2428 10563 2431
rect 10594 2428 10600 2440
rect 10551 2400 10600 2428
rect 10551 2397 10563 2400
rect 10505 2391 10563 2397
rect 10594 2388 10600 2400
rect 10652 2388 10658 2440
rect 10704 2428 10732 2527
rect 11146 2524 11152 2576
rect 11204 2524 11210 2576
rect 11330 2524 11336 2576
rect 11388 2564 11394 2576
rect 13173 2567 13231 2573
rect 13173 2564 13185 2567
rect 11388 2536 13185 2564
rect 11388 2524 11394 2536
rect 13173 2533 13185 2536
rect 13219 2533 13231 2567
rect 13173 2527 13231 2533
rect 11517 2499 11575 2505
rect 11517 2465 11529 2499
rect 11563 2496 11575 2499
rect 12805 2499 12863 2505
rect 11563 2468 12434 2496
rect 11563 2465 11575 2468
rect 11517 2459 11575 2465
rect 12406 2440 12434 2468
rect 12805 2465 12817 2499
rect 12851 2496 12863 2499
rect 13354 2496 13360 2508
rect 12851 2468 13360 2496
rect 12851 2465 12863 2468
rect 12805 2459 12863 2465
rect 13354 2456 13360 2468
rect 13412 2456 13418 2508
rect 13906 2456 13912 2508
rect 13964 2496 13970 2508
rect 13964 2468 14596 2496
rect 13964 2456 13970 2468
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 10704 2400 11713 2428
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 11882 2388 11888 2440
rect 11940 2388 11946 2440
rect 12406 2400 12440 2440
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 12989 2431 13047 2437
rect 12989 2397 13001 2431
rect 13035 2428 13047 2431
rect 13262 2428 13268 2440
rect 13035 2400 13268 2428
rect 13035 2397 13047 2400
rect 12989 2391 13047 2397
rect 13262 2388 13268 2400
rect 13320 2388 13326 2440
rect 13372 2428 13400 2456
rect 14568 2437 14596 2468
rect 14369 2431 14427 2437
rect 14369 2428 14381 2431
rect 13372 2400 14381 2428
rect 14369 2397 14381 2400
rect 14415 2397 14427 2431
rect 14369 2391 14427 2397
rect 14553 2431 14611 2437
rect 14553 2397 14565 2431
rect 14599 2397 14611 2431
rect 14553 2391 14611 2397
rect 15197 2431 15255 2437
rect 15197 2397 15209 2431
rect 15243 2397 15255 2431
rect 16114 2428 16120 2440
rect 16075 2400 16120 2428
rect 15197 2391 15255 2397
rect 10413 2363 10471 2369
rect 10413 2329 10425 2363
rect 10459 2360 10471 2363
rect 10962 2360 10968 2372
rect 10459 2332 10968 2360
rect 10459 2329 10471 2332
rect 10413 2323 10471 2329
rect 10962 2320 10968 2332
rect 11020 2320 11026 2372
rect 11900 2360 11928 2388
rect 15212 2360 15240 2391
rect 16114 2388 16120 2400
rect 16172 2388 16178 2440
rect 16684 2437 16712 2604
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 20898 2592 20904 2644
rect 20956 2632 20962 2644
rect 21085 2635 21143 2641
rect 21085 2632 21097 2635
rect 20956 2604 21097 2632
rect 20956 2592 20962 2604
rect 21085 2601 21097 2604
rect 21131 2632 21143 2635
rect 21726 2632 21732 2644
rect 21131 2604 21732 2632
rect 21131 2601 21143 2604
rect 21085 2595 21143 2601
rect 21726 2592 21732 2604
rect 21784 2632 21790 2644
rect 22005 2635 22063 2641
rect 22005 2632 22017 2635
rect 21784 2604 22017 2632
rect 21784 2592 21790 2604
rect 22005 2601 22017 2604
rect 22051 2601 22063 2635
rect 22186 2632 22192 2644
rect 22147 2604 22192 2632
rect 22005 2595 22063 2601
rect 22186 2592 22192 2604
rect 22244 2592 22250 2644
rect 23569 2635 23627 2641
rect 23569 2632 23581 2635
rect 22756 2604 23581 2632
rect 19242 2524 19248 2576
rect 19300 2564 19306 2576
rect 20165 2567 20223 2573
rect 20165 2564 20177 2567
rect 19300 2536 20177 2564
rect 19300 2524 19306 2536
rect 20165 2533 20177 2536
rect 20211 2533 20223 2567
rect 20165 2527 20223 2533
rect 20622 2524 20628 2576
rect 20680 2564 20686 2576
rect 22756 2564 22784 2604
rect 23569 2601 23581 2604
rect 23615 2601 23627 2635
rect 23569 2595 23627 2601
rect 20680 2536 22784 2564
rect 22833 2567 22891 2573
rect 20680 2524 20686 2536
rect 22833 2533 22845 2567
rect 22879 2533 22891 2567
rect 22833 2527 22891 2533
rect 19886 2496 19892 2508
rect 18156 2468 19892 2496
rect 18156 2437 18184 2468
rect 19886 2456 19892 2468
rect 19944 2456 19950 2508
rect 20070 2456 20076 2508
rect 20128 2496 20134 2508
rect 22848 2496 22876 2527
rect 23014 2524 23020 2576
rect 23072 2564 23078 2576
rect 25317 2567 25375 2573
rect 25317 2564 25329 2567
rect 23072 2536 25329 2564
rect 23072 2524 23078 2536
rect 25317 2533 25329 2536
rect 25363 2533 25375 2567
rect 25317 2527 25375 2533
rect 23290 2496 23296 2508
rect 20128 2468 22876 2496
rect 22940 2468 23296 2496
rect 20128 2456 20134 2468
rect 16669 2431 16727 2437
rect 16669 2397 16681 2431
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 17405 2431 17463 2437
rect 17405 2397 17417 2431
rect 17451 2397 17463 2431
rect 17405 2391 17463 2397
rect 18141 2431 18199 2437
rect 18141 2397 18153 2431
rect 18187 2397 18199 2431
rect 18141 2391 18199 2397
rect 19245 2431 19303 2437
rect 19245 2397 19257 2431
rect 19291 2428 19303 2431
rect 19610 2428 19616 2440
rect 19291 2400 19616 2428
rect 19291 2397 19303 2400
rect 19245 2391 19303 2397
rect 11900 2332 15240 2360
rect 17420 2360 17448 2391
rect 19610 2388 19616 2400
rect 19668 2388 19674 2440
rect 19981 2431 20039 2437
rect 19981 2397 19993 2431
rect 20027 2428 20039 2431
rect 20806 2428 20812 2440
rect 20027 2400 20812 2428
rect 20027 2397 20039 2400
rect 19981 2391 20039 2397
rect 20806 2388 20812 2400
rect 20864 2388 20870 2440
rect 22646 2428 22652 2440
rect 22607 2400 22652 2428
rect 22646 2388 22652 2400
rect 22704 2388 22710 2440
rect 18230 2360 18236 2372
rect 17420 2332 18236 2360
rect 18230 2320 18236 2332
rect 18288 2320 18294 2372
rect 20714 2320 20720 2372
rect 20772 2360 20778 2372
rect 20901 2363 20959 2369
rect 20901 2360 20913 2363
rect 20772 2332 20913 2360
rect 20772 2320 20778 2332
rect 20901 2329 20913 2332
rect 20947 2329 20959 2363
rect 20901 2323 20959 2329
rect 20990 2320 20996 2372
rect 21048 2360 21054 2372
rect 21101 2363 21159 2369
rect 21101 2360 21113 2363
rect 21048 2332 21113 2360
rect 21048 2320 21054 2332
rect 21101 2329 21113 2332
rect 21147 2360 21159 2363
rect 21821 2363 21879 2369
rect 21147 2332 21395 2360
rect 21147 2329 21159 2332
rect 21101 2323 21159 2329
rect 11054 2292 11060 2304
rect 9646 2264 11060 2292
rect 11054 2252 11060 2264
rect 11112 2252 11118 2304
rect 11882 2292 11888 2304
rect 11843 2264 11888 2292
rect 11882 2252 11888 2264
rect 11940 2252 11946 2304
rect 12158 2252 12164 2304
rect 12216 2292 12222 2304
rect 16758 2292 16764 2304
rect 12216 2264 16764 2292
rect 12216 2252 12222 2264
rect 16758 2252 16764 2264
rect 16816 2252 16822 2304
rect 16850 2252 16856 2304
rect 16908 2292 16914 2304
rect 16908 2264 16953 2292
rect 16908 2252 16914 2264
rect 17310 2252 17316 2304
rect 17368 2292 17374 2304
rect 17589 2295 17647 2301
rect 17589 2292 17601 2295
rect 17368 2264 17601 2292
rect 17368 2252 17374 2264
rect 17589 2261 17601 2264
rect 17635 2261 17647 2295
rect 17589 2255 17647 2261
rect 17862 2252 17868 2304
rect 17920 2292 17926 2304
rect 18325 2295 18383 2301
rect 18325 2292 18337 2295
rect 17920 2264 18337 2292
rect 17920 2252 17926 2264
rect 18325 2261 18337 2264
rect 18371 2261 18383 2295
rect 18325 2255 18383 2261
rect 18414 2252 18420 2304
rect 18472 2292 18478 2304
rect 19429 2295 19487 2301
rect 19429 2292 19441 2295
rect 18472 2264 19441 2292
rect 18472 2252 18478 2264
rect 19429 2261 19441 2264
rect 19475 2261 19487 2295
rect 21266 2292 21272 2304
rect 21227 2264 21272 2292
rect 19429 2255 19487 2261
rect 21266 2252 21272 2264
rect 21324 2252 21330 2304
rect 21367 2292 21395 2332
rect 21821 2329 21833 2363
rect 21867 2360 21879 2363
rect 22940 2360 22968 2468
rect 23290 2456 23296 2468
rect 23348 2456 23354 2508
rect 23934 2456 23940 2508
rect 23992 2496 23998 2508
rect 23992 2468 25912 2496
rect 23992 2456 23998 2468
rect 23198 2388 23204 2440
rect 23256 2428 23262 2440
rect 23385 2431 23443 2437
rect 23385 2428 23397 2431
rect 23256 2400 23397 2428
rect 23256 2388 23262 2400
rect 23385 2397 23397 2400
rect 23431 2397 23443 2431
rect 23385 2391 23443 2397
rect 24302 2388 24308 2440
rect 24360 2428 24366 2440
rect 24397 2431 24455 2437
rect 24397 2428 24409 2431
rect 24360 2400 24409 2428
rect 24360 2388 24366 2400
rect 24397 2397 24409 2400
rect 24443 2397 24455 2431
rect 25130 2428 25136 2440
rect 25091 2400 25136 2428
rect 24397 2391 24455 2397
rect 25130 2388 25136 2400
rect 25188 2388 25194 2440
rect 25884 2437 25912 2468
rect 25869 2431 25927 2437
rect 25869 2397 25881 2431
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 27157 2363 27215 2369
rect 21867 2332 22968 2360
rect 23308 2332 26096 2360
rect 21867 2329 21879 2332
rect 21821 2323 21879 2329
rect 22021 2295 22079 2301
rect 22021 2292 22033 2295
rect 21367 2264 22033 2292
rect 22021 2261 22033 2264
rect 22067 2261 22079 2295
rect 22021 2255 22079 2261
rect 22186 2252 22192 2304
rect 22244 2292 22250 2304
rect 23308 2292 23336 2332
rect 22244 2264 23336 2292
rect 22244 2252 22250 2264
rect 23382 2252 23388 2304
rect 23440 2292 23446 2304
rect 26068 2301 26096 2332
rect 27157 2329 27169 2363
rect 27203 2360 27215 2363
rect 28994 2360 29000 2372
rect 27203 2332 29000 2360
rect 27203 2329 27215 2332
rect 27157 2323 27215 2329
rect 28994 2320 29000 2332
rect 29052 2320 29058 2372
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 23440 2264 24593 2292
rect 23440 2252 23446 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 26053 2295 26111 2301
rect 26053 2261 26065 2295
rect 26099 2261 26111 2295
rect 27246 2292 27252 2304
rect 27207 2264 27252 2292
rect 26053 2255 26111 2261
rect 27246 2252 27252 2264
rect 27304 2252 27310 2304
rect 1104 2202 28060 2224
rect 1104 2150 9935 2202
rect 9987 2150 9999 2202
rect 10051 2150 10063 2202
rect 10115 2150 10127 2202
rect 10179 2150 10191 2202
rect 10243 2150 18920 2202
rect 18972 2150 18984 2202
rect 19036 2150 19048 2202
rect 19100 2150 19112 2202
rect 19164 2150 19176 2202
rect 19228 2150 28060 2202
rect 1104 2128 28060 2150
rect 3142 2048 3148 2100
rect 3200 2088 3206 2100
rect 7006 2088 7012 2100
rect 3200 2060 7012 2088
rect 3200 2048 3206 2060
rect 7006 2048 7012 2060
rect 7064 2048 7070 2100
rect 16758 2048 16764 2100
rect 16816 2088 16822 2100
rect 27246 2088 27252 2100
rect 16816 2060 27252 2088
rect 16816 2048 16822 2060
rect 27246 2048 27252 2060
rect 27304 2048 27310 2100
rect 2130 1980 2136 2032
rect 2188 2020 2194 2032
rect 9030 2020 9036 2032
rect 2188 1992 9036 2020
rect 2188 1980 2194 1992
rect 9030 1980 9036 1992
rect 9088 1980 9094 2032
rect 16850 1980 16856 2032
rect 16908 2020 16914 2032
rect 27062 2020 27068 2032
rect 16908 1992 27068 2020
rect 16908 1980 16914 1992
rect 27062 1980 27068 1992
rect 27120 1980 27126 2032
rect 3786 1912 3792 1964
rect 3844 1952 3850 1964
rect 11882 1952 11888 1964
rect 3844 1924 11888 1952
rect 3844 1912 3850 1924
rect 11882 1912 11888 1924
rect 11940 1912 11946 1964
rect 16758 1912 16764 1964
rect 16816 1952 16822 1964
rect 17126 1952 17132 1964
rect 16816 1924 17132 1952
rect 16816 1912 16822 1924
rect 17126 1912 17132 1924
rect 17184 1912 17190 1964
rect 19518 1912 19524 1964
rect 19576 1952 19582 1964
rect 20346 1952 20352 1964
rect 19576 1924 20352 1952
rect 19576 1912 19582 1924
rect 20346 1912 20352 1924
rect 20404 1912 20410 1964
rect 21266 1912 21272 1964
rect 21324 1952 21330 1964
rect 24118 1952 24124 1964
rect 21324 1924 24124 1952
rect 21324 1912 21330 1924
rect 24118 1912 24124 1924
rect 24176 1912 24182 1964
rect 21082 1436 21088 1488
rect 21140 1476 21146 1488
rect 23382 1476 23388 1488
rect 21140 1448 23388 1476
rect 21140 1436 21146 1448
rect 23382 1436 23388 1448
rect 23440 1436 23446 1488
rect 21634 1368 21640 1420
rect 21692 1408 21698 1420
rect 23014 1408 23020 1420
rect 21692 1380 23020 1408
rect 21692 1368 21698 1380
rect 23014 1368 23020 1380
rect 23072 1368 23078 1420
rect 18782 1028 18788 1080
rect 18840 1068 18846 1080
rect 19242 1068 19248 1080
rect 18840 1040 19248 1068
rect 18840 1028 18846 1040
rect 19242 1028 19248 1040
rect 19300 1028 19306 1080
<< via1 >>
rect 5442 28806 5494 28858
rect 5506 28806 5558 28858
rect 5570 28806 5622 28858
rect 5634 28806 5686 28858
rect 5698 28806 5750 28858
rect 14428 28806 14480 28858
rect 14492 28806 14544 28858
rect 14556 28806 14608 28858
rect 14620 28806 14672 28858
rect 14684 28806 14736 28858
rect 23413 28806 23465 28858
rect 23477 28806 23529 28858
rect 23541 28806 23593 28858
rect 23605 28806 23657 28858
rect 23669 28806 23721 28858
rect 12808 28704 12860 28756
rect 9128 28636 9180 28688
rect 15752 28704 15804 28756
rect 16672 28704 16724 28756
rect 13544 28636 13596 28688
rect 18328 28636 18380 28688
rect 20168 28636 20220 28688
rect 8300 28500 8352 28552
rect 8392 28543 8444 28552
rect 8392 28509 8401 28543
rect 8401 28509 8435 28543
rect 8435 28509 8444 28543
rect 8392 28500 8444 28509
rect 10508 28500 10560 28552
rect 11336 28543 11388 28552
rect 11336 28509 11345 28543
rect 11345 28509 11379 28543
rect 11379 28509 11388 28543
rect 11336 28500 11388 28509
rect 14004 28568 14056 28620
rect 19248 28568 19300 28620
rect 22100 28636 22152 28688
rect 8576 28475 8628 28484
rect 8576 28441 8585 28475
rect 8585 28441 8619 28475
rect 8619 28441 8628 28475
rect 8576 28432 8628 28441
rect 8760 28475 8812 28484
rect 8760 28441 8769 28475
rect 8769 28441 8803 28475
rect 8803 28441 8812 28475
rect 8760 28432 8812 28441
rect 13176 28543 13228 28552
rect 13176 28509 13185 28543
rect 13185 28509 13219 28543
rect 13219 28509 13228 28543
rect 13176 28500 13228 28509
rect 13728 28500 13780 28552
rect 15016 28543 15068 28552
rect 15016 28509 15025 28543
rect 15025 28509 15059 28543
rect 15059 28509 15068 28543
rect 15016 28500 15068 28509
rect 16488 28543 16540 28552
rect 16488 28509 16497 28543
rect 16497 28509 16531 28543
rect 16531 28509 16540 28543
rect 16488 28500 16540 28509
rect 17592 28500 17644 28552
rect 18144 28543 18196 28552
rect 18144 28509 18153 28543
rect 18153 28509 18187 28543
rect 18187 28509 18196 28543
rect 18144 28500 18196 28509
rect 18696 28543 18748 28552
rect 18696 28509 18705 28543
rect 18705 28509 18739 28543
rect 18739 28509 18748 28543
rect 18696 28500 18748 28509
rect 19800 28500 19852 28552
rect 20628 28500 20680 28552
rect 21640 28543 21692 28552
rect 21640 28509 21649 28543
rect 21649 28509 21683 28543
rect 21683 28509 21692 28543
rect 21640 28500 21692 28509
rect 22928 28500 22980 28552
rect 27344 28543 27396 28552
rect 27344 28509 27353 28543
rect 27353 28509 27387 28543
rect 27387 28509 27396 28543
rect 27344 28500 27396 28509
rect 4344 28364 4396 28416
rect 7104 28364 7156 28416
rect 7472 28364 7524 28416
rect 10416 28364 10468 28416
rect 10968 28364 11020 28416
rect 11152 28407 11204 28416
rect 11152 28373 11161 28407
rect 11161 28373 11195 28407
rect 11195 28373 11204 28407
rect 11152 28364 11204 28373
rect 11980 28364 12032 28416
rect 12164 28407 12216 28416
rect 12164 28373 12173 28407
rect 12173 28373 12207 28407
rect 12207 28373 12216 28407
rect 12164 28364 12216 28373
rect 13084 28407 13136 28416
rect 13084 28373 13093 28407
rect 13093 28373 13127 28407
rect 13127 28373 13136 28407
rect 13084 28364 13136 28373
rect 13820 28364 13872 28416
rect 14832 28407 14884 28416
rect 14832 28373 14841 28407
rect 14841 28373 14875 28407
rect 14875 28373 14884 28407
rect 14832 28364 14884 28373
rect 15568 28407 15620 28416
rect 15568 28373 15577 28407
rect 15577 28373 15611 28407
rect 15611 28373 15620 28407
rect 15568 28364 15620 28373
rect 21824 28432 21876 28484
rect 16856 28364 16908 28416
rect 17316 28407 17368 28416
rect 17316 28373 17325 28407
rect 17325 28373 17359 28407
rect 17359 28373 17368 28407
rect 17316 28364 17368 28373
rect 18604 28364 18656 28416
rect 19616 28364 19668 28416
rect 20720 28407 20772 28416
rect 20720 28373 20729 28407
rect 20729 28373 20763 28407
rect 20763 28373 20772 28407
rect 20720 28364 20772 28373
rect 22192 28364 22244 28416
rect 27068 28364 27120 28416
rect 9935 28262 9987 28314
rect 9999 28262 10051 28314
rect 10063 28262 10115 28314
rect 10127 28262 10179 28314
rect 10191 28262 10243 28314
rect 18920 28262 18972 28314
rect 18984 28262 19036 28314
rect 19048 28262 19100 28314
rect 19112 28262 19164 28314
rect 19176 28262 19228 28314
rect 4344 28203 4396 28212
rect 4344 28169 4353 28203
rect 4353 28169 4387 28203
rect 4387 28169 4396 28203
rect 4344 28160 4396 28169
rect 5908 28160 5960 28212
rect 4252 28092 4304 28144
rect 12808 28160 12860 28212
rect 16120 28160 16172 28212
rect 3884 27820 3936 27872
rect 5264 28024 5316 28076
rect 9680 28092 9732 28144
rect 9864 28067 9916 28076
rect 9864 28033 9898 28067
rect 9898 28033 9916 28067
rect 9864 28024 9916 28033
rect 6552 27956 6604 28008
rect 10968 27956 11020 28008
rect 12532 28024 12584 28076
rect 13912 27956 13964 28008
rect 16764 28024 16816 28076
rect 16948 28067 17000 28076
rect 16948 28033 16982 28067
rect 16982 28033 17000 28067
rect 16948 28024 17000 28033
rect 19708 28092 19760 28144
rect 18604 28024 18656 28076
rect 19616 28024 19668 28076
rect 22284 28024 22336 28076
rect 23296 28024 23348 28076
rect 26884 28024 26936 28076
rect 27160 28067 27212 28076
rect 27160 28033 27169 28067
rect 27169 28033 27203 28067
rect 27203 28033 27212 28067
rect 27160 28024 27212 28033
rect 27804 27956 27856 28008
rect 6828 27888 6880 27940
rect 25872 27888 25924 27940
rect 5816 27863 5868 27872
rect 5816 27829 5825 27863
rect 5825 27829 5859 27863
rect 5859 27829 5868 27863
rect 5816 27820 5868 27829
rect 8576 27863 8628 27872
rect 8576 27829 8585 27863
rect 8585 27829 8619 27863
rect 8619 27829 8628 27863
rect 8576 27820 8628 27829
rect 9220 27820 9272 27872
rect 10692 27820 10744 27872
rect 13176 27820 13228 27872
rect 13544 27820 13596 27872
rect 15292 27820 15344 27872
rect 18052 27863 18104 27872
rect 18052 27829 18061 27863
rect 18061 27829 18095 27863
rect 18095 27829 18104 27863
rect 18052 27820 18104 27829
rect 19432 27820 19484 27872
rect 20352 27863 20404 27872
rect 20352 27829 20361 27863
rect 20361 27829 20395 27863
rect 20395 27829 20404 27863
rect 20352 27820 20404 27829
rect 20996 27863 21048 27872
rect 20996 27829 21005 27863
rect 21005 27829 21039 27863
rect 21039 27829 21048 27863
rect 20996 27820 21048 27829
rect 22376 27863 22428 27872
rect 22376 27829 22385 27863
rect 22385 27829 22419 27863
rect 22419 27829 22428 27863
rect 22376 27820 22428 27829
rect 22744 27820 22796 27872
rect 23296 27863 23348 27872
rect 23296 27829 23305 27863
rect 23305 27829 23339 27863
rect 23339 27829 23348 27863
rect 23296 27820 23348 27829
rect 23848 27820 23900 27872
rect 26608 27820 26660 27872
rect 5442 27718 5494 27770
rect 5506 27718 5558 27770
rect 5570 27718 5622 27770
rect 5634 27718 5686 27770
rect 5698 27718 5750 27770
rect 14428 27718 14480 27770
rect 14492 27718 14544 27770
rect 14556 27718 14608 27770
rect 14620 27718 14672 27770
rect 14684 27718 14736 27770
rect 23413 27718 23465 27770
rect 23477 27718 23529 27770
rect 23541 27718 23593 27770
rect 23605 27718 23657 27770
rect 23669 27718 23721 27770
rect 4344 27548 4396 27600
rect 5448 27548 5500 27600
rect 5540 27548 5592 27600
rect 5816 27548 5868 27600
rect 6644 27616 6696 27668
rect 4160 27480 4212 27532
rect 4988 27480 5040 27532
rect 2596 27455 2648 27464
rect 2596 27421 2605 27455
rect 2605 27421 2639 27455
rect 2639 27421 2648 27455
rect 2596 27412 2648 27421
rect 3700 27412 3752 27464
rect 4712 27455 4764 27464
rect 4712 27421 4721 27455
rect 4721 27421 4755 27455
rect 4755 27421 4764 27455
rect 4712 27412 4764 27421
rect 6000 27412 6052 27464
rect 6460 27455 6512 27464
rect 6460 27421 6469 27455
rect 6469 27421 6503 27455
rect 6503 27421 6512 27455
rect 6460 27412 6512 27421
rect 8116 27412 8168 27464
rect 9680 27616 9732 27668
rect 10968 27616 11020 27668
rect 13084 27616 13136 27668
rect 18144 27616 18196 27668
rect 21640 27616 21692 27668
rect 21824 27616 21876 27668
rect 27620 27616 27672 27668
rect 13912 27548 13964 27600
rect 18236 27548 18288 27600
rect 25228 27548 25280 27600
rect 27160 27548 27212 27600
rect 5172 27344 5224 27396
rect 6368 27344 6420 27396
rect 9128 27344 9180 27396
rect 10968 27412 11020 27464
rect 11152 27412 11204 27464
rect 13544 27455 13596 27464
rect 13544 27421 13553 27455
rect 13553 27421 13587 27455
rect 13587 27421 13596 27455
rect 13544 27412 13596 27421
rect 14004 27480 14056 27532
rect 18696 27480 18748 27532
rect 21824 27523 21876 27532
rect 13820 27412 13872 27464
rect 13912 27455 13964 27464
rect 13912 27421 13921 27455
rect 13921 27421 13955 27455
rect 13955 27421 13964 27455
rect 13912 27412 13964 27421
rect 2504 27276 2556 27328
rect 3056 27319 3108 27328
rect 3056 27285 3065 27319
rect 3065 27285 3099 27319
rect 3099 27285 3108 27319
rect 3056 27276 3108 27285
rect 3700 27276 3752 27328
rect 4344 27276 4396 27328
rect 6828 27276 6880 27328
rect 7840 27319 7892 27328
rect 7840 27285 7849 27319
rect 7849 27285 7883 27319
rect 7883 27285 7892 27319
rect 7840 27276 7892 27285
rect 8024 27276 8076 27328
rect 14096 27344 14148 27396
rect 16028 27412 16080 27464
rect 10324 27319 10376 27328
rect 10324 27285 10333 27319
rect 10333 27285 10367 27319
rect 10367 27285 10376 27319
rect 10324 27276 10376 27285
rect 12440 27319 12492 27328
rect 12440 27285 12449 27319
rect 12449 27285 12483 27319
rect 12483 27285 12492 27319
rect 12440 27276 12492 27285
rect 12716 27276 12768 27328
rect 14924 27319 14976 27328
rect 14924 27285 14933 27319
rect 14933 27285 14967 27319
rect 14967 27285 14976 27319
rect 14924 27276 14976 27285
rect 15200 27319 15252 27328
rect 15200 27285 15209 27319
rect 15209 27285 15243 27319
rect 15243 27285 15252 27319
rect 15200 27276 15252 27285
rect 15660 27319 15712 27328
rect 15660 27285 15669 27319
rect 15669 27285 15703 27319
rect 15703 27285 15712 27319
rect 15660 27276 15712 27285
rect 18512 27455 18564 27464
rect 17132 27344 17184 27396
rect 18512 27421 18521 27455
rect 18521 27421 18555 27455
rect 18555 27421 18564 27455
rect 18512 27412 18564 27421
rect 19892 27412 19944 27464
rect 21824 27489 21833 27523
rect 21833 27489 21867 27523
rect 21867 27489 21876 27523
rect 21824 27480 21876 27489
rect 23204 27480 23256 27532
rect 21180 27412 21232 27464
rect 22100 27455 22152 27464
rect 22100 27421 22134 27455
rect 22134 27421 22152 27455
rect 20352 27344 20404 27396
rect 22100 27412 22152 27421
rect 22468 27344 22520 27396
rect 16580 27276 16632 27328
rect 17040 27276 17092 27328
rect 20076 27276 20128 27328
rect 21548 27276 21600 27328
rect 23756 27412 23808 27464
rect 24584 27455 24636 27464
rect 24584 27421 24593 27455
rect 24593 27421 24627 27455
rect 24627 27421 24636 27455
rect 24584 27412 24636 27421
rect 24216 27344 24268 27396
rect 24308 27344 24360 27396
rect 26056 27412 26108 27464
rect 26976 27412 27028 27464
rect 27160 27412 27212 27464
rect 23020 27276 23072 27328
rect 23940 27276 23992 27328
rect 24492 27276 24544 27328
rect 25136 27276 25188 27328
rect 25780 27319 25832 27328
rect 25780 27285 25789 27319
rect 25789 27285 25823 27319
rect 25823 27285 25832 27319
rect 25780 27276 25832 27285
rect 26332 27276 26384 27328
rect 27252 27319 27304 27328
rect 27252 27285 27261 27319
rect 27261 27285 27295 27319
rect 27295 27285 27304 27319
rect 27252 27276 27304 27285
rect 9935 27174 9987 27226
rect 9999 27174 10051 27226
rect 10063 27174 10115 27226
rect 10127 27174 10179 27226
rect 10191 27174 10243 27226
rect 18920 27174 18972 27226
rect 18984 27174 19036 27226
rect 19048 27174 19100 27226
rect 19112 27174 19164 27226
rect 19176 27174 19228 27226
rect 2596 27072 2648 27124
rect 4068 27072 4120 27124
rect 4160 27072 4212 27124
rect 5264 27115 5316 27124
rect 1400 26936 1452 26988
rect 2872 26936 2924 26988
rect 4252 27004 4304 27056
rect 1860 26868 1912 26920
rect 4528 26936 4580 26988
rect 5264 27081 5273 27115
rect 5273 27081 5307 27115
rect 5307 27081 5316 27115
rect 5264 27072 5316 27081
rect 5816 27072 5868 27124
rect 6368 27115 6420 27124
rect 6368 27081 6377 27115
rect 6377 27081 6411 27115
rect 6411 27081 6420 27115
rect 6368 27072 6420 27081
rect 5540 26979 5592 26988
rect 5540 26945 5549 26979
rect 5549 26945 5583 26979
rect 5583 26945 5592 26979
rect 5540 26936 5592 26945
rect 6092 26936 6144 26988
rect 7012 27072 7064 27124
rect 11336 27072 11388 27124
rect 12532 27115 12584 27124
rect 12532 27081 12541 27115
rect 12541 27081 12575 27115
rect 12575 27081 12584 27115
rect 12532 27072 12584 27081
rect 15660 27072 15712 27124
rect 7288 27004 7340 27056
rect 7564 27004 7616 27056
rect 10876 27004 10928 27056
rect 6184 26868 6236 26920
rect 7196 26936 7248 26988
rect 8576 26936 8628 26988
rect 9220 26979 9272 26988
rect 9220 26945 9229 26979
rect 9229 26945 9263 26979
rect 9263 26945 9272 26979
rect 9220 26936 9272 26945
rect 9404 26936 9456 26988
rect 10692 26936 10744 26988
rect 11520 26979 11572 26988
rect 11520 26945 11529 26979
rect 11529 26945 11563 26979
rect 11563 26945 11572 26979
rect 11520 26936 11572 26945
rect 12716 26979 12768 26988
rect 7472 26868 7524 26920
rect 7840 26868 7892 26920
rect 1676 26732 1728 26784
rect 2872 26732 2924 26784
rect 7564 26800 7616 26852
rect 8116 26868 8168 26920
rect 10600 26868 10652 26920
rect 11428 26868 11480 26920
rect 12716 26945 12725 26979
rect 12725 26945 12759 26979
rect 12759 26945 12768 26979
rect 12716 26936 12768 26945
rect 12900 27004 12952 27056
rect 18512 27072 18564 27124
rect 27160 27115 27212 27124
rect 13176 26868 13228 26920
rect 13820 26936 13872 26988
rect 14004 26979 14056 26988
rect 14004 26945 14013 26979
rect 14013 26945 14047 26979
rect 14047 26945 14056 26979
rect 14004 26936 14056 26945
rect 14740 26979 14792 26988
rect 14740 26945 14774 26979
rect 14774 26945 14792 26979
rect 19340 27004 19392 27056
rect 14740 26936 14792 26945
rect 16764 26936 16816 26988
rect 17684 26936 17736 26988
rect 18696 26979 18748 26988
rect 18696 26945 18705 26979
rect 18705 26945 18739 26979
rect 18739 26945 18748 26979
rect 18696 26936 18748 26945
rect 4896 26732 4948 26784
rect 5080 26732 5132 26784
rect 5356 26732 5408 26784
rect 8668 26732 8720 26784
rect 9680 26732 9732 26784
rect 11152 26732 11204 26784
rect 13268 26800 13320 26852
rect 12072 26732 12124 26784
rect 14280 26732 14332 26784
rect 17960 26868 18012 26920
rect 19616 26868 19668 26920
rect 20352 27004 20404 27056
rect 27160 27081 27169 27115
rect 27169 27081 27203 27115
rect 27203 27081 27212 27115
rect 27160 27072 27212 27081
rect 19892 26979 19944 26988
rect 19892 26945 19901 26979
rect 19901 26945 19935 26979
rect 19935 26945 19944 26979
rect 19892 26936 19944 26945
rect 21272 26936 21324 26988
rect 22008 26979 22060 26988
rect 22008 26945 22017 26979
rect 22017 26945 22051 26979
rect 22051 26945 22060 26979
rect 22652 26979 22704 26988
rect 22008 26936 22060 26945
rect 22652 26945 22661 26979
rect 22661 26945 22695 26979
rect 22695 26945 22704 26979
rect 22652 26936 22704 26945
rect 22836 26936 22888 26988
rect 23848 26936 23900 26988
rect 24216 26936 24268 26988
rect 25964 26936 26016 26988
rect 26424 26979 26476 26988
rect 26424 26945 26433 26979
rect 26433 26945 26467 26979
rect 26467 26945 26476 26979
rect 26424 26936 26476 26945
rect 15384 26732 15436 26784
rect 15844 26775 15896 26784
rect 15844 26741 15853 26775
rect 15853 26741 15887 26775
rect 15887 26741 15896 26775
rect 15844 26732 15896 26741
rect 15936 26732 15988 26784
rect 21456 26800 21508 26852
rect 22284 26800 22336 26852
rect 18144 26732 18196 26784
rect 20812 26732 20864 26784
rect 21640 26732 21692 26784
rect 23112 26775 23164 26784
rect 23112 26741 23121 26775
rect 23121 26741 23155 26775
rect 23155 26741 23164 26775
rect 23112 26732 23164 26741
rect 24216 26732 24268 26784
rect 25688 26732 25740 26784
rect 26240 26775 26292 26784
rect 26240 26741 26249 26775
rect 26249 26741 26283 26775
rect 26283 26741 26292 26775
rect 26240 26732 26292 26741
rect 5442 26630 5494 26682
rect 5506 26630 5558 26682
rect 5570 26630 5622 26682
rect 5634 26630 5686 26682
rect 5698 26630 5750 26682
rect 14428 26630 14480 26682
rect 14492 26630 14544 26682
rect 14556 26630 14608 26682
rect 14620 26630 14672 26682
rect 14684 26630 14736 26682
rect 23413 26630 23465 26682
rect 23477 26630 23529 26682
rect 23541 26630 23593 26682
rect 23605 26630 23657 26682
rect 23669 26630 23721 26682
rect 4528 26571 4580 26580
rect 4528 26537 4537 26571
rect 4537 26537 4571 26571
rect 4571 26537 4580 26571
rect 4528 26528 4580 26537
rect 5816 26528 5868 26580
rect 7472 26528 7524 26580
rect 8208 26528 8260 26580
rect 8300 26528 8352 26580
rect 9864 26528 9916 26580
rect 10048 26528 10100 26580
rect 11428 26528 11480 26580
rect 14280 26528 14332 26580
rect 14832 26528 14884 26580
rect 16028 26528 16080 26580
rect 19800 26571 19852 26580
rect 19800 26537 19809 26571
rect 19809 26537 19843 26571
rect 19843 26537 19852 26571
rect 19800 26528 19852 26537
rect 21456 26571 21508 26580
rect 21456 26537 21465 26571
rect 21465 26537 21499 26571
rect 21499 26537 21508 26571
rect 21456 26528 21508 26537
rect 1584 26460 1636 26512
rect 3424 26460 3476 26512
rect 3516 26324 3568 26376
rect 4160 26367 4212 26376
rect 2688 26256 2740 26308
rect 4160 26333 4169 26367
rect 4169 26333 4203 26367
rect 4203 26333 4212 26367
rect 4160 26324 4212 26333
rect 4896 26392 4948 26444
rect 4804 26367 4856 26376
rect 4804 26333 4813 26367
rect 4813 26333 4847 26367
rect 4847 26333 4856 26367
rect 5172 26460 5224 26512
rect 4804 26324 4856 26333
rect 4068 26256 4120 26308
rect 5356 26392 5408 26444
rect 5448 26392 5500 26444
rect 5264 26367 5316 26376
rect 5264 26333 5273 26367
rect 5273 26333 5307 26367
rect 5307 26333 5316 26367
rect 5264 26324 5316 26333
rect 5632 26324 5684 26376
rect 6092 26324 6144 26376
rect 6184 26367 6236 26376
rect 6184 26333 6193 26367
rect 6193 26333 6227 26367
rect 6227 26333 6236 26367
rect 6184 26324 6236 26333
rect 7472 26324 7524 26376
rect 8392 26460 8444 26512
rect 8024 26392 8076 26444
rect 10324 26460 10376 26512
rect 14004 26460 14056 26512
rect 10048 26392 10100 26444
rect 12532 26392 12584 26444
rect 12900 26435 12952 26444
rect 12900 26401 12909 26435
rect 12909 26401 12943 26435
rect 12943 26401 12952 26435
rect 12900 26392 12952 26401
rect 2964 26188 3016 26240
rect 4896 26188 4948 26240
rect 5908 26188 5960 26240
rect 6460 26188 6512 26240
rect 8668 26256 8720 26308
rect 10416 26367 10468 26376
rect 10416 26333 10425 26367
rect 10425 26333 10459 26367
rect 10459 26333 10468 26367
rect 10416 26324 10468 26333
rect 7196 26188 7248 26240
rect 7472 26188 7524 26240
rect 9772 26188 9824 26240
rect 10416 26188 10468 26240
rect 10600 26367 10652 26376
rect 10600 26333 10609 26367
rect 10609 26333 10643 26367
rect 10643 26333 10652 26367
rect 10600 26324 10652 26333
rect 10876 26324 10928 26376
rect 11428 26314 11480 26366
rect 12256 26324 12308 26376
rect 14096 26367 14148 26376
rect 14096 26333 14105 26367
rect 14105 26333 14139 26367
rect 14139 26333 14148 26367
rect 14096 26324 14148 26333
rect 16488 26460 16540 26512
rect 14556 26367 14608 26376
rect 14556 26333 14565 26367
rect 14565 26333 14599 26367
rect 14599 26333 14608 26367
rect 14556 26324 14608 26333
rect 18788 26392 18840 26444
rect 22652 26528 22704 26580
rect 27712 26528 27764 26580
rect 26516 26460 26568 26512
rect 20536 26392 20588 26444
rect 21824 26392 21876 26444
rect 13360 26256 13412 26308
rect 17500 26324 17552 26376
rect 17684 26324 17736 26376
rect 17960 26367 18012 26376
rect 17960 26333 17969 26367
rect 17969 26333 18003 26367
rect 18003 26333 18012 26367
rect 17960 26324 18012 26333
rect 19432 26367 19484 26376
rect 17776 26299 17828 26308
rect 17776 26265 17785 26299
rect 17785 26265 17819 26299
rect 17819 26265 17828 26299
rect 17776 26256 17828 26265
rect 18052 26256 18104 26308
rect 18420 26256 18472 26308
rect 19432 26333 19441 26367
rect 19441 26333 19475 26367
rect 19475 26333 19484 26367
rect 19432 26324 19484 26333
rect 19616 26367 19668 26376
rect 19616 26333 19625 26367
rect 19625 26333 19659 26367
rect 19659 26333 19668 26367
rect 19616 26324 19668 26333
rect 19800 26324 19852 26376
rect 20444 26367 20496 26376
rect 20444 26333 20453 26367
rect 20453 26333 20487 26367
rect 20487 26333 20496 26367
rect 20444 26324 20496 26333
rect 21180 26367 21232 26376
rect 21180 26333 21189 26367
rect 21189 26333 21223 26367
rect 21223 26333 21232 26367
rect 21180 26324 21232 26333
rect 20076 26256 20128 26308
rect 25412 26324 25464 26376
rect 26700 26324 26752 26376
rect 10784 26188 10836 26240
rect 11428 26188 11480 26240
rect 14004 26188 14056 26240
rect 15384 26188 15436 26240
rect 15936 26188 15988 26240
rect 17684 26188 17736 26240
rect 19248 26188 19300 26240
rect 22376 26256 22428 26308
rect 24492 26256 24544 26308
rect 25504 26256 25556 26308
rect 22284 26188 22336 26240
rect 22744 26188 22796 26240
rect 24032 26188 24084 26240
rect 9935 26086 9987 26138
rect 9999 26086 10051 26138
rect 10063 26086 10115 26138
rect 10127 26086 10179 26138
rect 10191 26086 10243 26138
rect 18920 26086 18972 26138
rect 18984 26086 19036 26138
rect 19048 26086 19100 26138
rect 19112 26086 19164 26138
rect 19176 26086 19228 26138
rect 4804 25984 4856 26036
rect 4068 25848 4120 25900
rect 4160 25891 4212 25900
rect 4160 25857 4169 25891
rect 4169 25857 4203 25891
rect 4203 25857 4212 25891
rect 4160 25848 4212 25857
rect 4528 25891 4580 25900
rect 4528 25857 4537 25891
rect 4537 25857 4571 25891
rect 4571 25857 4580 25891
rect 5264 25916 5316 25968
rect 7196 25984 7248 26036
rect 7840 25984 7892 26036
rect 8668 26027 8720 26036
rect 8668 25993 8677 26027
rect 8677 25993 8711 26027
rect 8711 25993 8720 26027
rect 8668 25984 8720 25993
rect 4528 25848 4580 25857
rect 5448 25848 5500 25900
rect 7472 25916 7524 25968
rect 10876 25984 10928 26036
rect 11520 25984 11572 26036
rect 12440 25984 12492 26036
rect 1400 25780 1452 25832
rect 1860 25823 1912 25832
rect 1860 25789 1869 25823
rect 1869 25789 1903 25823
rect 1903 25789 1912 25823
rect 1860 25780 1912 25789
rect 4436 25780 4488 25832
rect 4620 25780 4672 25832
rect 7564 25848 7616 25900
rect 8852 25891 8904 25900
rect 8852 25857 8861 25891
rect 8861 25857 8895 25891
rect 8895 25857 8904 25891
rect 8852 25848 8904 25857
rect 9588 25891 9640 25900
rect 9588 25857 9597 25891
rect 9597 25857 9631 25891
rect 9631 25857 9640 25891
rect 9588 25848 9640 25857
rect 9680 25891 9732 25900
rect 9680 25857 9689 25891
rect 9689 25857 9723 25891
rect 9723 25857 9732 25891
rect 9680 25848 9732 25857
rect 6828 25712 6880 25764
rect 8852 25712 8904 25764
rect 10784 25916 10836 25968
rect 12440 25848 12492 25900
rect 12808 25984 12860 26036
rect 13820 25984 13872 26036
rect 14096 26027 14148 26036
rect 14096 25993 14105 26027
rect 14105 25993 14139 26027
rect 14139 25993 14148 26027
rect 14096 25984 14148 25993
rect 12624 25916 12676 25968
rect 17500 25984 17552 26036
rect 14280 25916 14332 25968
rect 12992 25891 13044 25900
rect 12992 25857 13001 25891
rect 13001 25857 13035 25891
rect 13035 25857 13044 25891
rect 12992 25848 13044 25857
rect 13268 25891 13320 25900
rect 13268 25857 13277 25891
rect 13277 25857 13311 25891
rect 13311 25857 13320 25891
rect 13268 25848 13320 25857
rect 13912 25891 13964 25900
rect 13912 25857 13921 25891
rect 13921 25857 13955 25891
rect 13955 25857 13964 25891
rect 13912 25848 13964 25857
rect 18696 25916 18748 25968
rect 15844 25848 15896 25900
rect 14004 25780 14056 25832
rect 17684 25848 17736 25900
rect 17960 25891 18012 25900
rect 17960 25857 17969 25891
rect 17969 25857 18003 25891
rect 18003 25857 18012 25891
rect 19340 25984 19392 26036
rect 20444 25984 20496 26036
rect 22008 25984 22060 26036
rect 22284 25984 22336 26036
rect 17960 25848 18012 25857
rect 19248 25848 19300 25900
rect 20904 25916 20956 25968
rect 22100 25959 22152 25968
rect 22100 25925 22109 25959
rect 22109 25925 22143 25959
rect 22143 25925 22152 25959
rect 22100 25916 22152 25925
rect 22744 25916 22796 25968
rect 24032 25984 24084 26036
rect 24584 26027 24636 26036
rect 24584 25993 24593 26027
rect 24593 25993 24627 26027
rect 24627 25993 24636 26027
rect 24584 25984 24636 25993
rect 26424 25984 26476 26036
rect 18144 25780 18196 25832
rect 18604 25780 18656 25832
rect 19616 25780 19668 25832
rect 19800 25891 19852 25900
rect 19800 25857 19809 25891
rect 19809 25857 19843 25891
rect 19843 25857 19852 25891
rect 19800 25848 19852 25857
rect 19984 25848 20036 25900
rect 20628 25891 20680 25900
rect 20628 25857 20637 25891
rect 20637 25857 20671 25891
rect 20671 25857 20680 25891
rect 20628 25848 20680 25857
rect 21088 25891 21140 25900
rect 21088 25857 21097 25891
rect 21097 25857 21131 25891
rect 21131 25857 21140 25891
rect 21088 25848 21140 25857
rect 21180 25848 21232 25900
rect 21824 25891 21876 25900
rect 21824 25857 21833 25891
rect 21833 25857 21867 25891
rect 21867 25857 21876 25891
rect 21824 25848 21876 25857
rect 21916 25848 21968 25900
rect 23204 25891 23256 25900
rect 20812 25780 20864 25832
rect 1308 25644 1360 25696
rect 1584 25644 1636 25696
rect 4804 25644 4856 25696
rect 4896 25644 4948 25696
rect 6276 25644 6328 25696
rect 6460 25687 6512 25696
rect 6460 25653 6469 25687
rect 6469 25653 6503 25687
rect 6503 25653 6512 25687
rect 6460 25644 6512 25653
rect 7288 25644 7340 25696
rect 9864 25644 9916 25696
rect 12256 25644 12308 25696
rect 13728 25712 13780 25764
rect 17408 25712 17460 25764
rect 18512 25712 18564 25764
rect 14832 25644 14884 25696
rect 15108 25687 15160 25696
rect 15108 25653 15117 25687
rect 15117 25653 15151 25687
rect 15151 25653 15160 25687
rect 15108 25644 15160 25653
rect 15936 25687 15988 25696
rect 15936 25653 15945 25687
rect 15945 25653 15979 25687
rect 15979 25653 15988 25687
rect 15936 25644 15988 25653
rect 16488 25644 16540 25696
rect 19800 25644 19852 25696
rect 20536 25644 20588 25696
rect 23204 25857 23213 25891
rect 23213 25857 23247 25891
rect 23247 25857 23256 25891
rect 23204 25848 23256 25857
rect 23296 25848 23348 25900
rect 24124 25916 24176 25968
rect 24952 25848 25004 25900
rect 26424 25848 26476 25900
rect 27160 25891 27212 25900
rect 27160 25857 27169 25891
rect 27169 25857 27203 25891
rect 27203 25857 27212 25891
rect 27160 25848 27212 25857
rect 24216 25823 24268 25832
rect 24216 25789 24225 25823
rect 24225 25789 24259 25823
rect 24259 25789 24268 25823
rect 24216 25780 24268 25789
rect 26148 25780 26200 25832
rect 22284 25644 22336 25696
rect 24860 25644 24912 25696
rect 26792 25644 26844 25696
rect 5442 25542 5494 25594
rect 5506 25542 5558 25594
rect 5570 25542 5622 25594
rect 5634 25542 5686 25594
rect 5698 25542 5750 25594
rect 14428 25542 14480 25594
rect 14492 25542 14544 25594
rect 14556 25542 14608 25594
rect 14620 25542 14672 25594
rect 14684 25542 14736 25594
rect 23413 25542 23465 25594
rect 23477 25542 23529 25594
rect 23541 25542 23593 25594
rect 23605 25542 23657 25594
rect 23669 25542 23721 25594
rect 2964 25440 3016 25492
rect 4068 25440 4120 25492
rect 4620 25440 4672 25492
rect 5172 25440 5224 25492
rect 9588 25440 9640 25492
rect 12440 25483 12492 25492
rect 12440 25449 12449 25483
rect 12449 25449 12483 25483
rect 12483 25449 12492 25483
rect 12440 25440 12492 25449
rect 4160 25372 4212 25424
rect 7472 25372 7524 25424
rect 8024 25372 8076 25424
rect 10324 25372 10376 25424
rect 4804 25347 4856 25356
rect 4804 25313 4813 25347
rect 4813 25313 4847 25347
rect 4847 25313 4856 25347
rect 4804 25304 4856 25313
rect 3240 25279 3292 25288
rect 3240 25245 3249 25279
rect 3249 25245 3283 25279
rect 3283 25245 3292 25279
rect 3240 25236 3292 25245
rect 5908 25304 5960 25356
rect 5080 25279 5132 25288
rect 3332 25168 3384 25220
rect 5080 25245 5089 25279
rect 5089 25245 5123 25279
rect 5123 25245 5132 25279
rect 5080 25236 5132 25245
rect 5724 25279 5776 25288
rect 5724 25245 5733 25279
rect 5733 25245 5767 25279
rect 5767 25245 5776 25279
rect 5724 25236 5776 25245
rect 6092 25236 6144 25288
rect 6828 25279 6880 25288
rect 6828 25245 6837 25279
rect 6837 25245 6871 25279
rect 6871 25245 6880 25279
rect 6828 25236 6880 25245
rect 9404 25279 9456 25288
rect 9404 25245 9413 25279
rect 9413 25245 9447 25279
rect 9447 25245 9456 25279
rect 9404 25236 9456 25245
rect 12440 25304 12492 25356
rect 12992 25440 13044 25492
rect 13084 25440 13136 25492
rect 14280 25372 14332 25424
rect 12808 25347 12860 25356
rect 12808 25313 12817 25347
rect 12817 25313 12851 25347
rect 12851 25313 12860 25347
rect 12808 25304 12860 25313
rect 15108 25440 15160 25492
rect 14832 25372 14884 25424
rect 15292 25372 15344 25424
rect 16304 25372 16356 25424
rect 19616 25440 19668 25492
rect 22468 25440 22520 25492
rect 24952 25483 25004 25492
rect 24952 25449 24961 25483
rect 24961 25449 24995 25483
rect 24995 25449 25004 25483
rect 24952 25440 25004 25449
rect 17868 25372 17920 25424
rect 17960 25304 18012 25356
rect 6368 25168 6420 25220
rect 7564 25168 7616 25220
rect 3056 25143 3108 25152
rect 3056 25109 3065 25143
rect 3065 25109 3099 25143
rect 3099 25109 3108 25143
rect 3056 25100 3108 25109
rect 4252 25100 4304 25152
rect 4712 25100 4764 25152
rect 5356 25100 5408 25152
rect 10968 25236 11020 25288
rect 11796 25236 11848 25288
rect 12900 25279 12952 25288
rect 10876 25168 10928 25220
rect 12900 25245 12909 25279
rect 12909 25245 12943 25279
rect 12943 25245 12952 25279
rect 12900 25236 12952 25245
rect 13268 25236 13320 25288
rect 15844 25236 15896 25288
rect 16396 25236 16448 25288
rect 22744 25372 22796 25424
rect 20352 25347 20404 25356
rect 20352 25313 20361 25347
rect 20361 25313 20395 25347
rect 20395 25313 20404 25347
rect 20352 25304 20404 25313
rect 19892 25236 19944 25288
rect 21088 25236 21140 25288
rect 21364 25279 21416 25288
rect 21364 25245 21373 25279
rect 21373 25245 21407 25279
rect 21407 25245 21416 25279
rect 21364 25236 21416 25245
rect 21824 25279 21876 25288
rect 21824 25245 21833 25279
rect 21833 25245 21867 25279
rect 21867 25245 21876 25279
rect 21824 25236 21876 25245
rect 22284 25304 22336 25356
rect 24124 25304 24176 25356
rect 25412 25347 25464 25356
rect 22744 25236 22796 25288
rect 24400 25279 24452 25288
rect 24400 25245 24409 25279
rect 24409 25245 24443 25279
rect 24443 25245 24452 25279
rect 24400 25236 24452 25245
rect 24584 25279 24636 25288
rect 24584 25245 24593 25279
rect 24593 25245 24627 25279
rect 24627 25245 24636 25279
rect 24584 25236 24636 25245
rect 25412 25313 25421 25347
rect 25421 25313 25455 25347
rect 25455 25313 25464 25347
rect 25412 25304 25464 25313
rect 24952 25236 25004 25288
rect 26240 25236 26292 25288
rect 14188 25211 14240 25220
rect 14188 25177 14197 25211
rect 14197 25177 14231 25211
rect 14231 25177 14240 25211
rect 14188 25168 14240 25177
rect 16856 25168 16908 25220
rect 20812 25168 20864 25220
rect 22008 25211 22060 25220
rect 22008 25177 22017 25211
rect 22017 25177 22051 25211
rect 22051 25177 22060 25211
rect 22008 25168 22060 25177
rect 22468 25168 22520 25220
rect 24676 25211 24728 25220
rect 24676 25177 24681 25211
rect 24681 25177 24715 25211
rect 24715 25177 24728 25211
rect 24676 25168 24728 25177
rect 10968 25100 11020 25152
rect 15200 25100 15252 25152
rect 16948 25143 17000 25152
rect 16948 25109 16957 25143
rect 16957 25109 16991 25143
rect 16991 25109 17000 25143
rect 16948 25100 17000 25109
rect 20168 25143 20220 25152
rect 20168 25109 20177 25143
rect 20177 25109 20211 25143
rect 20211 25109 20220 25143
rect 20168 25100 20220 25109
rect 21732 25100 21784 25152
rect 23020 25100 23072 25152
rect 9935 24998 9987 25050
rect 9999 24998 10051 25050
rect 10063 24998 10115 25050
rect 10127 24998 10179 25050
rect 10191 24998 10243 25050
rect 18920 24998 18972 25050
rect 18984 24998 19036 25050
rect 19048 24998 19100 25050
rect 19112 24998 19164 25050
rect 19176 24998 19228 25050
rect 2412 24803 2464 24812
rect 2412 24769 2421 24803
rect 2421 24769 2455 24803
rect 2455 24769 2464 24803
rect 2412 24760 2464 24769
rect 3516 24828 3568 24880
rect 3976 24828 4028 24880
rect 1308 24692 1360 24744
rect 4068 24760 4120 24812
rect 5816 24896 5868 24948
rect 6460 24896 6512 24948
rect 9312 24896 9364 24948
rect 9772 24896 9824 24948
rect 10876 24939 10928 24948
rect 10876 24905 10885 24939
rect 10885 24905 10919 24939
rect 10919 24905 10928 24939
rect 10876 24896 10928 24905
rect 12440 24896 12492 24948
rect 4804 24828 4856 24880
rect 7472 24871 7524 24880
rect 4896 24760 4948 24812
rect 5540 24803 5592 24812
rect 5540 24769 5549 24803
rect 5549 24769 5583 24803
rect 5583 24769 5592 24803
rect 5540 24760 5592 24769
rect 5724 24803 5776 24812
rect 5724 24769 5733 24803
rect 5733 24769 5767 24803
rect 5767 24769 5776 24803
rect 5724 24760 5776 24769
rect 5908 24760 5960 24812
rect 7472 24837 7481 24871
rect 7481 24837 7515 24871
rect 7515 24837 7524 24871
rect 7472 24828 7524 24837
rect 7656 24803 7708 24812
rect 3424 24692 3476 24744
rect 2412 24624 2464 24676
rect 3148 24624 3200 24676
rect 3700 24692 3752 24744
rect 5632 24692 5684 24744
rect 6184 24692 6236 24744
rect 6460 24735 6512 24744
rect 6460 24701 6469 24735
rect 6469 24701 6503 24735
rect 6503 24701 6512 24735
rect 6460 24692 6512 24701
rect 3792 24624 3844 24676
rect 6092 24624 6144 24676
rect 7656 24769 7665 24803
rect 7665 24769 7699 24803
rect 7699 24769 7708 24803
rect 7656 24760 7708 24769
rect 7748 24803 7800 24812
rect 7748 24769 7757 24803
rect 7757 24769 7791 24803
rect 7791 24769 7800 24803
rect 7748 24760 7800 24769
rect 8760 24760 8812 24812
rect 9588 24803 9640 24812
rect 6920 24692 6972 24744
rect 1952 24556 2004 24608
rect 2964 24556 3016 24608
rect 3424 24599 3476 24608
rect 3424 24565 3433 24599
rect 3433 24565 3467 24599
rect 3467 24565 3476 24599
rect 3424 24556 3476 24565
rect 3700 24556 3752 24608
rect 4160 24556 4212 24608
rect 6184 24556 6236 24608
rect 7840 24624 7892 24676
rect 8484 24735 8536 24744
rect 8484 24701 8493 24735
rect 8493 24701 8527 24735
rect 8527 24701 8536 24735
rect 9588 24769 9597 24803
rect 9597 24769 9631 24803
rect 9631 24769 9640 24803
rect 9588 24760 9640 24769
rect 8484 24692 8536 24701
rect 9680 24692 9732 24744
rect 10324 24760 10376 24812
rect 10784 24803 10836 24812
rect 10784 24769 10793 24803
rect 10793 24769 10827 24803
rect 10827 24769 10836 24803
rect 10784 24760 10836 24769
rect 10876 24760 10928 24812
rect 11152 24760 11204 24812
rect 12624 24828 12676 24880
rect 13084 24896 13136 24948
rect 18696 24939 18748 24948
rect 18696 24905 18705 24939
rect 18705 24905 18739 24939
rect 18739 24905 18748 24939
rect 18696 24896 18748 24905
rect 12072 24760 12124 24812
rect 12348 24803 12400 24812
rect 10692 24692 10744 24744
rect 12348 24769 12357 24803
rect 12357 24769 12391 24803
rect 12391 24769 12400 24803
rect 12348 24760 12400 24769
rect 13544 24760 13596 24812
rect 14188 24760 14240 24812
rect 15200 24803 15252 24812
rect 15200 24769 15209 24803
rect 15209 24769 15243 24803
rect 15243 24769 15252 24803
rect 15200 24760 15252 24769
rect 12624 24692 12676 24744
rect 12808 24692 12860 24744
rect 6920 24556 6972 24608
rect 9864 24624 9916 24676
rect 12072 24624 12124 24676
rect 12256 24667 12308 24676
rect 12256 24633 12265 24667
rect 12265 24633 12299 24667
rect 12299 24633 12308 24667
rect 12256 24624 12308 24633
rect 13176 24667 13228 24676
rect 13176 24633 13185 24667
rect 13185 24633 13219 24667
rect 13219 24633 13228 24667
rect 13176 24624 13228 24633
rect 17500 24760 17552 24812
rect 17684 24803 17736 24812
rect 17684 24769 17693 24803
rect 17693 24769 17727 24803
rect 17727 24769 17736 24803
rect 17684 24760 17736 24769
rect 15384 24624 15436 24676
rect 11520 24556 11572 24608
rect 12348 24556 12400 24608
rect 12900 24556 12952 24608
rect 13636 24556 13688 24608
rect 13912 24556 13964 24608
rect 15660 24556 15712 24608
rect 16856 24556 16908 24608
rect 17224 24692 17276 24744
rect 18604 24828 18656 24880
rect 19524 24896 19576 24948
rect 20352 24896 20404 24948
rect 21180 24896 21232 24948
rect 22008 24939 22060 24948
rect 22008 24905 22017 24939
rect 22017 24905 22051 24939
rect 22051 24905 22060 24939
rect 22008 24896 22060 24905
rect 18236 24760 18288 24812
rect 22468 24871 22520 24880
rect 20076 24760 20128 24812
rect 19248 24735 19300 24744
rect 19248 24701 19257 24735
rect 19257 24701 19291 24735
rect 19291 24701 19300 24735
rect 19248 24692 19300 24701
rect 21180 24760 21232 24812
rect 22468 24837 22477 24871
rect 22477 24837 22511 24871
rect 22511 24837 22520 24871
rect 22468 24828 22520 24837
rect 23204 24828 23256 24880
rect 22376 24803 22428 24812
rect 22376 24769 22385 24803
rect 22385 24769 22419 24803
rect 22419 24769 22428 24803
rect 22376 24760 22428 24769
rect 22560 24760 22612 24812
rect 20536 24735 20588 24744
rect 20536 24701 20545 24735
rect 20545 24701 20579 24735
rect 20579 24701 20588 24735
rect 20536 24692 20588 24701
rect 23204 24692 23256 24744
rect 24400 24760 24452 24812
rect 24768 24803 24820 24812
rect 24768 24769 24777 24803
rect 24777 24769 24811 24803
rect 24811 24769 24820 24803
rect 24768 24760 24820 24769
rect 23848 24692 23900 24744
rect 24952 24803 25004 24812
rect 24952 24769 24961 24803
rect 24961 24769 24995 24803
rect 24995 24769 25004 24803
rect 24952 24760 25004 24769
rect 25044 24692 25096 24744
rect 26240 24760 26292 24812
rect 19432 24556 19484 24608
rect 21088 24599 21140 24608
rect 21088 24565 21097 24599
rect 21097 24565 21131 24599
rect 21131 24565 21140 24599
rect 21088 24556 21140 24565
rect 21272 24624 21324 24676
rect 27988 24760 28040 24812
rect 24952 24556 25004 24608
rect 25320 24556 25372 24608
rect 25596 24599 25648 24608
rect 25596 24565 25605 24599
rect 25605 24565 25639 24599
rect 25639 24565 25648 24599
rect 25596 24556 25648 24565
rect 27068 24556 27120 24608
rect 27528 24556 27580 24608
rect 5442 24454 5494 24506
rect 5506 24454 5558 24506
rect 5570 24454 5622 24506
rect 5634 24454 5686 24506
rect 5698 24454 5750 24506
rect 14428 24454 14480 24506
rect 14492 24454 14544 24506
rect 14556 24454 14608 24506
rect 14620 24454 14672 24506
rect 14684 24454 14736 24506
rect 23413 24454 23465 24506
rect 23477 24454 23529 24506
rect 23541 24454 23593 24506
rect 23605 24454 23657 24506
rect 23669 24454 23721 24506
rect 204 24352 256 24404
rect 3240 24352 3292 24404
rect 3516 24352 3568 24404
rect 5264 24352 5316 24404
rect 5908 24395 5960 24404
rect 5908 24361 5917 24395
rect 5917 24361 5951 24395
rect 5951 24361 5960 24395
rect 5908 24352 5960 24361
rect 7748 24352 7800 24404
rect 8300 24352 8352 24404
rect 10784 24352 10836 24404
rect 12532 24352 12584 24404
rect 14832 24395 14884 24404
rect 14832 24361 14841 24395
rect 14841 24361 14875 24395
rect 14875 24361 14884 24395
rect 14832 24352 14884 24361
rect 17224 24352 17276 24404
rect 17776 24352 17828 24404
rect 18788 24352 18840 24404
rect 19432 24352 19484 24404
rect 20720 24352 20772 24404
rect 21916 24352 21968 24404
rect 22560 24352 22612 24404
rect 22744 24352 22796 24404
rect 2964 24284 3016 24336
rect 4528 24284 4580 24336
rect 5816 24284 5868 24336
rect 6184 24284 6236 24336
rect 7656 24284 7708 24336
rect 16856 24284 16908 24336
rect 17684 24284 17736 24336
rect 23296 24352 23348 24404
rect 25504 24395 25556 24404
rect 25504 24361 25513 24395
rect 25513 24361 25547 24395
rect 25547 24361 25556 24395
rect 25504 24352 25556 24361
rect 25964 24352 26016 24404
rect 27160 24352 27212 24404
rect 23388 24284 23440 24336
rect 1400 24259 1452 24268
rect 1400 24225 1409 24259
rect 1409 24225 1443 24259
rect 1443 24225 1452 24259
rect 1400 24216 1452 24225
rect 3148 24216 3200 24268
rect 4712 24216 4764 24268
rect 5356 24259 5408 24268
rect 5356 24225 5365 24259
rect 5365 24225 5399 24259
rect 5399 24225 5408 24259
rect 5356 24216 5408 24225
rect 6920 24216 6972 24268
rect 8116 24216 8168 24268
rect 8484 24216 8536 24268
rect 9864 24216 9916 24268
rect 10968 24216 11020 24268
rect 15844 24259 15896 24268
rect 15844 24225 15853 24259
rect 15853 24225 15887 24259
rect 15887 24225 15896 24259
rect 15844 24216 15896 24225
rect 17224 24259 17276 24268
rect 17224 24225 17233 24259
rect 17233 24225 17267 24259
rect 17267 24225 17276 24259
rect 17224 24216 17276 24225
rect 3792 24191 3844 24200
rect 3792 24157 3801 24191
rect 3801 24157 3835 24191
rect 3835 24157 3844 24191
rect 3792 24148 3844 24157
rect 3976 24191 4028 24200
rect 3976 24157 3985 24191
rect 3985 24157 4019 24191
rect 4019 24157 4028 24191
rect 3976 24148 4028 24157
rect 6368 24148 6420 24200
rect 7932 24148 7984 24200
rect 8024 24148 8076 24200
rect 3240 24080 3292 24132
rect 4620 24080 4672 24132
rect 5080 24123 5132 24132
rect 5080 24089 5089 24123
rect 5089 24089 5123 24123
rect 5123 24089 5132 24123
rect 5080 24080 5132 24089
rect 6644 24080 6696 24132
rect 2964 24012 3016 24064
rect 4068 24012 4120 24064
rect 4252 24012 4304 24064
rect 5908 24012 5960 24064
rect 6368 24055 6420 24064
rect 6368 24021 6377 24055
rect 6377 24021 6411 24055
rect 6411 24021 6420 24055
rect 6368 24012 6420 24021
rect 7840 24012 7892 24064
rect 8300 24012 8352 24064
rect 9036 24148 9088 24200
rect 9956 24148 10008 24200
rect 10140 24191 10192 24200
rect 10140 24157 10149 24191
rect 10149 24157 10183 24191
rect 10183 24157 10192 24191
rect 10416 24191 10468 24200
rect 10140 24148 10192 24157
rect 10416 24157 10425 24191
rect 10425 24157 10459 24191
rect 10459 24157 10468 24191
rect 10416 24148 10468 24157
rect 11152 24191 11204 24200
rect 11152 24157 11161 24191
rect 11161 24157 11195 24191
rect 11195 24157 11204 24191
rect 11152 24148 11204 24157
rect 11704 24148 11756 24200
rect 13176 24191 13228 24200
rect 11612 24080 11664 24132
rect 9588 24012 9640 24064
rect 12624 24080 12676 24132
rect 13176 24157 13185 24191
rect 13185 24157 13219 24191
rect 13219 24157 13228 24191
rect 13176 24148 13228 24157
rect 14188 24148 14240 24200
rect 14740 24191 14792 24200
rect 14740 24157 14749 24191
rect 14749 24157 14783 24191
rect 14783 24157 14792 24191
rect 14740 24148 14792 24157
rect 15200 24148 15252 24200
rect 16672 24148 16724 24200
rect 16948 24148 17000 24200
rect 18236 24191 18288 24200
rect 13268 24055 13320 24064
rect 13268 24021 13277 24055
rect 13277 24021 13311 24055
rect 13311 24021 13320 24055
rect 13268 24012 13320 24021
rect 15936 24080 15988 24132
rect 18236 24157 18245 24191
rect 18245 24157 18279 24191
rect 18279 24157 18288 24191
rect 18236 24148 18288 24157
rect 19616 24216 19668 24268
rect 19800 24259 19852 24268
rect 19800 24225 19809 24259
rect 19809 24225 19843 24259
rect 19843 24225 19852 24259
rect 19800 24216 19852 24225
rect 20168 24216 20220 24268
rect 21640 24259 21692 24268
rect 19524 24148 19576 24200
rect 20444 24148 20496 24200
rect 21640 24225 21649 24259
rect 21649 24225 21683 24259
rect 21683 24225 21692 24259
rect 21640 24216 21692 24225
rect 22560 24216 22612 24268
rect 22744 24216 22796 24268
rect 25412 24216 25464 24268
rect 25964 24259 26016 24268
rect 25964 24225 25973 24259
rect 25973 24225 26007 24259
rect 26007 24225 26016 24259
rect 25964 24216 26016 24225
rect 21916 24148 21968 24200
rect 24492 24148 24544 24200
rect 25320 24191 25372 24200
rect 17500 24080 17552 24132
rect 21272 24080 21324 24132
rect 21456 24123 21508 24132
rect 21456 24089 21465 24123
rect 21465 24089 21499 24123
rect 21499 24089 21508 24123
rect 21456 24080 21508 24089
rect 21824 24080 21876 24132
rect 22836 24080 22888 24132
rect 24124 24080 24176 24132
rect 25320 24157 25329 24191
rect 25329 24157 25363 24191
rect 25363 24157 25372 24191
rect 25320 24148 25372 24157
rect 26516 24148 26568 24200
rect 26148 24080 26200 24132
rect 15108 24012 15160 24064
rect 18236 24012 18288 24064
rect 18420 24012 18472 24064
rect 19340 24012 19392 24064
rect 20260 24012 20312 24064
rect 20720 24012 20772 24064
rect 21916 24012 21968 24064
rect 22284 24055 22336 24064
rect 22284 24021 22293 24055
rect 22293 24021 22327 24055
rect 22327 24021 22336 24055
rect 22284 24012 22336 24021
rect 22376 24012 22428 24064
rect 23388 24055 23440 24064
rect 23388 24021 23397 24055
rect 23397 24021 23431 24055
rect 23431 24021 23440 24055
rect 23388 24012 23440 24021
rect 24032 24012 24084 24064
rect 25044 24012 25096 24064
rect 25504 24012 25556 24064
rect 9935 23910 9987 23962
rect 9999 23910 10051 23962
rect 10063 23910 10115 23962
rect 10127 23910 10179 23962
rect 10191 23910 10243 23962
rect 18920 23910 18972 23962
rect 18984 23910 19036 23962
rect 19048 23910 19100 23962
rect 19112 23910 19164 23962
rect 19176 23910 19228 23962
rect 4252 23808 4304 23860
rect 5356 23808 5408 23860
rect 2136 23715 2188 23724
rect 2136 23681 2145 23715
rect 2145 23681 2179 23715
rect 2179 23681 2188 23715
rect 2136 23672 2188 23681
rect 3424 23715 3476 23724
rect 3424 23681 3433 23715
rect 3433 23681 3467 23715
rect 3467 23681 3476 23715
rect 3424 23672 3476 23681
rect 3608 23647 3660 23656
rect 3608 23613 3617 23647
rect 3617 23613 3651 23647
rect 3651 23613 3660 23647
rect 3608 23604 3660 23613
rect 6092 23808 6144 23860
rect 7012 23808 7064 23860
rect 7656 23808 7708 23860
rect 7840 23808 7892 23860
rect 8944 23808 8996 23860
rect 9220 23808 9272 23860
rect 4068 23672 4120 23724
rect 5264 23672 5316 23724
rect 3240 23536 3292 23588
rect 2780 23511 2832 23520
rect 2780 23477 2789 23511
rect 2789 23477 2823 23511
rect 2823 23477 2832 23511
rect 2780 23468 2832 23477
rect 3608 23468 3660 23520
rect 4436 23468 4488 23520
rect 5356 23604 5408 23656
rect 7288 23672 7340 23724
rect 8208 23740 8260 23792
rect 8392 23740 8444 23792
rect 9036 23740 9088 23792
rect 9128 23740 9180 23792
rect 7564 23672 7616 23724
rect 6920 23604 6972 23656
rect 7656 23604 7708 23656
rect 7932 23604 7984 23656
rect 9588 23715 9640 23724
rect 9588 23681 9597 23715
rect 9597 23681 9631 23715
rect 9631 23681 9640 23715
rect 9588 23672 9640 23681
rect 10416 23740 10468 23792
rect 11152 23740 11204 23792
rect 11612 23808 11664 23860
rect 10784 23715 10836 23724
rect 8944 23647 8996 23656
rect 8944 23613 8953 23647
rect 8953 23613 8987 23647
rect 8987 23613 8996 23647
rect 8944 23604 8996 23613
rect 9128 23647 9180 23656
rect 9128 23613 9137 23647
rect 9137 23613 9171 23647
rect 9171 23613 9180 23647
rect 9128 23604 9180 23613
rect 9312 23604 9364 23656
rect 10784 23681 10793 23715
rect 10793 23681 10827 23715
rect 10827 23681 10836 23715
rect 10784 23672 10836 23681
rect 13728 23808 13780 23860
rect 15660 23851 15712 23860
rect 15660 23817 15685 23851
rect 15685 23817 15712 23851
rect 15660 23808 15712 23817
rect 17868 23808 17920 23860
rect 19248 23808 19300 23860
rect 20536 23808 20588 23860
rect 22560 23808 22612 23860
rect 23204 23851 23256 23860
rect 15384 23740 15436 23792
rect 18512 23783 18564 23792
rect 18512 23749 18521 23783
rect 18521 23749 18555 23783
rect 18555 23749 18564 23783
rect 18512 23740 18564 23749
rect 19156 23740 19208 23792
rect 23204 23817 23213 23851
rect 23213 23817 23247 23851
rect 23247 23817 23256 23851
rect 23204 23808 23256 23817
rect 24768 23808 24820 23860
rect 12532 23715 12584 23724
rect 12532 23681 12566 23715
rect 12566 23681 12584 23715
rect 10232 23604 10284 23656
rect 10600 23604 10652 23656
rect 12532 23672 12584 23681
rect 13544 23672 13596 23724
rect 14740 23672 14792 23724
rect 17224 23715 17276 23724
rect 17224 23681 17233 23715
rect 17233 23681 17267 23715
rect 17267 23681 17276 23715
rect 17224 23672 17276 23681
rect 11704 23604 11756 23656
rect 11888 23604 11940 23656
rect 8024 23536 8076 23588
rect 8484 23468 8536 23520
rect 9036 23511 9088 23520
rect 9036 23477 9045 23511
rect 9045 23477 9079 23511
rect 9079 23477 9088 23511
rect 9036 23468 9088 23477
rect 11520 23468 11572 23520
rect 16672 23604 16724 23656
rect 18512 23604 18564 23656
rect 18696 23647 18748 23656
rect 18696 23613 18705 23647
rect 18705 23613 18739 23647
rect 18739 23613 18748 23647
rect 18696 23604 18748 23613
rect 14280 23536 14332 23588
rect 19524 23672 19576 23724
rect 19708 23672 19760 23724
rect 19892 23672 19944 23724
rect 19248 23604 19300 23656
rect 21640 23672 21692 23724
rect 19524 23536 19576 23588
rect 13728 23468 13780 23520
rect 14004 23468 14056 23520
rect 16948 23468 17000 23520
rect 18052 23468 18104 23520
rect 18236 23468 18288 23520
rect 20904 23604 20956 23656
rect 21916 23647 21968 23656
rect 21916 23613 21925 23647
rect 21925 23613 21959 23647
rect 21959 23613 21968 23647
rect 21916 23604 21968 23613
rect 21180 23536 21232 23588
rect 22008 23511 22060 23520
rect 22008 23477 22017 23511
rect 22017 23477 22051 23511
rect 22051 23477 22060 23511
rect 22008 23468 22060 23477
rect 25320 23740 25372 23792
rect 22376 23672 22428 23724
rect 23112 23672 23164 23724
rect 23388 23672 23440 23724
rect 24768 23672 24820 23724
rect 25688 23808 25740 23860
rect 25504 23783 25556 23792
rect 25504 23749 25513 23783
rect 25513 23749 25547 23783
rect 25547 23749 25556 23783
rect 27160 23783 27212 23792
rect 25504 23740 25556 23749
rect 27160 23749 27169 23783
rect 27169 23749 27203 23783
rect 27203 23749 27212 23783
rect 27160 23740 27212 23749
rect 23296 23604 23348 23656
rect 24400 23604 24452 23656
rect 25596 23647 25648 23656
rect 25596 23613 25605 23647
rect 25605 23613 25639 23647
rect 25639 23613 25648 23647
rect 25596 23604 25648 23613
rect 25688 23536 25740 23588
rect 27436 23536 27488 23588
rect 22560 23468 22612 23520
rect 25320 23468 25372 23520
rect 5442 23366 5494 23418
rect 5506 23366 5558 23418
rect 5570 23366 5622 23418
rect 5634 23366 5686 23418
rect 5698 23366 5750 23418
rect 14428 23366 14480 23418
rect 14492 23366 14544 23418
rect 14556 23366 14608 23418
rect 14620 23366 14672 23418
rect 14684 23366 14736 23418
rect 23413 23366 23465 23418
rect 23477 23366 23529 23418
rect 23541 23366 23593 23418
rect 23605 23366 23657 23418
rect 23669 23366 23721 23418
rect 3792 23264 3844 23316
rect 5908 23307 5960 23316
rect 5908 23273 5917 23307
rect 5917 23273 5951 23307
rect 5951 23273 5960 23307
rect 5908 23264 5960 23273
rect 6368 23264 6420 23316
rect 6920 23264 6972 23316
rect 10784 23264 10836 23316
rect 12532 23264 12584 23316
rect 13728 23264 13780 23316
rect 5356 23196 5408 23248
rect 6460 23196 6512 23248
rect 7564 23196 7616 23248
rect 7932 23196 7984 23248
rect 8484 23196 8536 23248
rect 8852 23196 8904 23248
rect 4436 23128 4488 23180
rect 2044 22924 2096 22976
rect 2964 23060 3016 23112
rect 3148 23060 3200 23112
rect 4252 23060 4304 23112
rect 5080 23060 5132 23112
rect 7840 23128 7892 23180
rect 7196 23060 7248 23112
rect 7656 23103 7708 23112
rect 7656 23069 7665 23103
rect 7665 23069 7699 23103
rect 7699 23069 7708 23103
rect 7656 23060 7708 23069
rect 8024 23103 8076 23112
rect 8024 23069 8033 23103
rect 8033 23069 8067 23103
rect 8067 23069 8076 23103
rect 8024 23060 8076 23069
rect 8116 23103 8168 23112
rect 8116 23069 8125 23103
rect 8125 23069 8159 23103
rect 8159 23069 8168 23103
rect 9220 23128 9272 23180
rect 10692 23196 10744 23248
rect 16396 23264 16448 23316
rect 18052 23264 18104 23316
rect 20628 23264 20680 23316
rect 22008 23264 22060 23316
rect 22560 23307 22612 23316
rect 22560 23273 22569 23307
rect 22569 23273 22603 23307
rect 22603 23273 22612 23307
rect 22560 23264 22612 23273
rect 22744 23307 22796 23316
rect 22744 23273 22753 23307
rect 22753 23273 22787 23307
rect 22787 23273 22796 23307
rect 22744 23264 22796 23273
rect 22836 23264 22888 23316
rect 24584 23264 24636 23316
rect 9312 23103 9364 23112
rect 8116 23060 8168 23069
rect 9312 23069 9321 23103
rect 9321 23069 9355 23103
rect 9355 23069 9364 23103
rect 9312 23060 9364 23069
rect 9588 23060 9640 23112
rect 10508 23128 10560 23180
rect 10876 23128 10928 23180
rect 9864 23060 9916 23112
rect 11060 23103 11112 23112
rect 4988 23035 5040 23044
rect 4988 23001 4997 23035
rect 4997 23001 5031 23035
rect 5031 23001 5040 23035
rect 4988 22992 5040 23001
rect 5356 22992 5408 23044
rect 7564 22992 7616 23044
rect 8576 22992 8628 23044
rect 8852 22992 8904 23044
rect 9036 22992 9088 23044
rect 11060 23069 11069 23103
rect 11069 23069 11103 23103
rect 11103 23069 11112 23103
rect 11060 23060 11112 23069
rect 11520 23103 11572 23112
rect 11520 23069 11529 23103
rect 11529 23069 11563 23103
rect 11563 23069 11572 23103
rect 11520 23060 11572 23069
rect 11704 23103 11756 23112
rect 11704 23069 11713 23103
rect 11713 23069 11747 23103
rect 11747 23069 11756 23103
rect 11704 23060 11756 23069
rect 12256 23060 12308 23112
rect 12532 23103 12584 23112
rect 12532 23069 12541 23103
rect 12541 23069 12575 23103
rect 12575 23069 12584 23103
rect 14004 23128 14056 23180
rect 18696 23128 18748 23180
rect 19892 23128 19944 23180
rect 12532 23060 12584 23069
rect 13544 23103 13596 23112
rect 13544 23069 13553 23103
rect 13553 23069 13587 23103
rect 13587 23069 13596 23103
rect 13544 23060 13596 23069
rect 14280 23060 14332 23112
rect 15108 23060 15160 23112
rect 15476 23060 15528 23112
rect 15660 23103 15712 23112
rect 15660 23069 15669 23103
rect 15669 23069 15703 23103
rect 15703 23069 15712 23103
rect 15660 23060 15712 23069
rect 16488 23060 16540 23112
rect 16856 23060 16908 23112
rect 18328 23103 18380 23112
rect 18328 23069 18337 23103
rect 18337 23069 18371 23103
rect 18371 23069 18380 23103
rect 18328 23060 18380 23069
rect 18512 23103 18564 23112
rect 18512 23069 18521 23103
rect 18521 23069 18555 23103
rect 18555 23069 18564 23103
rect 18512 23060 18564 23069
rect 19524 23103 19576 23112
rect 12624 22992 12676 23044
rect 14096 23035 14148 23044
rect 14096 23001 14105 23035
rect 14105 23001 14139 23035
rect 14139 23001 14148 23035
rect 14096 22992 14148 23001
rect 2596 22924 2648 22976
rect 2964 22967 3016 22976
rect 2964 22933 2973 22967
rect 2973 22933 3007 22967
rect 3007 22933 3016 22967
rect 2964 22924 3016 22933
rect 3516 22924 3568 22976
rect 3976 22924 4028 22976
rect 5908 22924 5960 22976
rect 7656 22924 7708 22976
rect 12348 22924 12400 22976
rect 13544 22967 13596 22976
rect 13544 22933 13553 22967
rect 13553 22933 13587 22967
rect 13587 22933 13596 22967
rect 13544 22924 13596 22933
rect 14280 22967 14332 22976
rect 14280 22933 14289 22967
rect 14289 22933 14323 22967
rect 14323 22933 14332 22967
rect 14280 22924 14332 22933
rect 14464 22967 14516 22976
rect 14464 22933 14473 22967
rect 14473 22933 14507 22967
rect 14507 22933 14516 22967
rect 14464 22924 14516 22933
rect 19156 22992 19208 23044
rect 19524 23069 19533 23103
rect 19533 23069 19567 23103
rect 19567 23069 19576 23103
rect 19524 23060 19576 23069
rect 19708 22992 19760 23044
rect 20904 23196 20956 23248
rect 21180 23196 21232 23248
rect 21088 23128 21140 23180
rect 20904 23103 20956 23112
rect 20904 23069 20913 23103
rect 20913 23069 20947 23103
rect 20947 23069 20956 23103
rect 20904 23060 20956 23069
rect 21548 23128 21600 23180
rect 21916 23128 21968 23180
rect 22192 23128 22244 23180
rect 23296 23171 23348 23180
rect 23296 23137 23305 23171
rect 23305 23137 23339 23171
rect 23339 23137 23348 23171
rect 23296 23128 23348 23137
rect 25596 23196 25648 23248
rect 25964 23171 26016 23180
rect 25964 23137 25973 23171
rect 25973 23137 26007 23171
rect 26007 23137 26016 23171
rect 25964 23128 26016 23137
rect 21640 23103 21692 23112
rect 21640 23069 21649 23103
rect 21649 23069 21683 23103
rect 21683 23069 21692 23103
rect 21640 23060 21692 23069
rect 21456 22992 21508 23044
rect 23112 23060 23164 23112
rect 24768 23103 24820 23112
rect 24768 23069 24777 23103
rect 24777 23069 24811 23103
rect 24811 23069 24820 23103
rect 24768 23060 24820 23069
rect 22376 22992 22428 23044
rect 23388 22992 23440 23044
rect 26332 22992 26384 23044
rect 19616 22924 19668 22976
rect 22468 22924 22520 22976
rect 24216 22924 24268 22976
rect 24584 22924 24636 22976
rect 25504 22924 25556 22976
rect 9935 22822 9987 22874
rect 9999 22822 10051 22874
rect 10063 22822 10115 22874
rect 10127 22822 10179 22874
rect 10191 22822 10243 22874
rect 18920 22822 18972 22874
rect 18984 22822 19036 22874
rect 19048 22822 19100 22874
rect 19112 22822 19164 22874
rect 19176 22822 19228 22874
rect 2964 22720 3016 22772
rect 3976 22720 4028 22772
rect 3792 22652 3844 22704
rect 4068 22627 4120 22636
rect 4068 22593 4077 22627
rect 4077 22593 4111 22627
rect 4111 22593 4120 22627
rect 4068 22584 4120 22593
rect 5356 22720 5408 22772
rect 6276 22720 6328 22772
rect 6828 22720 6880 22772
rect 7288 22720 7340 22772
rect 8024 22720 8076 22772
rect 8300 22720 8352 22772
rect 4436 22652 4488 22704
rect 7012 22652 7064 22704
rect 5448 22627 5500 22636
rect 4160 22516 4212 22568
rect 4344 22448 4396 22500
rect 4528 22448 4580 22500
rect 5448 22593 5457 22627
rect 5457 22593 5491 22627
rect 5491 22593 5500 22627
rect 5448 22584 5500 22593
rect 7196 22584 7248 22636
rect 7472 22584 7524 22636
rect 9864 22720 9916 22772
rect 11060 22720 11112 22772
rect 12900 22720 12952 22772
rect 17684 22720 17736 22772
rect 17960 22720 18012 22772
rect 18512 22720 18564 22772
rect 18604 22720 18656 22772
rect 19432 22720 19484 22772
rect 19800 22720 19852 22772
rect 20628 22720 20680 22772
rect 20812 22720 20864 22772
rect 21640 22720 21692 22772
rect 22744 22720 22796 22772
rect 24124 22720 24176 22772
rect 24400 22720 24452 22772
rect 25504 22763 25556 22772
rect 25504 22729 25513 22763
rect 25513 22729 25547 22763
rect 25547 22729 25556 22763
rect 25504 22720 25556 22729
rect 26976 22720 27028 22772
rect 6092 22516 6144 22568
rect 6644 22516 6696 22568
rect 6920 22516 6972 22568
rect 9404 22584 9456 22636
rect 9772 22627 9824 22636
rect 9772 22593 9781 22627
rect 9781 22593 9815 22627
rect 9815 22593 9824 22627
rect 9772 22584 9824 22593
rect 11888 22652 11940 22704
rect 8208 22516 8260 22568
rect 8576 22516 8628 22568
rect 10324 22584 10376 22636
rect 10232 22516 10284 22568
rect 10416 22516 10468 22568
rect 10876 22516 10928 22568
rect 5448 22448 5500 22500
rect 7932 22448 7984 22500
rect 2412 22380 2464 22432
rect 4804 22380 4856 22432
rect 4896 22380 4948 22432
rect 5264 22380 5316 22432
rect 6552 22423 6604 22432
rect 6552 22389 6561 22423
rect 6561 22389 6595 22423
rect 6595 22389 6604 22423
rect 6552 22380 6604 22389
rect 7012 22380 7064 22432
rect 7472 22380 7524 22432
rect 8116 22380 8168 22432
rect 8668 22423 8720 22432
rect 8668 22389 8677 22423
rect 8677 22389 8711 22423
rect 8711 22389 8720 22423
rect 8668 22380 8720 22389
rect 9496 22448 9548 22500
rect 11336 22584 11388 22636
rect 12072 22584 12124 22636
rect 13544 22652 13596 22704
rect 15200 22652 15252 22704
rect 15476 22652 15528 22704
rect 12532 22584 12584 22636
rect 14096 22627 14148 22636
rect 14096 22593 14105 22627
rect 14105 22593 14139 22627
rect 14139 22593 14148 22627
rect 14096 22584 14148 22593
rect 14188 22627 14240 22636
rect 14188 22593 14197 22627
rect 14197 22593 14231 22627
rect 14231 22593 14240 22627
rect 14188 22584 14240 22593
rect 14464 22584 14516 22636
rect 15660 22584 15712 22636
rect 19708 22652 19760 22704
rect 20352 22652 20404 22704
rect 22192 22652 22244 22704
rect 22652 22652 22704 22704
rect 25320 22652 25372 22704
rect 12164 22559 12216 22568
rect 12164 22525 12173 22559
rect 12173 22525 12207 22559
rect 12207 22525 12216 22559
rect 12164 22516 12216 22525
rect 12440 22559 12492 22568
rect 12440 22525 12449 22559
rect 12449 22525 12483 22559
rect 12483 22525 12492 22559
rect 12440 22516 12492 22525
rect 12992 22559 13044 22568
rect 12992 22525 13001 22559
rect 13001 22525 13035 22559
rect 13035 22525 13044 22559
rect 12992 22516 13044 22525
rect 16488 22516 16540 22568
rect 17960 22584 18012 22636
rect 18236 22584 18288 22636
rect 19432 22584 19484 22636
rect 21548 22584 21600 22636
rect 22376 22584 22428 22636
rect 22560 22584 22612 22636
rect 23848 22584 23900 22636
rect 27160 22627 27212 22636
rect 27160 22593 27169 22627
rect 27169 22593 27203 22627
rect 27203 22593 27212 22627
rect 27160 22584 27212 22593
rect 16028 22448 16080 22500
rect 14004 22380 14056 22432
rect 16488 22380 16540 22432
rect 19800 22516 19852 22568
rect 20352 22516 20404 22568
rect 20536 22516 20588 22568
rect 20812 22516 20864 22568
rect 23388 22516 23440 22568
rect 25044 22516 25096 22568
rect 25872 22516 25924 22568
rect 26148 22516 26200 22568
rect 26792 22516 26844 22568
rect 18972 22423 19024 22432
rect 18972 22389 18981 22423
rect 18981 22389 19015 22423
rect 19015 22389 19024 22423
rect 18972 22380 19024 22389
rect 19524 22448 19576 22500
rect 20904 22448 20956 22500
rect 21640 22380 21692 22432
rect 22560 22448 22612 22500
rect 23112 22448 23164 22500
rect 23296 22380 23348 22432
rect 25872 22380 25924 22432
rect 5442 22278 5494 22330
rect 5506 22278 5558 22330
rect 5570 22278 5622 22330
rect 5634 22278 5686 22330
rect 5698 22278 5750 22330
rect 14428 22278 14480 22330
rect 14492 22278 14544 22330
rect 14556 22278 14608 22330
rect 14620 22278 14672 22330
rect 14684 22278 14736 22330
rect 23413 22278 23465 22330
rect 23477 22278 23529 22330
rect 23541 22278 23593 22330
rect 23605 22278 23657 22330
rect 23669 22278 23721 22330
rect 4068 22176 4120 22228
rect 3148 22108 3200 22160
rect 4988 22176 5040 22228
rect 5540 22108 5592 22160
rect 2320 21836 2372 21888
rect 2688 21836 2740 21888
rect 3424 21972 3476 22024
rect 3976 21972 4028 22024
rect 4252 22015 4304 22024
rect 4252 21981 4261 22015
rect 4261 21981 4295 22015
rect 4295 21981 4304 22015
rect 4252 21972 4304 21981
rect 4620 22015 4672 22024
rect 4620 21981 4629 22015
rect 4629 21981 4663 22015
rect 4663 21981 4672 22015
rect 4620 21972 4672 21981
rect 6092 22040 6144 22092
rect 5356 22015 5408 22024
rect 5356 21981 5365 22015
rect 5365 21981 5399 22015
rect 5399 21981 5408 22015
rect 5356 21972 5408 21981
rect 5540 22015 5592 22024
rect 5540 21981 5549 22015
rect 5549 21981 5583 22015
rect 5583 21981 5592 22015
rect 8208 22176 8260 22228
rect 8668 22176 8720 22228
rect 7472 22108 7524 22160
rect 5540 21972 5592 21981
rect 4988 21904 5040 21956
rect 5908 21904 5960 21956
rect 6920 22015 6972 22024
rect 6920 21981 6929 22015
rect 6929 21981 6963 22015
rect 6963 21981 6972 22015
rect 7380 22040 7432 22092
rect 9772 22040 9824 22092
rect 10140 22108 10192 22160
rect 6920 21972 6972 21981
rect 7288 21947 7340 21956
rect 7288 21913 7297 21947
rect 7297 21913 7331 21947
rect 7331 21913 7340 21947
rect 7288 21904 7340 21913
rect 7656 21972 7708 22024
rect 8300 21972 8352 22024
rect 8944 22015 8996 22024
rect 8944 21981 8953 22015
rect 8953 21981 8987 22015
rect 8987 21981 8996 22015
rect 8944 21972 8996 21981
rect 9680 22015 9732 22024
rect 9680 21981 9689 22015
rect 9689 21981 9723 22015
rect 9723 21981 9732 22015
rect 9680 21972 9732 21981
rect 10324 22040 10376 22092
rect 10416 22083 10468 22092
rect 10416 22049 10425 22083
rect 10425 22049 10459 22083
rect 10459 22049 10468 22083
rect 10416 22040 10468 22049
rect 12992 22176 13044 22228
rect 14004 22176 14056 22228
rect 14188 22176 14240 22228
rect 12164 22108 12216 22160
rect 11612 22040 11664 22092
rect 11888 22083 11940 22092
rect 11888 22049 11897 22083
rect 11897 22049 11931 22083
rect 11931 22049 11940 22083
rect 11888 22040 11940 22049
rect 14096 22108 14148 22160
rect 14372 22108 14424 22160
rect 18972 22176 19024 22228
rect 19616 22176 19668 22228
rect 18328 22108 18380 22160
rect 20536 22176 20588 22228
rect 25688 22176 25740 22228
rect 26148 22176 26200 22228
rect 27160 22176 27212 22228
rect 23480 22108 23532 22160
rect 23848 22108 23900 22160
rect 26056 22108 26108 22160
rect 10232 22015 10284 22024
rect 10232 21981 10241 22015
rect 10241 21981 10275 22015
rect 10275 21981 10284 22015
rect 10232 21972 10284 21981
rect 10600 21972 10652 22024
rect 8668 21904 8720 21956
rect 10968 21947 11020 21956
rect 10968 21913 10977 21947
rect 10977 21913 11011 21947
rect 11011 21913 11020 21947
rect 10968 21904 11020 21913
rect 12072 21972 12124 22024
rect 12808 21972 12860 22024
rect 12532 21904 12584 21956
rect 13912 21972 13964 22024
rect 14096 21972 14148 22024
rect 15108 22040 15160 22092
rect 15292 22040 15344 22092
rect 15844 22083 15896 22092
rect 15844 22049 15853 22083
rect 15853 22049 15887 22083
rect 15887 22049 15896 22083
rect 15844 22040 15896 22049
rect 16488 22040 16540 22092
rect 17868 22040 17920 22092
rect 20904 22040 20956 22092
rect 22008 22040 22060 22092
rect 23388 22040 23440 22092
rect 14372 22015 14424 22024
rect 14372 21981 14381 22015
rect 14381 21981 14415 22015
rect 14415 21981 14424 22015
rect 14372 21972 14424 21981
rect 14740 21972 14792 22024
rect 16304 21972 16356 22024
rect 17960 21972 18012 22024
rect 18236 21972 18288 22024
rect 19892 22015 19944 22024
rect 3240 21836 3292 21888
rect 3516 21836 3568 21888
rect 5080 21836 5132 21888
rect 6644 21879 6696 21888
rect 6644 21845 6653 21879
rect 6653 21845 6687 21879
rect 6687 21845 6696 21879
rect 6644 21836 6696 21845
rect 6828 21836 6880 21888
rect 8484 21836 8536 21888
rect 11796 21836 11848 21888
rect 12440 21836 12492 21888
rect 12624 21836 12676 21888
rect 13084 21836 13136 21888
rect 14096 21836 14148 21888
rect 14832 21904 14884 21956
rect 16856 21904 16908 21956
rect 19892 21981 19901 22015
rect 19901 21981 19935 22015
rect 19935 21981 19944 22015
rect 19892 21972 19944 21981
rect 21640 22015 21692 22024
rect 21640 21981 21649 22015
rect 21649 21981 21683 22015
rect 21683 21981 21692 22015
rect 21640 21972 21692 21981
rect 23572 21972 23624 22024
rect 26792 22040 26844 22092
rect 25872 22015 25924 22024
rect 25872 21981 25881 22015
rect 25881 21981 25915 22015
rect 25915 21981 25924 22015
rect 25872 21972 25924 21981
rect 26056 22015 26108 22024
rect 26056 21981 26065 22015
rect 26065 21981 26099 22015
rect 26099 21981 26108 22015
rect 26056 21972 26108 21981
rect 16120 21836 16172 21888
rect 19616 21904 19668 21956
rect 20904 21904 20956 21956
rect 24676 21904 24728 21956
rect 18052 21836 18104 21888
rect 21824 21836 21876 21888
rect 23112 21879 23164 21888
rect 23112 21845 23121 21879
rect 23121 21845 23155 21879
rect 23155 21845 23164 21879
rect 23112 21836 23164 21845
rect 23664 21836 23716 21888
rect 24032 21836 24084 21888
rect 24768 21836 24820 21888
rect 25044 21904 25096 21956
rect 25504 21904 25556 21956
rect 26240 21904 26292 21956
rect 26792 21904 26844 21956
rect 25596 21836 25648 21888
rect 25688 21836 25740 21888
rect 9935 21734 9987 21786
rect 9999 21734 10051 21786
rect 10063 21734 10115 21786
rect 10127 21734 10179 21786
rect 10191 21734 10243 21786
rect 18920 21734 18972 21786
rect 18984 21734 19036 21786
rect 19048 21734 19100 21786
rect 19112 21734 19164 21786
rect 19176 21734 19228 21786
rect 2872 21632 2924 21684
rect 3240 21632 3292 21684
rect 4068 21675 4120 21684
rect 3148 21564 3200 21616
rect 4068 21641 4077 21675
rect 4077 21641 4111 21675
rect 4111 21641 4120 21675
rect 4068 21632 4120 21641
rect 4160 21632 4212 21684
rect 4896 21632 4948 21684
rect 7380 21632 7432 21684
rect 7656 21675 7708 21684
rect 7656 21641 7665 21675
rect 7665 21641 7699 21675
rect 7699 21641 7708 21675
rect 7656 21632 7708 21641
rect 3608 21496 3660 21548
rect 4252 21496 4304 21548
rect 4528 21496 4580 21548
rect 3240 21360 3292 21412
rect 2596 21292 2648 21344
rect 4160 21428 4212 21480
rect 4988 21564 5040 21616
rect 6644 21564 6696 21616
rect 4804 21496 4856 21548
rect 5080 21539 5132 21548
rect 5080 21505 5089 21539
rect 5089 21505 5123 21539
rect 5123 21505 5132 21539
rect 5080 21496 5132 21505
rect 5540 21496 5592 21548
rect 6644 21428 6696 21480
rect 6828 21539 6880 21548
rect 6828 21505 6837 21539
rect 6837 21505 6871 21539
rect 6871 21505 6880 21539
rect 7012 21539 7064 21548
rect 6828 21496 6880 21505
rect 7012 21505 7021 21539
rect 7021 21505 7055 21539
rect 7055 21505 7064 21539
rect 7012 21496 7064 21505
rect 7472 21564 7524 21616
rect 10416 21632 10468 21684
rect 10600 21632 10652 21684
rect 7196 21496 7248 21548
rect 7748 21496 7800 21548
rect 7840 21496 7892 21548
rect 8116 21539 8168 21548
rect 8116 21505 8125 21539
rect 8125 21505 8159 21539
rect 8159 21505 8168 21539
rect 8116 21496 8168 21505
rect 8576 21564 8628 21616
rect 8944 21564 8996 21616
rect 6920 21428 6972 21480
rect 7472 21428 7524 21480
rect 8484 21496 8536 21548
rect 9404 21539 9456 21548
rect 9404 21505 9413 21539
rect 9413 21505 9447 21539
rect 9447 21505 9456 21539
rect 9404 21496 9456 21505
rect 9588 21564 9640 21616
rect 11336 21632 11388 21684
rect 12164 21632 12216 21684
rect 13452 21632 13504 21684
rect 9864 21496 9916 21548
rect 10600 21539 10652 21548
rect 10600 21505 10609 21539
rect 10609 21505 10643 21539
rect 10643 21505 10652 21539
rect 10600 21496 10652 21505
rect 9588 21471 9640 21480
rect 9588 21437 9605 21471
rect 9605 21437 9640 21471
rect 9588 21428 9640 21437
rect 9680 21428 9732 21480
rect 11520 21428 11572 21480
rect 12348 21564 12400 21616
rect 13820 21496 13872 21548
rect 14832 21496 14884 21548
rect 18788 21564 18840 21616
rect 16120 21539 16172 21548
rect 16120 21505 16129 21539
rect 16129 21505 16163 21539
rect 16163 21505 16172 21539
rect 16120 21496 16172 21505
rect 17960 21539 18012 21548
rect 17960 21505 17969 21539
rect 17969 21505 18003 21539
rect 18003 21505 18012 21539
rect 17960 21496 18012 21505
rect 18052 21496 18104 21548
rect 19892 21632 19944 21684
rect 20628 21632 20680 21684
rect 23388 21632 23440 21684
rect 23664 21632 23716 21684
rect 24768 21632 24820 21684
rect 25688 21675 25740 21684
rect 20812 21607 20864 21616
rect 20812 21573 20821 21607
rect 20821 21573 20855 21607
rect 20855 21573 20864 21607
rect 22008 21607 22060 21616
rect 20812 21564 20864 21573
rect 22008 21573 22017 21607
rect 22017 21573 22051 21607
rect 22051 21573 22060 21607
rect 22008 21564 22060 21573
rect 8668 21360 8720 21412
rect 4896 21292 4948 21344
rect 4988 21292 5040 21344
rect 7196 21292 7248 21344
rect 7380 21292 7432 21344
rect 9680 21292 9732 21344
rect 10692 21360 10744 21412
rect 9864 21292 9916 21344
rect 10876 21292 10928 21344
rect 11336 21292 11388 21344
rect 11520 21292 11572 21344
rect 12256 21428 12308 21480
rect 17868 21471 17920 21480
rect 17868 21437 17877 21471
rect 17877 21437 17911 21471
rect 17911 21437 17920 21471
rect 17868 21428 17920 21437
rect 19616 21471 19668 21480
rect 19616 21437 19625 21471
rect 19625 21437 19659 21471
rect 19659 21437 19668 21471
rect 21824 21496 21876 21548
rect 22100 21496 22152 21548
rect 22652 21564 22704 21616
rect 23112 21564 23164 21616
rect 22560 21496 22612 21548
rect 23388 21496 23440 21548
rect 24584 21564 24636 21616
rect 24860 21564 24912 21616
rect 25688 21641 25697 21675
rect 25697 21641 25731 21675
rect 25731 21641 25740 21675
rect 25688 21632 25740 21641
rect 25964 21632 26016 21684
rect 25596 21564 25648 21616
rect 26148 21564 26200 21616
rect 19616 21428 19668 21437
rect 19892 21428 19944 21480
rect 20536 21428 20588 21480
rect 23572 21428 23624 21480
rect 14280 21292 14332 21344
rect 15016 21292 15068 21344
rect 17224 21335 17276 21344
rect 17224 21301 17233 21335
rect 17233 21301 17267 21335
rect 17267 21301 17276 21335
rect 17224 21292 17276 21301
rect 18972 21335 19024 21344
rect 18972 21301 18981 21335
rect 18981 21301 19015 21335
rect 19015 21301 19024 21335
rect 18972 21292 19024 21301
rect 23204 21360 23256 21412
rect 24768 21496 24820 21548
rect 25044 21496 25096 21548
rect 26056 21496 26108 21548
rect 26240 21539 26292 21548
rect 26240 21505 26249 21539
rect 26249 21505 26283 21539
rect 26283 21505 26292 21539
rect 26240 21496 26292 21505
rect 26976 21539 27028 21548
rect 26976 21505 26985 21539
rect 26985 21505 27019 21539
rect 27019 21505 27028 21539
rect 26976 21496 27028 21505
rect 26608 21428 26660 21480
rect 24676 21360 24728 21412
rect 19432 21292 19484 21344
rect 20628 21292 20680 21344
rect 20904 21335 20956 21344
rect 20904 21301 20913 21335
rect 20913 21301 20947 21335
rect 20947 21301 20956 21335
rect 20904 21292 20956 21301
rect 21640 21292 21692 21344
rect 23848 21335 23900 21344
rect 23848 21301 23857 21335
rect 23857 21301 23891 21335
rect 23891 21301 23900 21335
rect 23848 21292 23900 21301
rect 25688 21292 25740 21344
rect 5442 21190 5494 21242
rect 5506 21190 5558 21242
rect 5570 21190 5622 21242
rect 5634 21190 5686 21242
rect 5698 21190 5750 21242
rect 14428 21190 14480 21242
rect 14492 21190 14544 21242
rect 14556 21190 14608 21242
rect 14620 21190 14672 21242
rect 14684 21190 14736 21242
rect 23413 21190 23465 21242
rect 23477 21190 23529 21242
rect 23541 21190 23593 21242
rect 23605 21190 23657 21242
rect 23669 21190 23721 21242
rect 4988 21088 5040 21140
rect 6644 21088 6696 21140
rect 7656 21131 7708 21140
rect 7656 21097 7665 21131
rect 7665 21097 7699 21131
rect 7699 21097 7708 21131
rect 7656 21088 7708 21097
rect 8392 21088 8444 21140
rect 10692 21131 10744 21140
rect 10692 21097 10701 21131
rect 10701 21097 10735 21131
rect 10735 21097 10744 21131
rect 10692 21088 10744 21097
rect 14004 21088 14056 21140
rect 16856 21131 16908 21140
rect 1216 21020 1268 21072
rect 2228 20884 2280 20936
rect 3976 21020 4028 21072
rect 3148 20884 3200 20936
rect 4160 20952 4212 21004
rect 3792 20884 3844 20936
rect 6184 20952 6236 21004
rect 4804 20884 4856 20936
rect 10140 21063 10192 21072
rect 10140 21029 10149 21063
rect 10149 21029 10183 21063
rect 10183 21029 10192 21063
rect 10140 21020 10192 21029
rect 10324 21020 10376 21072
rect 2872 20816 2924 20868
rect 2320 20748 2372 20800
rect 2412 20748 2464 20800
rect 4712 20816 4764 20868
rect 3240 20791 3292 20800
rect 3240 20757 3249 20791
rect 3249 20757 3283 20791
rect 3283 20757 3292 20791
rect 3240 20748 3292 20757
rect 3608 20748 3660 20800
rect 3792 20791 3844 20800
rect 3792 20757 3801 20791
rect 3801 20757 3835 20791
rect 3835 20757 3844 20791
rect 3792 20748 3844 20757
rect 5356 20791 5408 20800
rect 5356 20757 5365 20791
rect 5365 20757 5399 20791
rect 5399 20757 5408 20791
rect 5356 20748 5408 20757
rect 5448 20748 5500 20800
rect 7288 20952 7340 21004
rect 7472 20927 7524 20936
rect 7472 20893 7481 20927
rect 7481 20893 7515 20927
rect 7515 20893 7524 20927
rect 7472 20884 7524 20893
rect 7932 20884 7984 20936
rect 8944 20927 8996 20936
rect 8944 20893 8953 20927
rect 8953 20893 8987 20927
rect 8987 20893 8996 20927
rect 8944 20884 8996 20893
rect 9588 20927 9640 20936
rect 8024 20816 8076 20868
rect 9588 20893 9597 20927
rect 9597 20893 9631 20927
rect 9631 20893 9640 20927
rect 9588 20884 9640 20893
rect 9680 20884 9732 20936
rect 9956 20927 10008 20936
rect 9956 20893 9965 20927
rect 9965 20893 9999 20927
rect 9999 20893 10008 20927
rect 9956 20884 10008 20893
rect 10600 20927 10652 20936
rect 10600 20893 10609 20927
rect 10609 20893 10643 20927
rect 10643 20893 10652 20927
rect 10600 20884 10652 20893
rect 10876 20884 10928 20936
rect 11336 20884 11388 20936
rect 11796 20884 11848 20936
rect 6736 20748 6788 20800
rect 7196 20748 7248 20800
rect 7564 20748 7616 20800
rect 9036 20748 9088 20800
rect 9680 20748 9732 20800
rect 11520 20791 11572 20800
rect 11520 20757 11529 20791
rect 11529 20757 11563 20791
rect 11563 20757 11572 20791
rect 11520 20748 11572 20757
rect 11888 20816 11940 20868
rect 13084 20884 13136 20936
rect 16856 21097 16865 21131
rect 16865 21097 16899 21131
rect 16899 21097 16908 21131
rect 16856 21088 16908 21097
rect 18972 21088 19024 21140
rect 20812 21088 20864 21140
rect 21088 21088 21140 21140
rect 22376 21131 22428 21140
rect 22376 21097 22385 21131
rect 22385 21097 22419 21131
rect 22419 21097 22428 21131
rect 22376 21088 22428 21097
rect 23756 21131 23808 21140
rect 23756 21097 23765 21131
rect 23765 21097 23799 21131
rect 23799 21097 23808 21131
rect 23756 21088 23808 21097
rect 24400 21088 24452 21140
rect 18328 21020 18380 21072
rect 19892 21020 19944 21072
rect 23112 21020 23164 21072
rect 16304 20884 16356 20936
rect 16764 20884 16816 20936
rect 17224 20884 17276 20936
rect 18052 20884 18104 20936
rect 13820 20816 13872 20868
rect 15200 20816 15252 20868
rect 19616 20884 19668 20936
rect 19432 20816 19484 20868
rect 20352 20884 20404 20936
rect 20536 20884 20588 20936
rect 21916 20952 21968 21004
rect 21088 20927 21140 20936
rect 21088 20893 21097 20927
rect 21097 20893 21131 20927
rect 21131 20893 21140 20927
rect 21088 20884 21140 20893
rect 21180 20927 21232 20936
rect 21180 20893 21189 20927
rect 21189 20893 21223 20927
rect 21223 20893 21232 20927
rect 21824 20927 21876 20936
rect 21180 20884 21232 20893
rect 21824 20893 21833 20927
rect 21833 20893 21867 20927
rect 21867 20893 21876 20927
rect 21824 20884 21876 20893
rect 22008 20884 22060 20936
rect 20996 20816 21048 20868
rect 23296 20952 23348 21004
rect 23756 20952 23808 21004
rect 24124 20952 24176 21004
rect 24400 20952 24452 21004
rect 24952 20952 25004 21004
rect 25964 20995 26016 21004
rect 25964 20961 25973 20995
rect 25973 20961 26007 20995
rect 26007 20961 26016 20995
rect 25964 20952 26016 20961
rect 22560 20927 22612 20936
rect 22560 20893 22569 20927
rect 22569 20893 22603 20927
rect 22603 20893 22612 20927
rect 22560 20884 22612 20893
rect 23848 20884 23900 20936
rect 25780 20884 25832 20936
rect 25320 20816 25372 20868
rect 12164 20748 12216 20800
rect 13544 20748 13596 20800
rect 17592 20748 17644 20800
rect 17868 20791 17920 20800
rect 17868 20757 17877 20791
rect 17877 20757 17911 20791
rect 17911 20757 17920 20791
rect 17868 20748 17920 20757
rect 20352 20748 20404 20800
rect 21364 20748 21416 20800
rect 21640 20791 21692 20800
rect 21640 20757 21649 20791
rect 21649 20757 21683 20791
rect 21683 20757 21692 20791
rect 21640 20748 21692 20757
rect 22008 20748 22060 20800
rect 24216 20748 24268 20800
rect 25044 20748 25096 20800
rect 25596 20748 25648 20800
rect 26148 20748 26200 20800
rect 9935 20646 9987 20698
rect 9999 20646 10051 20698
rect 10063 20646 10115 20698
rect 10127 20646 10179 20698
rect 10191 20646 10243 20698
rect 18920 20646 18972 20698
rect 18984 20646 19036 20698
rect 19048 20646 19100 20698
rect 19112 20646 19164 20698
rect 19176 20646 19228 20698
rect 6920 20587 6972 20596
rect 2688 20408 2740 20460
rect 4896 20451 4948 20460
rect 1492 20340 1544 20392
rect 1676 20340 1728 20392
rect 2228 20340 2280 20392
rect 4896 20417 4905 20451
rect 4905 20417 4939 20451
rect 4939 20417 4948 20451
rect 4896 20408 4948 20417
rect 5448 20476 5500 20528
rect 6092 20408 6144 20460
rect 6184 20340 6236 20392
rect 6920 20553 6929 20587
rect 6929 20553 6963 20587
rect 6963 20553 6972 20587
rect 6920 20544 6972 20553
rect 8852 20544 8904 20596
rect 8024 20476 8076 20528
rect 9036 20476 9088 20528
rect 9588 20476 9640 20528
rect 10600 20476 10652 20528
rect 11244 20476 11296 20528
rect 6736 20451 6788 20460
rect 6736 20417 6745 20451
rect 6745 20417 6779 20451
rect 6779 20417 6788 20451
rect 6736 20408 6788 20417
rect 7564 20408 7616 20460
rect 7656 20451 7708 20460
rect 7656 20417 7665 20451
rect 7665 20417 7699 20451
rect 7699 20417 7708 20451
rect 7656 20408 7708 20417
rect 7840 20408 7892 20460
rect 9220 20408 9272 20460
rect 9772 20451 9824 20460
rect 9772 20417 9781 20451
rect 9781 20417 9815 20451
rect 9815 20417 9824 20451
rect 9772 20408 9824 20417
rect 10600 20340 10652 20392
rect 4528 20272 4580 20324
rect 1492 20204 1544 20256
rect 2872 20204 2924 20256
rect 4068 20204 4120 20256
rect 7472 20272 7524 20324
rect 6644 20247 6696 20256
rect 6644 20213 6653 20247
rect 6653 20213 6687 20247
rect 6687 20213 6696 20247
rect 6644 20204 6696 20213
rect 7012 20204 7064 20256
rect 8852 20272 8904 20324
rect 11796 20408 11848 20460
rect 11888 20383 11940 20392
rect 11888 20349 11897 20383
rect 11897 20349 11931 20383
rect 11931 20349 11940 20383
rect 11888 20340 11940 20349
rect 11152 20272 11204 20324
rect 12348 20451 12400 20460
rect 12348 20417 12362 20451
rect 12362 20417 12396 20451
rect 12396 20417 12400 20451
rect 12348 20408 12400 20417
rect 12900 20544 12952 20596
rect 16948 20544 17000 20596
rect 17408 20544 17460 20596
rect 19708 20544 19760 20596
rect 13084 20519 13136 20528
rect 13084 20485 13093 20519
rect 13093 20485 13127 20519
rect 13127 20485 13136 20519
rect 13084 20476 13136 20485
rect 14004 20476 14056 20528
rect 12808 20340 12860 20392
rect 13820 20408 13872 20460
rect 15660 20476 15712 20528
rect 14188 20451 14240 20460
rect 14188 20417 14222 20451
rect 14222 20417 14240 20451
rect 14188 20408 14240 20417
rect 15292 20408 15344 20460
rect 16764 20408 16816 20460
rect 17040 20451 17092 20460
rect 17040 20417 17049 20451
rect 17049 20417 17083 20451
rect 17083 20417 17092 20451
rect 17040 20408 17092 20417
rect 17868 20476 17920 20528
rect 17960 20476 18012 20528
rect 18604 20476 18656 20528
rect 20996 20544 21048 20596
rect 21364 20544 21416 20596
rect 24032 20587 24084 20596
rect 18052 20451 18104 20460
rect 18052 20417 18086 20451
rect 18086 20417 18104 20451
rect 15844 20340 15896 20392
rect 12624 20272 12676 20324
rect 13544 20272 13596 20324
rect 9312 20204 9364 20256
rect 12072 20204 12124 20256
rect 13820 20204 13872 20256
rect 15108 20204 15160 20256
rect 16028 20272 16080 20324
rect 16396 20340 16448 20392
rect 18052 20408 18104 20417
rect 19524 20408 19576 20460
rect 19892 20451 19944 20460
rect 19892 20417 19901 20451
rect 19901 20417 19935 20451
rect 19935 20417 19944 20451
rect 19892 20408 19944 20417
rect 20628 20408 20680 20460
rect 21824 20408 21876 20460
rect 21916 20408 21968 20460
rect 24032 20553 24041 20587
rect 24041 20553 24075 20587
rect 24075 20553 24084 20587
rect 24032 20544 24084 20553
rect 27344 20587 27396 20596
rect 27344 20553 27353 20587
rect 27353 20553 27387 20587
rect 27387 20553 27396 20587
rect 27344 20544 27396 20553
rect 22192 20408 22244 20460
rect 22376 20451 22428 20460
rect 22376 20417 22385 20451
rect 22385 20417 22419 20451
rect 22419 20417 22428 20451
rect 22376 20408 22428 20417
rect 17224 20340 17276 20392
rect 24860 20476 24912 20528
rect 25044 20476 25096 20528
rect 23848 20408 23900 20460
rect 24952 20408 25004 20460
rect 25596 20451 25648 20460
rect 25596 20417 25605 20451
rect 25605 20417 25639 20451
rect 25639 20417 25648 20451
rect 25596 20408 25648 20417
rect 25780 20408 25832 20460
rect 15476 20204 15528 20256
rect 16580 20204 16632 20256
rect 19156 20247 19208 20256
rect 19156 20213 19165 20247
rect 19165 20213 19199 20247
rect 19199 20213 19208 20247
rect 19156 20204 19208 20213
rect 19432 20204 19484 20256
rect 24216 20383 24268 20392
rect 24216 20349 24225 20383
rect 24225 20349 24259 20383
rect 24259 20349 24268 20383
rect 24216 20340 24268 20349
rect 24952 20272 25004 20324
rect 26332 20340 26384 20392
rect 21364 20204 21416 20256
rect 24124 20204 24176 20256
rect 5442 20102 5494 20154
rect 5506 20102 5558 20154
rect 5570 20102 5622 20154
rect 5634 20102 5686 20154
rect 5698 20102 5750 20154
rect 14428 20102 14480 20154
rect 14492 20102 14544 20154
rect 14556 20102 14608 20154
rect 14620 20102 14672 20154
rect 14684 20102 14736 20154
rect 23413 20102 23465 20154
rect 23477 20102 23529 20154
rect 23541 20102 23593 20154
rect 23605 20102 23657 20154
rect 23669 20102 23721 20154
rect 1860 20000 1912 20052
rect 3608 20000 3660 20052
rect 4068 20000 4120 20052
rect 5264 20043 5316 20052
rect 2412 19932 2464 19984
rect 4436 19975 4488 19984
rect 4436 19941 4445 19975
rect 4445 19941 4479 19975
rect 4479 19941 4488 19975
rect 4436 19932 4488 19941
rect 5264 20009 5273 20043
rect 5273 20009 5307 20043
rect 5307 20009 5316 20043
rect 5264 20000 5316 20009
rect 7656 20000 7708 20052
rect 8116 20000 8168 20052
rect 11520 20000 11572 20052
rect 8484 19932 8536 19984
rect 4068 19864 4120 19916
rect 6184 19864 6236 19916
rect 6828 19864 6880 19916
rect 7656 19864 7708 19916
rect 8576 19864 8628 19916
rect 8944 19864 8996 19916
rect 4252 19771 4304 19780
rect 4252 19737 4261 19771
rect 4261 19737 4295 19771
rect 4295 19737 4304 19771
rect 4252 19728 4304 19737
rect 1124 19660 1176 19712
rect 3056 19703 3108 19712
rect 3056 19669 3065 19703
rect 3065 19669 3099 19703
rect 3099 19669 3108 19703
rect 3056 19660 3108 19669
rect 3608 19660 3660 19712
rect 5264 19796 5316 19848
rect 6092 19839 6144 19848
rect 4896 19728 4948 19780
rect 6092 19805 6101 19839
rect 6101 19805 6135 19839
rect 6135 19805 6144 19839
rect 6092 19796 6144 19805
rect 6644 19796 6696 19848
rect 13452 20000 13504 20052
rect 14004 20000 14056 20052
rect 15200 20043 15252 20052
rect 15200 20009 15209 20043
rect 15209 20009 15243 20043
rect 15243 20009 15252 20043
rect 15200 20000 15252 20009
rect 6920 19728 6972 19780
rect 7380 19728 7432 19780
rect 9036 19728 9088 19780
rect 7472 19660 7524 19712
rect 8392 19660 8444 19712
rect 9496 19796 9548 19848
rect 9588 19839 9640 19848
rect 9588 19805 9597 19839
rect 9597 19805 9631 19839
rect 9631 19805 9640 19839
rect 10324 19839 10376 19848
rect 9588 19796 9640 19805
rect 10324 19805 10333 19839
rect 10333 19805 10367 19839
rect 10367 19805 10376 19839
rect 10324 19796 10376 19805
rect 9864 19728 9916 19780
rect 12072 19796 12124 19848
rect 14280 19932 14332 19984
rect 12808 19864 12860 19916
rect 14372 19907 14424 19916
rect 13268 19796 13320 19848
rect 14372 19873 14381 19907
rect 14381 19873 14415 19907
rect 14415 19873 14424 19907
rect 14372 19864 14424 19873
rect 17040 20000 17092 20052
rect 18052 20000 18104 20052
rect 18696 20000 18748 20052
rect 19340 20000 19392 20052
rect 21088 20000 21140 20052
rect 21364 20043 21416 20052
rect 21364 20009 21373 20043
rect 21373 20009 21407 20043
rect 21407 20009 21416 20043
rect 21364 20000 21416 20009
rect 22376 20000 22428 20052
rect 24308 20000 24360 20052
rect 15660 19932 15712 19984
rect 14280 19839 14332 19848
rect 10876 19728 10928 19780
rect 12256 19660 12308 19712
rect 12900 19660 12952 19712
rect 13728 19728 13780 19780
rect 14280 19805 14289 19839
rect 14289 19805 14323 19839
rect 14323 19805 14332 19839
rect 14280 19796 14332 19805
rect 14464 19839 14516 19848
rect 14464 19805 14473 19839
rect 14473 19805 14507 19839
rect 14507 19805 14516 19839
rect 14464 19796 14516 19805
rect 15016 19796 15068 19848
rect 15660 19839 15712 19848
rect 15660 19805 15669 19839
rect 15669 19805 15703 19839
rect 15703 19805 15712 19839
rect 18052 19864 18104 19916
rect 19708 19864 19760 19916
rect 15660 19796 15712 19805
rect 16304 19839 16356 19848
rect 16304 19805 16313 19839
rect 16313 19805 16347 19839
rect 16347 19805 16356 19839
rect 16304 19796 16356 19805
rect 16580 19839 16632 19848
rect 16580 19805 16614 19839
rect 16614 19805 16632 19839
rect 16580 19796 16632 19805
rect 17040 19796 17092 19848
rect 18328 19839 18380 19848
rect 16488 19728 16540 19780
rect 14648 19660 14700 19712
rect 15108 19660 15160 19712
rect 15292 19660 15344 19712
rect 15844 19660 15896 19712
rect 16580 19660 16632 19712
rect 16764 19660 16816 19712
rect 17684 19703 17736 19712
rect 17684 19669 17693 19703
rect 17693 19669 17727 19703
rect 17727 19669 17736 19703
rect 17684 19660 17736 19669
rect 18328 19805 18337 19839
rect 18337 19805 18371 19839
rect 18371 19805 18380 19839
rect 18328 19796 18380 19805
rect 19156 19796 19208 19848
rect 19432 19839 19484 19848
rect 19432 19805 19441 19839
rect 19441 19805 19475 19839
rect 19475 19805 19484 19839
rect 19432 19796 19484 19805
rect 19984 19796 20036 19848
rect 22560 19932 22612 19984
rect 26332 20000 26384 20052
rect 22100 19864 22152 19916
rect 20352 19839 20404 19848
rect 20352 19805 20361 19839
rect 20361 19805 20395 19839
rect 20395 19805 20404 19839
rect 20352 19796 20404 19805
rect 22284 19796 22336 19848
rect 23112 19864 23164 19916
rect 23572 19864 23624 19916
rect 24768 19864 24820 19916
rect 25228 19864 25280 19916
rect 25964 19907 26016 19916
rect 25964 19873 25973 19907
rect 25973 19873 26007 19907
rect 26007 19873 26016 19907
rect 25964 19864 26016 19873
rect 22652 19839 22704 19848
rect 22652 19805 22661 19839
rect 22661 19805 22695 19839
rect 22695 19805 22704 19839
rect 22652 19796 22704 19805
rect 22192 19728 22244 19780
rect 24216 19796 24268 19848
rect 24308 19796 24360 19848
rect 24492 19796 24544 19848
rect 27252 19796 27304 19848
rect 25872 19728 25924 19780
rect 19800 19660 19852 19712
rect 20628 19660 20680 19712
rect 23296 19660 23348 19712
rect 24768 19703 24820 19712
rect 24768 19669 24777 19703
rect 24777 19669 24811 19703
rect 24811 19669 24820 19703
rect 24768 19660 24820 19669
rect 25044 19660 25096 19712
rect 25228 19703 25280 19712
rect 25228 19669 25237 19703
rect 25237 19669 25271 19703
rect 25271 19669 25280 19703
rect 25228 19660 25280 19669
rect 25596 19660 25648 19712
rect 9935 19558 9987 19610
rect 9999 19558 10051 19610
rect 10063 19558 10115 19610
rect 10127 19558 10179 19610
rect 10191 19558 10243 19610
rect 18920 19558 18972 19610
rect 18984 19558 19036 19610
rect 19048 19558 19100 19610
rect 19112 19558 19164 19610
rect 19176 19558 19228 19610
rect 1860 19456 1912 19508
rect 3608 19456 3660 19508
rect 4436 19456 4488 19508
rect 4896 19456 4948 19508
rect 6092 19456 6144 19508
rect 7288 19456 7340 19508
rect 8300 19456 8352 19508
rect 13268 19456 13320 19508
rect 13452 19456 13504 19508
rect 14004 19456 14056 19508
rect 14464 19456 14516 19508
rect 15936 19456 15988 19508
rect 17684 19456 17736 19508
rect 18328 19456 18380 19508
rect 2504 19363 2556 19372
rect 2504 19329 2513 19363
rect 2513 19329 2547 19363
rect 2547 19329 2556 19363
rect 2504 19320 2556 19329
rect 3148 19363 3200 19372
rect 3148 19329 3157 19363
rect 3157 19329 3191 19363
rect 3191 19329 3200 19363
rect 3148 19320 3200 19329
rect 3608 19363 3660 19372
rect 3608 19329 3617 19363
rect 3617 19329 3651 19363
rect 3651 19329 3660 19363
rect 3608 19320 3660 19329
rect 6092 19320 6144 19372
rect 2688 19184 2740 19236
rect 5264 19184 5316 19236
rect 7564 19252 7616 19304
rect 7288 19184 7340 19236
rect 2596 19116 2648 19168
rect 4620 19116 4672 19168
rect 6920 19116 6972 19168
rect 7012 19116 7064 19168
rect 7840 19320 7892 19372
rect 8116 19363 8168 19372
rect 8116 19329 8125 19363
rect 8125 19329 8159 19363
rect 8159 19329 8168 19363
rect 8116 19320 8168 19329
rect 9036 19363 9088 19372
rect 9036 19329 9070 19363
rect 9070 19329 9088 19363
rect 9036 19320 9088 19329
rect 9588 19388 9640 19440
rect 10232 19320 10284 19372
rect 8392 19252 8444 19304
rect 10692 19431 10744 19440
rect 10692 19397 10701 19431
rect 10701 19397 10735 19431
rect 10735 19397 10744 19431
rect 10692 19388 10744 19397
rect 10968 19388 11020 19440
rect 11612 19320 11664 19372
rect 11888 19363 11940 19372
rect 11888 19329 11897 19363
rect 11897 19329 11931 19363
rect 11931 19329 11940 19363
rect 11888 19320 11940 19329
rect 12072 19320 12124 19372
rect 12992 19388 13044 19440
rect 12624 19363 12676 19372
rect 12624 19329 12633 19363
rect 12633 19329 12667 19363
rect 12667 19329 12676 19363
rect 12624 19320 12676 19329
rect 12808 19363 12860 19372
rect 12808 19329 12817 19363
rect 12817 19329 12851 19363
rect 12851 19329 12860 19363
rect 13820 19363 13872 19372
rect 12808 19320 12860 19329
rect 13820 19329 13843 19363
rect 13843 19329 13872 19363
rect 13820 19320 13872 19329
rect 14188 19363 14240 19372
rect 12440 19252 12492 19304
rect 14188 19329 14197 19363
rect 14197 19329 14231 19363
rect 14231 19329 14240 19363
rect 14188 19320 14240 19329
rect 16304 19388 16356 19440
rect 19616 19456 19668 19508
rect 20628 19456 20680 19508
rect 14832 19320 14884 19372
rect 15752 19294 15804 19346
rect 16120 19320 16172 19372
rect 16764 19320 16816 19372
rect 17408 19363 17460 19372
rect 17408 19329 17417 19363
rect 17417 19329 17451 19363
rect 17451 19329 17460 19363
rect 17408 19320 17460 19329
rect 17868 19320 17920 19372
rect 18696 19320 18748 19372
rect 18880 19363 18932 19372
rect 18880 19329 18889 19363
rect 18889 19329 18923 19363
rect 18923 19329 18932 19363
rect 18880 19320 18932 19329
rect 16488 19252 16540 19304
rect 17224 19252 17276 19304
rect 18328 19252 18380 19304
rect 8576 19184 8628 19236
rect 8116 19116 8168 19168
rect 9956 19116 10008 19168
rect 10324 19184 10376 19236
rect 10232 19116 10284 19168
rect 10784 19159 10836 19168
rect 10784 19125 10793 19159
rect 10793 19125 10827 19159
rect 10827 19125 10836 19159
rect 10784 19116 10836 19125
rect 11520 19159 11572 19168
rect 11520 19125 11529 19159
rect 11529 19125 11563 19159
rect 11563 19125 11572 19159
rect 11520 19116 11572 19125
rect 11888 19116 11940 19168
rect 12532 19184 12584 19236
rect 13728 19184 13780 19236
rect 12440 19116 12492 19168
rect 13084 19116 13136 19168
rect 13360 19116 13412 19168
rect 14464 19184 14516 19236
rect 17868 19184 17920 19236
rect 19064 19184 19116 19236
rect 14096 19116 14148 19168
rect 16488 19116 16540 19168
rect 18328 19116 18380 19168
rect 20076 19320 20128 19372
rect 22376 19456 22428 19508
rect 23020 19456 23072 19508
rect 22192 19388 22244 19440
rect 23204 19388 23256 19440
rect 22652 19320 22704 19372
rect 23296 19320 23348 19372
rect 23848 19320 23900 19372
rect 24124 19431 24176 19440
rect 24124 19397 24133 19431
rect 24133 19397 24167 19431
rect 24167 19397 24176 19431
rect 24124 19388 24176 19397
rect 24492 19388 24544 19440
rect 24768 19388 24820 19440
rect 26424 19456 26476 19508
rect 26884 19456 26936 19508
rect 23664 19252 23716 19304
rect 22652 19184 22704 19236
rect 23112 19184 23164 19236
rect 23572 19184 23624 19236
rect 23848 19184 23900 19236
rect 25780 19320 25832 19372
rect 26056 19320 26108 19372
rect 25320 19252 25372 19304
rect 26332 19252 26384 19304
rect 19616 19159 19668 19168
rect 19616 19125 19625 19159
rect 19625 19125 19659 19159
rect 19659 19125 19668 19159
rect 19616 19116 19668 19125
rect 20076 19116 20128 19168
rect 22284 19116 22336 19168
rect 24032 19116 24084 19168
rect 24216 19116 24268 19168
rect 24952 19116 25004 19168
rect 25044 19116 25096 19168
rect 25320 19116 25372 19168
rect 5442 19014 5494 19066
rect 5506 19014 5558 19066
rect 5570 19014 5622 19066
rect 5634 19014 5686 19066
rect 5698 19014 5750 19066
rect 14428 19014 14480 19066
rect 14492 19014 14544 19066
rect 14556 19014 14608 19066
rect 14620 19014 14672 19066
rect 14684 19014 14736 19066
rect 23413 19014 23465 19066
rect 23477 19014 23529 19066
rect 23541 19014 23593 19066
rect 23605 19014 23657 19066
rect 23669 19014 23721 19066
rect 3608 18912 3660 18964
rect 8484 18912 8536 18964
rect 9036 18912 9088 18964
rect 6828 18887 6880 18896
rect 3148 18776 3200 18828
rect 6828 18853 6837 18887
rect 6837 18853 6871 18887
rect 6871 18853 6880 18887
rect 6828 18844 6880 18853
rect 6920 18844 6972 18896
rect 11888 18912 11940 18964
rect 14004 18912 14056 18964
rect 14096 18912 14148 18964
rect 7564 18819 7616 18828
rect 1400 18708 1452 18760
rect 1860 18708 1912 18760
rect 2688 18708 2740 18760
rect 7564 18785 7573 18819
rect 7573 18785 7607 18819
rect 7607 18785 7616 18819
rect 7564 18776 7616 18785
rect 10692 18844 10744 18896
rect 10876 18887 10928 18896
rect 10876 18853 10885 18887
rect 10885 18853 10919 18887
rect 10919 18853 10928 18887
rect 10876 18844 10928 18853
rect 4896 18708 4948 18760
rect 5356 18708 5408 18760
rect 6552 18708 6604 18760
rect 1860 18572 1912 18624
rect 2228 18572 2280 18624
rect 3424 18572 3476 18624
rect 4436 18572 4488 18624
rect 5540 18640 5592 18692
rect 7012 18708 7064 18760
rect 7288 18751 7340 18760
rect 7288 18717 7297 18751
rect 7297 18717 7331 18751
rect 7331 18717 7340 18751
rect 7288 18708 7340 18717
rect 9956 18708 10008 18760
rect 6920 18640 6972 18692
rect 10692 18708 10744 18760
rect 12256 18844 12308 18896
rect 11612 18776 11664 18828
rect 14188 18844 14240 18896
rect 13084 18776 13136 18828
rect 14004 18776 14056 18828
rect 14280 18776 14332 18828
rect 16488 18912 16540 18964
rect 21916 18955 21968 18964
rect 16212 18844 16264 18896
rect 18328 18844 18380 18896
rect 18880 18844 18932 18896
rect 21916 18921 21925 18955
rect 21925 18921 21959 18955
rect 21959 18921 21968 18955
rect 21916 18912 21968 18921
rect 26792 18912 26844 18964
rect 27252 18955 27304 18964
rect 27252 18921 27261 18955
rect 27261 18921 27295 18955
rect 27295 18921 27304 18955
rect 27252 18912 27304 18921
rect 10600 18640 10652 18692
rect 10876 18640 10928 18692
rect 12072 18708 12124 18760
rect 12164 18751 12216 18760
rect 12164 18717 12173 18751
rect 12173 18717 12207 18751
rect 12207 18717 12216 18751
rect 12532 18751 12584 18760
rect 12164 18708 12216 18717
rect 12532 18717 12541 18751
rect 12541 18717 12575 18751
rect 12575 18717 12584 18751
rect 12532 18708 12584 18717
rect 11612 18640 11664 18692
rect 6092 18572 6144 18624
rect 6368 18572 6420 18624
rect 9496 18572 9548 18624
rect 12624 18572 12676 18624
rect 13820 18708 13872 18760
rect 14096 18751 14148 18760
rect 14096 18717 14105 18751
rect 14105 18717 14139 18751
rect 14139 18717 14148 18751
rect 14096 18708 14148 18717
rect 15016 18708 15068 18760
rect 15936 18708 15988 18760
rect 12992 18640 13044 18692
rect 15200 18572 15252 18624
rect 16488 18751 16540 18760
rect 16488 18717 16497 18751
rect 16497 18717 16531 18751
rect 16531 18717 16540 18751
rect 16488 18708 16540 18717
rect 22100 18776 22152 18828
rect 23204 18776 23256 18828
rect 17408 18708 17460 18760
rect 17776 18751 17828 18760
rect 17776 18717 17785 18751
rect 17785 18717 17819 18751
rect 17819 18717 17828 18751
rect 17776 18708 17828 18717
rect 17868 18708 17920 18760
rect 18420 18708 18472 18760
rect 18788 18708 18840 18760
rect 19515 18717 19547 18736
rect 19547 18717 19567 18736
rect 19515 18684 19567 18717
rect 17040 18572 17092 18624
rect 17224 18572 17276 18624
rect 22008 18708 22060 18760
rect 24308 18708 24360 18760
rect 24860 18708 24912 18760
rect 20904 18640 20956 18692
rect 25136 18640 25188 18692
rect 19892 18572 19944 18624
rect 21364 18572 21416 18624
rect 22284 18615 22336 18624
rect 22284 18581 22293 18615
rect 22293 18581 22327 18615
rect 22327 18581 22336 18615
rect 22284 18572 22336 18581
rect 22376 18615 22428 18624
rect 22376 18581 22385 18615
rect 22385 18581 22419 18615
rect 22419 18581 22428 18615
rect 23112 18615 23164 18624
rect 22376 18572 22428 18581
rect 23112 18581 23121 18615
rect 23121 18581 23155 18615
rect 23155 18581 23164 18615
rect 23112 18572 23164 18581
rect 24952 18572 25004 18624
rect 9935 18470 9987 18522
rect 9999 18470 10051 18522
rect 10063 18470 10115 18522
rect 10127 18470 10179 18522
rect 10191 18470 10243 18522
rect 18920 18470 18972 18522
rect 18984 18470 19036 18522
rect 19048 18470 19100 18522
rect 19112 18470 19164 18522
rect 19176 18470 19228 18522
rect 1952 18368 2004 18420
rect 2228 18368 2280 18420
rect 5356 18368 5408 18420
rect 3608 18300 3660 18352
rect 2504 18232 2556 18284
rect 1952 18207 2004 18216
rect 1952 18173 1961 18207
rect 1961 18173 1995 18207
rect 1995 18173 2004 18207
rect 1952 18164 2004 18173
rect 4160 18232 4212 18284
rect 4620 18232 4672 18284
rect 5356 18275 5408 18284
rect 5356 18241 5365 18275
rect 5365 18241 5399 18275
rect 5399 18241 5408 18275
rect 5356 18232 5408 18241
rect 5540 18343 5592 18352
rect 5540 18309 5549 18343
rect 5549 18309 5583 18343
rect 5583 18309 5592 18343
rect 5540 18300 5592 18309
rect 5908 18300 5960 18352
rect 6828 18300 6880 18352
rect 7288 18368 7340 18420
rect 5724 18232 5776 18284
rect 6460 18232 6512 18284
rect 4896 18164 4948 18216
rect 6368 18207 6420 18216
rect 6368 18173 6377 18207
rect 6377 18173 6411 18207
rect 6411 18173 6420 18207
rect 6368 18164 6420 18173
rect 5908 18096 5960 18148
rect 7932 18368 7984 18420
rect 10324 18368 10376 18420
rect 10876 18368 10928 18420
rect 12072 18343 12124 18352
rect 9496 18275 9548 18284
rect 9496 18241 9505 18275
rect 9505 18241 9539 18275
rect 9539 18241 9548 18275
rect 9496 18232 9548 18241
rect 9588 18232 9640 18284
rect 10140 18232 10192 18284
rect 9220 18207 9272 18216
rect 9220 18173 9229 18207
rect 9229 18173 9263 18207
rect 9263 18173 9272 18207
rect 9220 18164 9272 18173
rect 10048 18096 10100 18148
rect 3884 18071 3936 18080
rect 3884 18037 3893 18071
rect 3893 18037 3927 18071
rect 3927 18037 3936 18071
rect 3884 18028 3936 18037
rect 4252 18028 4304 18080
rect 8760 18028 8812 18080
rect 10140 18028 10192 18080
rect 10876 18275 10928 18284
rect 10876 18241 10885 18275
rect 10885 18241 10919 18275
rect 10919 18241 10928 18275
rect 10876 18232 10928 18241
rect 12072 18309 12091 18343
rect 12091 18309 12124 18343
rect 13268 18368 13320 18420
rect 14832 18368 14884 18420
rect 15752 18368 15804 18420
rect 16488 18368 16540 18420
rect 17408 18368 17460 18420
rect 12072 18300 12124 18309
rect 11796 18275 11848 18284
rect 11796 18241 11805 18275
rect 11805 18241 11839 18275
rect 11839 18241 11848 18275
rect 11796 18232 11848 18241
rect 14004 18300 14056 18352
rect 12900 18275 12952 18284
rect 12900 18241 12909 18275
rect 12909 18241 12943 18275
rect 12943 18241 12952 18275
rect 12900 18232 12952 18241
rect 14096 18275 14148 18284
rect 14096 18241 14105 18275
rect 14105 18241 14139 18275
rect 14139 18241 14148 18275
rect 14096 18232 14148 18241
rect 15108 18275 15160 18284
rect 15108 18241 15117 18275
rect 15117 18241 15151 18275
rect 15151 18241 15160 18275
rect 15108 18232 15160 18241
rect 15200 18275 15252 18284
rect 15200 18241 15209 18275
rect 15209 18241 15243 18275
rect 15243 18241 15252 18275
rect 15200 18232 15252 18241
rect 11704 18164 11756 18216
rect 12072 18164 12124 18216
rect 13084 18164 13136 18216
rect 13820 18164 13872 18216
rect 15016 18164 15068 18216
rect 15936 18232 15988 18284
rect 17776 18232 17828 18284
rect 18328 18275 18380 18284
rect 16488 18164 16540 18216
rect 17868 18164 17920 18216
rect 18328 18241 18337 18275
rect 18337 18241 18371 18275
rect 18371 18241 18380 18275
rect 18328 18232 18380 18241
rect 18604 18368 18656 18420
rect 18880 18300 18932 18352
rect 19524 18368 19576 18420
rect 20536 18411 20588 18420
rect 20536 18377 20545 18411
rect 20545 18377 20579 18411
rect 20579 18377 20588 18411
rect 20536 18368 20588 18377
rect 20904 18368 20956 18420
rect 22100 18368 22152 18420
rect 24676 18368 24728 18420
rect 20812 18300 20864 18352
rect 23940 18300 23992 18352
rect 26516 18300 26568 18352
rect 18972 18232 19024 18284
rect 19432 18232 19484 18284
rect 19616 18275 19668 18284
rect 19616 18241 19625 18275
rect 19625 18241 19659 18275
rect 19659 18241 19668 18275
rect 19616 18232 19668 18241
rect 19708 18232 19760 18284
rect 20904 18275 20956 18284
rect 20904 18241 20913 18275
rect 20913 18241 20947 18275
rect 20947 18241 20956 18275
rect 20904 18232 20956 18241
rect 22192 18232 22244 18284
rect 26976 18275 27028 18284
rect 12624 18096 12676 18148
rect 18880 18164 18932 18216
rect 19892 18207 19944 18216
rect 19892 18173 19901 18207
rect 19901 18173 19935 18207
rect 19935 18173 19944 18207
rect 19892 18164 19944 18173
rect 19984 18164 20036 18216
rect 21824 18164 21876 18216
rect 26976 18241 26985 18275
rect 26985 18241 27019 18275
rect 27019 18241 27028 18275
rect 26976 18232 27028 18241
rect 27344 18232 27396 18284
rect 20812 18096 20864 18148
rect 21180 18096 21232 18148
rect 21916 18096 21968 18148
rect 24860 18164 24912 18216
rect 25044 18207 25096 18216
rect 25044 18173 25053 18207
rect 25053 18173 25087 18207
rect 25087 18173 25096 18207
rect 25044 18164 25096 18173
rect 27252 18164 27304 18216
rect 11152 18028 11204 18080
rect 11796 18028 11848 18080
rect 12532 18071 12584 18080
rect 12532 18037 12541 18071
rect 12541 18037 12575 18071
rect 12575 18037 12584 18071
rect 12532 18028 12584 18037
rect 13268 18028 13320 18080
rect 15200 18028 15252 18080
rect 17868 18028 17920 18080
rect 19984 18028 20036 18080
rect 21088 18028 21140 18080
rect 23940 18028 23992 18080
rect 25320 18028 25372 18080
rect 27160 18028 27212 18080
rect 5442 17926 5494 17978
rect 5506 17926 5558 17978
rect 5570 17926 5622 17978
rect 5634 17926 5686 17978
rect 5698 17926 5750 17978
rect 14428 17926 14480 17978
rect 14492 17926 14544 17978
rect 14556 17926 14608 17978
rect 14620 17926 14672 17978
rect 14684 17926 14736 17978
rect 23413 17926 23465 17978
rect 23477 17926 23529 17978
rect 23541 17926 23593 17978
rect 23605 17926 23657 17978
rect 23669 17926 23721 17978
rect 2596 17824 2648 17876
rect 6460 17867 6512 17876
rect 3608 17688 3660 17740
rect 4896 17688 4948 17740
rect 5632 17688 5684 17740
rect 6460 17833 6469 17867
rect 6469 17833 6503 17867
rect 6503 17833 6512 17867
rect 6460 17824 6512 17833
rect 1952 17620 2004 17672
rect 3884 17620 3936 17672
rect 5908 17620 5960 17672
rect 6644 17620 6696 17672
rect 8300 17824 8352 17876
rect 9404 17824 9456 17876
rect 11520 17824 11572 17876
rect 13176 17824 13228 17876
rect 13268 17824 13320 17876
rect 13728 17824 13780 17876
rect 14832 17824 14884 17876
rect 15660 17824 15712 17876
rect 15936 17824 15988 17876
rect 16396 17824 16448 17876
rect 17224 17824 17276 17876
rect 21824 17824 21876 17876
rect 23204 17824 23256 17876
rect 24032 17824 24084 17876
rect 15108 17756 15160 17808
rect 19064 17756 19116 17808
rect 20076 17756 20128 17808
rect 20720 17756 20772 17808
rect 8300 17688 8352 17740
rect 18880 17688 18932 17740
rect 19984 17688 20036 17740
rect 21548 17688 21600 17740
rect 3608 17552 3660 17604
rect 5356 17552 5408 17604
rect 8668 17620 8720 17672
rect 8944 17620 8996 17672
rect 10784 17620 10836 17672
rect 17960 17620 18012 17672
rect 18788 17620 18840 17672
rect 8576 17552 8628 17604
rect 9588 17552 9640 17604
rect 12532 17552 12584 17604
rect 13728 17552 13780 17604
rect 15016 17552 15068 17604
rect 16488 17552 16540 17604
rect 17592 17595 17644 17604
rect 17592 17561 17626 17595
rect 17626 17561 17644 17595
rect 17592 17552 17644 17561
rect 20812 17620 20864 17672
rect 4896 17484 4948 17536
rect 5540 17484 5592 17536
rect 5724 17484 5776 17536
rect 10508 17484 10560 17536
rect 10876 17527 10928 17536
rect 10876 17493 10885 17527
rect 10885 17493 10919 17527
rect 10919 17493 10928 17527
rect 10876 17484 10928 17493
rect 11520 17484 11572 17536
rect 11796 17484 11848 17536
rect 20628 17552 20680 17604
rect 21088 17663 21140 17672
rect 21088 17629 21097 17663
rect 21097 17629 21131 17663
rect 21131 17629 21140 17663
rect 21088 17620 21140 17629
rect 26884 17688 26936 17740
rect 21916 17620 21968 17672
rect 25044 17620 25096 17672
rect 25780 17620 25832 17672
rect 26516 17620 26568 17672
rect 22100 17552 22152 17604
rect 23112 17552 23164 17604
rect 24216 17552 24268 17604
rect 17776 17484 17828 17536
rect 21088 17484 21140 17536
rect 23296 17484 23348 17536
rect 24860 17484 24912 17536
rect 26332 17484 26384 17536
rect 26792 17484 26844 17536
rect 9935 17382 9987 17434
rect 9999 17382 10051 17434
rect 10063 17382 10115 17434
rect 10127 17382 10179 17434
rect 10191 17382 10243 17434
rect 18920 17382 18972 17434
rect 18984 17382 19036 17434
rect 19048 17382 19100 17434
rect 19112 17382 19164 17434
rect 19176 17382 19228 17434
rect 2504 17280 2556 17332
rect 3424 17212 3476 17264
rect 5724 17280 5776 17332
rect 9588 17323 9640 17332
rect 9588 17289 9597 17323
rect 9597 17289 9631 17323
rect 9631 17289 9640 17323
rect 9588 17280 9640 17289
rect 12164 17280 12216 17332
rect 13176 17280 13228 17332
rect 13728 17323 13780 17332
rect 13728 17289 13737 17323
rect 13737 17289 13771 17323
rect 13771 17289 13780 17323
rect 13728 17280 13780 17289
rect 4896 17212 4948 17264
rect 5540 17255 5592 17264
rect 5540 17221 5549 17255
rect 5549 17221 5583 17255
rect 5583 17221 5592 17255
rect 5540 17212 5592 17221
rect 5356 17187 5408 17196
rect 1952 17119 2004 17128
rect 1952 17085 1961 17119
rect 1961 17085 1995 17119
rect 1995 17085 2004 17119
rect 1952 17076 2004 17085
rect 4160 17076 4212 17128
rect 5356 17153 5365 17187
rect 5365 17153 5399 17187
rect 5399 17153 5408 17187
rect 5356 17144 5408 17153
rect 5632 17144 5684 17196
rect 6276 17144 6328 17196
rect 8300 17187 8352 17196
rect 8300 17153 8309 17187
rect 8309 17153 8343 17187
rect 8343 17153 8352 17187
rect 8300 17144 8352 17153
rect 9220 17144 9272 17196
rect 11336 17212 11388 17264
rect 11796 17212 11848 17264
rect 16764 17280 16816 17332
rect 17592 17323 17644 17332
rect 17592 17289 17601 17323
rect 17601 17289 17635 17323
rect 17635 17289 17644 17323
rect 17592 17280 17644 17289
rect 5816 17076 5868 17128
rect 6368 17119 6420 17128
rect 6368 17085 6377 17119
rect 6377 17085 6411 17119
rect 6411 17085 6420 17119
rect 6368 17076 6420 17085
rect 8576 17119 8628 17128
rect 8576 17085 8585 17119
rect 8585 17085 8619 17119
rect 8619 17085 8628 17119
rect 8576 17076 8628 17085
rect 4620 17008 4672 17060
rect 4528 16940 4580 16992
rect 4712 16940 4764 16992
rect 4988 16940 5040 16992
rect 7380 16940 7432 16992
rect 9680 16940 9732 16992
rect 10508 17144 10560 17196
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 12164 17187 12216 17196
rect 10968 17076 11020 17128
rect 12164 17153 12173 17187
rect 12173 17153 12207 17187
rect 12207 17153 12216 17187
rect 12164 17144 12216 17153
rect 12808 17187 12860 17196
rect 12808 17153 12817 17187
rect 12817 17153 12851 17187
rect 12851 17153 12860 17187
rect 12808 17144 12860 17153
rect 13084 17187 13136 17196
rect 13084 17153 13093 17187
rect 13093 17153 13127 17187
rect 13127 17153 13136 17187
rect 13084 17144 13136 17153
rect 13544 17144 13596 17196
rect 13728 17144 13780 17196
rect 14832 17212 14884 17264
rect 15016 17212 15068 17264
rect 19524 17280 19576 17332
rect 20812 17280 20864 17332
rect 24216 17323 24268 17332
rect 18788 17255 18840 17264
rect 14372 17187 14424 17196
rect 13268 17076 13320 17128
rect 14372 17153 14381 17187
rect 14381 17153 14415 17187
rect 14415 17153 14424 17187
rect 14372 17144 14424 17153
rect 18788 17221 18797 17255
rect 18797 17221 18831 17255
rect 18831 17221 18840 17255
rect 18788 17212 18840 17221
rect 19708 17212 19760 17264
rect 20168 17212 20220 17264
rect 15936 17187 15988 17196
rect 15936 17153 15945 17187
rect 15945 17153 15979 17187
rect 15979 17153 15988 17187
rect 15936 17144 15988 17153
rect 17316 17144 17368 17196
rect 18512 17144 18564 17196
rect 18696 17144 18748 17196
rect 16396 17076 16448 17128
rect 17224 17076 17276 17128
rect 17684 17076 17736 17128
rect 10968 16940 11020 16992
rect 12164 17008 12216 17060
rect 16488 17008 16540 17060
rect 17776 17008 17828 17060
rect 19340 17076 19392 17128
rect 20536 17144 20588 17196
rect 21180 17144 21232 17196
rect 22100 17212 22152 17264
rect 20076 17076 20128 17128
rect 21088 17076 21140 17128
rect 18972 17008 19024 17060
rect 20812 17008 20864 17060
rect 12532 16940 12584 16992
rect 16856 16940 16908 16992
rect 17316 16940 17368 16992
rect 18052 16940 18104 16992
rect 22100 17119 22152 17128
rect 22100 17085 22109 17119
rect 22109 17085 22143 17119
rect 22143 17085 22152 17119
rect 22652 17144 22704 17196
rect 23020 17187 23072 17196
rect 23020 17153 23029 17187
rect 23029 17153 23063 17187
rect 23063 17153 23072 17187
rect 23020 17144 23072 17153
rect 23204 17187 23256 17196
rect 23204 17153 23213 17187
rect 23213 17153 23247 17187
rect 23247 17153 23256 17187
rect 23204 17144 23256 17153
rect 24216 17289 24225 17323
rect 24225 17289 24259 17323
rect 24259 17289 24268 17323
rect 24216 17280 24268 17289
rect 26240 17280 26292 17332
rect 26700 17280 26752 17332
rect 26976 17280 27028 17332
rect 23664 17144 23716 17196
rect 24676 17187 24728 17196
rect 24676 17153 24685 17187
rect 24685 17153 24719 17187
rect 24719 17153 24728 17187
rect 24676 17144 24728 17153
rect 24860 17144 24912 17196
rect 25136 17144 25188 17196
rect 25964 17144 26016 17196
rect 22100 17076 22152 17085
rect 24032 17076 24084 17128
rect 24308 17076 24360 17128
rect 23296 16940 23348 16992
rect 26240 17076 26292 17128
rect 25964 17008 26016 17060
rect 26516 16940 26568 16992
rect 5442 16838 5494 16890
rect 5506 16838 5558 16890
rect 5570 16838 5622 16890
rect 5634 16838 5686 16890
rect 5698 16838 5750 16890
rect 14428 16838 14480 16890
rect 14492 16838 14544 16890
rect 14556 16838 14608 16890
rect 14620 16838 14672 16890
rect 14684 16838 14736 16890
rect 23413 16838 23465 16890
rect 23477 16838 23529 16890
rect 23541 16838 23593 16890
rect 23605 16838 23657 16890
rect 23669 16838 23721 16890
rect 3608 16736 3660 16788
rect 6276 16779 6328 16788
rect 6276 16745 6285 16779
rect 6285 16745 6319 16779
rect 6319 16745 6328 16779
rect 6276 16736 6328 16745
rect 11612 16736 11664 16788
rect 12808 16736 12860 16788
rect 15936 16736 15988 16788
rect 1032 16668 1084 16720
rect 1400 16668 1452 16720
rect 2872 16600 2924 16652
rect 3608 16600 3660 16652
rect 5816 16600 5868 16652
rect 8944 16600 8996 16652
rect 1400 16532 1452 16584
rect 1952 16532 2004 16584
rect 4252 16532 4304 16584
rect 4988 16575 5040 16584
rect 4988 16541 4997 16575
rect 4997 16541 5031 16575
rect 5031 16541 5040 16575
rect 4988 16532 5040 16541
rect 5172 16532 5224 16584
rect 7564 16532 7616 16584
rect 8392 16532 8444 16584
rect 9680 16532 9732 16584
rect 13544 16668 13596 16720
rect 14004 16668 14056 16720
rect 16212 16668 16264 16720
rect 13360 16532 13412 16584
rect 4068 16396 4120 16448
rect 5448 16439 5500 16448
rect 5448 16405 5457 16439
rect 5457 16405 5491 16439
rect 5491 16405 5500 16439
rect 5448 16396 5500 16405
rect 6276 16396 6328 16448
rect 6736 16396 6788 16448
rect 8208 16396 8260 16448
rect 9588 16464 9640 16516
rect 10692 16464 10744 16516
rect 10968 16464 11020 16516
rect 12164 16464 12216 16516
rect 15936 16600 15988 16652
rect 12440 16439 12492 16448
rect 12440 16405 12449 16439
rect 12449 16405 12483 16439
rect 12483 16405 12492 16439
rect 13728 16464 13780 16516
rect 14832 16532 14884 16584
rect 15384 16575 15436 16584
rect 15384 16541 15391 16575
rect 15391 16541 15436 16575
rect 15384 16532 15436 16541
rect 15660 16575 15712 16584
rect 15660 16541 15674 16575
rect 15674 16541 15708 16575
rect 15708 16541 15712 16575
rect 15660 16532 15712 16541
rect 14372 16507 14424 16516
rect 14372 16473 14381 16507
rect 14381 16473 14415 16507
rect 14415 16473 14424 16507
rect 14372 16464 14424 16473
rect 12440 16396 12492 16405
rect 15016 16464 15068 16516
rect 15752 16464 15804 16516
rect 15936 16464 15988 16516
rect 17316 16736 17368 16788
rect 19616 16736 19668 16788
rect 22008 16736 22060 16788
rect 25136 16779 25188 16788
rect 25136 16745 25145 16779
rect 25145 16745 25179 16779
rect 25179 16745 25188 16779
rect 25136 16736 25188 16745
rect 17224 16668 17276 16720
rect 18052 16668 18104 16720
rect 18512 16668 18564 16720
rect 16948 16532 17000 16584
rect 19340 16600 19392 16652
rect 20812 16668 20864 16720
rect 21824 16668 21876 16720
rect 22100 16668 22152 16720
rect 22652 16668 22704 16720
rect 24032 16668 24084 16720
rect 22928 16600 22980 16652
rect 23020 16600 23072 16652
rect 24216 16600 24268 16652
rect 25044 16600 25096 16652
rect 25964 16643 26016 16652
rect 25964 16609 25973 16643
rect 25973 16609 26007 16643
rect 26007 16609 26016 16643
rect 25964 16600 26016 16609
rect 17776 16532 17828 16584
rect 18144 16532 18196 16584
rect 18512 16532 18564 16584
rect 19432 16532 19484 16584
rect 21180 16575 21232 16584
rect 21180 16541 21189 16575
rect 21189 16541 21223 16575
rect 21223 16541 21232 16575
rect 21180 16532 21232 16541
rect 18788 16464 18840 16516
rect 22008 16532 22060 16584
rect 24400 16575 24452 16584
rect 24400 16541 24409 16575
rect 24409 16541 24443 16575
rect 24443 16541 24452 16575
rect 24400 16532 24452 16541
rect 26240 16575 26292 16584
rect 26240 16541 26274 16575
rect 26274 16541 26292 16575
rect 23204 16464 23256 16516
rect 24676 16464 24728 16516
rect 17408 16396 17460 16448
rect 17776 16396 17828 16448
rect 17868 16396 17920 16448
rect 18144 16396 18196 16448
rect 20168 16396 20220 16448
rect 21088 16396 21140 16448
rect 22008 16396 22060 16448
rect 24124 16396 24176 16448
rect 26240 16532 26292 16541
rect 25228 16396 25280 16448
rect 25872 16396 25924 16448
rect 9935 16294 9987 16346
rect 9999 16294 10051 16346
rect 10063 16294 10115 16346
rect 10127 16294 10179 16346
rect 10191 16294 10243 16346
rect 18920 16294 18972 16346
rect 18984 16294 19036 16346
rect 19048 16294 19100 16346
rect 19112 16294 19164 16346
rect 19176 16294 19228 16346
rect 4988 16192 5040 16244
rect 7564 16235 7616 16244
rect 7564 16201 7573 16235
rect 7573 16201 7607 16235
rect 7607 16201 7616 16235
rect 7564 16192 7616 16201
rect 8392 16235 8444 16244
rect 1952 16124 2004 16176
rect 2504 16099 2556 16108
rect 2504 16065 2513 16099
rect 2513 16065 2547 16099
rect 2547 16065 2556 16099
rect 2504 16056 2556 16065
rect 2780 16056 2832 16108
rect 3516 16099 3568 16108
rect 3516 16065 3525 16099
rect 3525 16065 3559 16099
rect 3559 16065 3568 16099
rect 3516 16056 3568 16065
rect 5816 16124 5868 16176
rect 5448 16056 5500 16108
rect 6736 16056 6788 16108
rect 7932 16124 7984 16176
rect 8392 16201 8401 16235
rect 8401 16201 8435 16235
rect 8435 16201 8444 16235
rect 8392 16192 8444 16201
rect 12256 16192 12308 16244
rect 8668 16124 8720 16176
rect 9404 16124 9456 16176
rect 13728 16192 13780 16244
rect 14372 16192 14424 16244
rect 8944 16099 8996 16108
rect 8944 16065 8953 16099
rect 8953 16065 8987 16099
rect 8987 16065 8996 16099
rect 8944 16056 8996 16065
rect 10784 16099 10836 16108
rect 10784 16065 10793 16099
rect 10793 16065 10827 16099
rect 10827 16065 10836 16099
rect 10784 16056 10836 16065
rect 11612 16056 11664 16108
rect 12164 16099 12216 16108
rect 12164 16065 12173 16099
rect 12173 16065 12207 16099
rect 12207 16065 12216 16099
rect 12164 16056 12216 16065
rect 13084 16056 13136 16108
rect 13544 16099 13596 16108
rect 13176 15988 13228 16040
rect 13544 16065 13553 16099
rect 13553 16065 13587 16099
rect 13587 16065 13596 16099
rect 13544 16056 13596 16065
rect 13820 16056 13872 16108
rect 14372 16099 14424 16108
rect 14372 16065 14381 16099
rect 14381 16065 14415 16099
rect 14415 16065 14424 16099
rect 14372 16056 14424 16065
rect 15016 15988 15068 16040
rect 2412 15852 2464 15904
rect 2872 15895 2924 15904
rect 2872 15861 2881 15895
rect 2881 15861 2915 15895
rect 2915 15861 2924 15895
rect 2872 15852 2924 15861
rect 3884 15852 3936 15904
rect 6368 15895 6420 15904
rect 6368 15861 6377 15895
rect 6377 15861 6411 15895
rect 6411 15861 6420 15895
rect 6368 15852 6420 15861
rect 7380 15895 7432 15904
rect 7380 15861 7389 15895
rect 7389 15861 7423 15895
rect 7423 15861 7432 15895
rect 7380 15852 7432 15861
rect 8208 15895 8260 15904
rect 8208 15861 8217 15895
rect 8217 15861 8251 15895
rect 8251 15861 8260 15895
rect 8208 15852 8260 15861
rect 10140 15920 10192 15972
rect 21824 16192 21876 16244
rect 16212 16124 16264 16176
rect 16856 16099 16908 16108
rect 16856 16065 16865 16099
rect 16865 16065 16899 16099
rect 16899 16065 16908 16099
rect 16856 16056 16908 16065
rect 17776 16056 17828 16108
rect 17960 16099 18012 16108
rect 17960 16065 17969 16099
rect 17969 16065 18003 16099
rect 18003 16065 18012 16099
rect 17960 16056 18012 16065
rect 18052 16056 18104 16108
rect 20628 16124 20680 16176
rect 23756 16192 23808 16244
rect 24032 16192 24084 16244
rect 24676 16192 24728 16244
rect 25780 16235 25832 16244
rect 19892 16056 19944 16108
rect 22928 16124 22980 16176
rect 16120 16031 16172 16040
rect 16120 15997 16129 16031
rect 16129 15997 16163 16031
rect 16163 15997 16172 16031
rect 16120 15988 16172 15997
rect 17132 16031 17184 16040
rect 17132 15997 17141 16031
rect 17141 15997 17175 16031
rect 17175 15997 17184 16031
rect 17132 15988 17184 15997
rect 15936 15920 15988 15972
rect 19340 15963 19392 15972
rect 9128 15852 9180 15904
rect 10324 15895 10376 15904
rect 10324 15861 10333 15895
rect 10333 15861 10367 15895
rect 10367 15861 10376 15895
rect 10324 15852 10376 15861
rect 13544 15852 13596 15904
rect 13912 15895 13964 15904
rect 13912 15861 13921 15895
rect 13921 15861 13955 15895
rect 13955 15861 13964 15895
rect 13912 15852 13964 15861
rect 16856 15852 16908 15904
rect 19340 15929 19349 15963
rect 19349 15929 19383 15963
rect 19383 15929 19392 15963
rect 19340 15920 19392 15929
rect 23204 16056 23256 16108
rect 25136 16124 25188 16176
rect 24400 16056 24452 16108
rect 24676 16056 24728 16108
rect 25412 16124 25464 16176
rect 25780 16201 25789 16235
rect 25789 16201 25823 16235
rect 25823 16201 25832 16235
rect 25780 16192 25832 16201
rect 26516 16192 26568 16244
rect 21916 16031 21968 16040
rect 21916 15997 21925 16031
rect 21925 15997 21959 16031
rect 21959 15997 21968 16031
rect 21916 15988 21968 15997
rect 23756 16031 23808 16040
rect 23756 15997 23765 16031
rect 23765 15997 23799 16031
rect 23799 15997 23808 16031
rect 23756 15988 23808 15997
rect 25872 16056 25924 16108
rect 26516 16056 26568 16108
rect 25688 15920 25740 15972
rect 21180 15895 21232 15904
rect 21180 15861 21189 15895
rect 21189 15861 21223 15895
rect 21223 15861 21232 15895
rect 21180 15852 21232 15861
rect 23112 15852 23164 15904
rect 26240 15895 26292 15904
rect 26240 15861 26249 15895
rect 26249 15861 26283 15895
rect 26283 15861 26292 15895
rect 26240 15852 26292 15861
rect 5442 15750 5494 15802
rect 5506 15750 5558 15802
rect 5570 15750 5622 15802
rect 5634 15750 5686 15802
rect 5698 15750 5750 15802
rect 14428 15750 14480 15802
rect 14492 15750 14544 15802
rect 14556 15750 14608 15802
rect 14620 15750 14672 15802
rect 14684 15750 14736 15802
rect 23413 15750 23465 15802
rect 23477 15750 23529 15802
rect 23541 15750 23593 15802
rect 23605 15750 23657 15802
rect 23669 15750 23721 15802
rect 2780 15691 2832 15700
rect 2780 15657 2789 15691
rect 2789 15657 2823 15691
rect 2823 15657 2832 15691
rect 4160 15691 4212 15700
rect 2780 15648 2832 15657
rect 4160 15657 4169 15691
rect 4169 15657 4203 15691
rect 4203 15657 4212 15691
rect 4160 15648 4212 15657
rect 4988 15691 5040 15700
rect 4988 15657 4997 15691
rect 4997 15657 5031 15691
rect 5031 15657 5040 15691
rect 4988 15648 5040 15657
rect 5172 15691 5224 15700
rect 5172 15657 5181 15691
rect 5181 15657 5215 15691
rect 5215 15657 5224 15691
rect 5172 15648 5224 15657
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 2504 15512 2556 15564
rect 5816 15648 5868 15700
rect 7380 15648 7432 15700
rect 7840 15648 7892 15700
rect 7932 15648 7984 15700
rect 10140 15648 10192 15700
rect 10600 15691 10652 15700
rect 10600 15657 10609 15691
rect 10609 15657 10643 15691
rect 10643 15657 10652 15691
rect 10600 15648 10652 15657
rect 13360 15648 13412 15700
rect 7472 15580 7524 15632
rect 7656 15580 7708 15632
rect 9220 15580 9272 15632
rect 10508 15580 10560 15632
rect 12348 15580 12400 15632
rect 7012 15512 7064 15564
rect 7840 15512 7892 15564
rect 10600 15512 10652 15564
rect 10784 15512 10836 15564
rect 11244 15512 11296 15564
rect 11796 15512 11848 15564
rect 12624 15512 12676 15564
rect 15108 15580 15160 15632
rect 12808 15512 12860 15564
rect 1860 15376 1912 15428
rect 4436 15376 4488 15428
rect 6368 15444 6420 15496
rect 6460 15444 6512 15496
rect 9588 15444 9640 15496
rect 10324 15444 10376 15496
rect 11152 15487 11204 15496
rect 11152 15453 11161 15487
rect 11161 15453 11195 15487
rect 11195 15453 11204 15487
rect 11152 15444 11204 15453
rect 13728 15444 13780 15496
rect 14188 15444 14240 15496
rect 14372 15444 14424 15496
rect 14740 15487 14792 15496
rect 14740 15453 14749 15487
rect 14749 15453 14783 15487
rect 14783 15453 14792 15487
rect 14740 15444 14792 15453
rect 15016 15487 15068 15496
rect 15016 15453 15025 15487
rect 15025 15453 15059 15487
rect 15059 15453 15068 15487
rect 15016 15444 15068 15453
rect 15844 15648 15896 15700
rect 16028 15691 16080 15700
rect 16028 15657 16037 15691
rect 16037 15657 16071 15691
rect 16071 15657 16080 15691
rect 16028 15648 16080 15657
rect 16212 15648 16264 15700
rect 16948 15648 17000 15700
rect 17776 15648 17828 15700
rect 19892 15648 19944 15700
rect 20904 15648 20956 15700
rect 22008 15648 22060 15700
rect 22192 15648 22244 15700
rect 23204 15691 23256 15700
rect 23204 15657 23213 15691
rect 23213 15657 23247 15691
rect 23247 15657 23256 15691
rect 23204 15648 23256 15657
rect 24308 15648 24360 15700
rect 25228 15648 25280 15700
rect 25412 15648 25464 15700
rect 26884 15648 26936 15700
rect 15384 15623 15436 15632
rect 15384 15589 15393 15623
rect 15393 15589 15427 15623
rect 15427 15589 15436 15623
rect 15384 15580 15436 15589
rect 15660 15444 15712 15496
rect 6828 15376 6880 15428
rect 2320 15308 2372 15360
rect 2596 15308 2648 15360
rect 5172 15308 5224 15360
rect 6368 15308 6420 15360
rect 14556 15376 14608 15428
rect 14648 15376 14700 15428
rect 19616 15580 19668 15632
rect 20628 15580 20680 15632
rect 15844 15512 15896 15564
rect 17960 15444 18012 15496
rect 20720 15512 20772 15564
rect 22100 15580 22152 15632
rect 20076 15444 20128 15496
rect 21180 15444 21232 15496
rect 22928 15580 22980 15632
rect 23204 15512 23256 15564
rect 23664 15555 23716 15564
rect 23664 15521 23673 15555
rect 23673 15521 23707 15555
rect 23707 15521 23716 15555
rect 23664 15512 23716 15521
rect 24676 15555 24728 15564
rect 24676 15521 24685 15555
rect 24685 15521 24719 15555
rect 24719 15521 24728 15555
rect 24676 15512 24728 15521
rect 25964 15555 26016 15564
rect 25964 15521 25973 15555
rect 25973 15521 26007 15555
rect 26007 15521 26016 15555
rect 25964 15512 26016 15521
rect 21824 15444 21876 15496
rect 22008 15487 22060 15496
rect 22008 15453 22017 15487
rect 22017 15453 22051 15487
rect 22051 15453 22060 15487
rect 22008 15444 22060 15453
rect 22192 15487 22244 15496
rect 22192 15453 22201 15487
rect 22201 15453 22235 15487
rect 22235 15453 22244 15487
rect 22192 15444 22244 15453
rect 21088 15376 21140 15428
rect 23296 15444 23348 15496
rect 23848 15444 23900 15496
rect 26332 15376 26384 15428
rect 8300 15308 8352 15360
rect 15936 15308 15988 15360
rect 16948 15308 17000 15360
rect 19340 15308 19392 15360
rect 20628 15308 20680 15360
rect 20720 15308 20772 15360
rect 22192 15308 22244 15360
rect 23848 15308 23900 15360
rect 25228 15308 25280 15360
rect 25872 15308 25924 15360
rect 9935 15206 9987 15258
rect 9999 15206 10051 15258
rect 10063 15206 10115 15258
rect 10127 15206 10179 15258
rect 10191 15206 10243 15258
rect 18920 15206 18972 15258
rect 18984 15206 19036 15258
rect 19048 15206 19100 15258
rect 19112 15206 19164 15258
rect 19176 15206 19228 15258
rect 1400 15104 1452 15156
rect 1676 15104 1728 15156
rect 1860 15147 1912 15156
rect 1860 15113 1869 15147
rect 1869 15113 1903 15147
rect 1903 15113 1912 15147
rect 1860 15104 1912 15113
rect 5172 15147 5224 15156
rect 2872 15036 2924 15088
rect 3792 14968 3844 15020
rect 5172 15113 5207 15147
rect 5207 15113 5224 15147
rect 5172 15104 5224 15113
rect 6460 15104 6512 15156
rect 6736 15147 6788 15156
rect 6736 15113 6745 15147
rect 6745 15113 6779 15147
rect 6779 15113 6788 15147
rect 6736 15104 6788 15113
rect 6828 15104 6880 15156
rect 8300 15104 8352 15156
rect 4436 15036 4488 15088
rect 9220 15104 9272 15156
rect 2688 14832 2740 14884
rect 4160 14832 4212 14884
rect 4344 14764 4396 14816
rect 6368 14764 6420 14816
rect 7932 14968 7984 15020
rect 8208 14968 8260 15020
rect 8300 14900 8352 14952
rect 8668 14968 8720 15020
rect 9772 15036 9824 15088
rect 13728 15104 13780 15156
rect 9680 14968 9732 15020
rect 10600 14968 10652 15020
rect 11336 14968 11388 15020
rect 10876 14900 10928 14952
rect 11428 14900 11480 14952
rect 12348 15036 12400 15088
rect 13360 15036 13412 15088
rect 15844 15147 15896 15156
rect 15844 15113 15869 15147
rect 15869 15113 15896 15147
rect 15844 15104 15896 15113
rect 19340 15104 19392 15156
rect 12624 14968 12676 15020
rect 13084 14968 13136 15020
rect 13728 14968 13780 15020
rect 11704 14900 11756 14952
rect 9864 14832 9916 14884
rect 10784 14832 10836 14884
rect 13268 14900 13320 14952
rect 12164 14832 12216 14884
rect 7840 14764 7892 14816
rect 9680 14764 9732 14816
rect 11336 14764 11388 14816
rect 11704 14807 11756 14816
rect 11704 14773 11713 14807
rect 11713 14773 11747 14807
rect 11747 14773 11756 14807
rect 11704 14764 11756 14773
rect 13084 14807 13136 14816
rect 13084 14773 13093 14807
rect 13093 14773 13127 14807
rect 13127 14773 13136 14807
rect 13084 14764 13136 14773
rect 14832 14968 14884 15020
rect 15384 14832 15436 14884
rect 15016 14807 15068 14816
rect 15016 14773 15025 14807
rect 15025 14773 15059 14807
rect 15059 14773 15068 14807
rect 15016 14764 15068 14773
rect 16580 14968 16632 15020
rect 16856 14968 16908 15020
rect 17408 14968 17460 15020
rect 17960 14968 18012 15020
rect 18696 14968 18748 15020
rect 17868 14900 17920 14952
rect 19892 14900 19944 14952
rect 20720 15036 20772 15088
rect 20812 14968 20864 15020
rect 21180 14900 21232 14952
rect 16212 14832 16264 14884
rect 16672 14832 16724 14884
rect 16856 14832 16908 14884
rect 22192 14968 22244 15020
rect 23112 15011 23164 15020
rect 23112 14977 23121 15011
rect 23121 14977 23155 15011
rect 23155 14977 23164 15011
rect 23112 14968 23164 14977
rect 24400 14968 24452 15020
rect 24676 14968 24728 15020
rect 25688 15011 25740 15020
rect 25688 14977 25697 15011
rect 25697 14977 25731 15011
rect 25731 14977 25740 15011
rect 25688 14968 25740 14977
rect 26148 14968 26200 15020
rect 22560 14900 22612 14952
rect 23296 14943 23348 14952
rect 23296 14909 23305 14943
rect 23305 14909 23339 14943
rect 23339 14909 23348 14943
rect 23296 14900 23348 14909
rect 16028 14764 16080 14816
rect 16396 14764 16448 14816
rect 23204 14832 23256 14884
rect 25136 14900 25188 14952
rect 23480 14832 23532 14884
rect 25872 14943 25924 14952
rect 25872 14909 25881 14943
rect 25881 14909 25915 14943
rect 25915 14909 25924 14943
rect 25872 14900 25924 14909
rect 19156 14764 19208 14816
rect 21088 14807 21140 14816
rect 21088 14773 21097 14807
rect 21097 14773 21131 14807
rect 21131 14773 21140 14807
rect 21088 14764 21140 14773
rect 21824 14807 21876 14816
rect 21824 14773 21833 14807
rect 21833 14773 21867 14807
rect 21867 14773 21876 14807
rect 21824 14764 21876 14773
rect 22928 14764 22980 14816
rect 24216 14764 24268 14816
rect 5442 14662 5494 14714
rect 5506 14662 5558 14714
rect 5570 14662 5622 14714
rect 5634 14662 5686 14714
rect 5698 14662 5750 14714
rect 14428 14662 14480 14714
rect 14492 14662 14544 14714
rect 14556 14662 14608 14714
rect 14620 14662 14672 14714
rect 14684 14662 14736 14714
rect 23413 14662 23465 14714
rect 23477 14662 23529 14714
rect 23541 14662 23593 14714
rect 23605 14662 23657 14714
rect 23669 14662 23721 14714
rect 3792 14603 3844 14612
rect 3792 14569 3801 14603
rect 3801 14569 3835 14603
rect 3835 14569 3844 14603
rect 3792 14560 3844 14569
rect 8852 14560 8904 14612
rect 9036 14560 9088 14612
rect 9772 14560 9824 14612
rect 9864 14492 9916 14544
rect 4344 14424 4396 14476
rect 8392 14424 8444 14476
rect 2044 14356 2096 14408
rect 4160 14356 4212 14408
rect 4252 14356 4304 14408
rect 1676 14331 1728 14340
rect 1676 14297 1710 14331
rect 1710 14297 1728 14331
rect 1676 14288 1728 14297
rect 3148 14288 3200 14340
rect 6276 14356 6328 14408
rect 7196 14356 7248 14408
rect 7748 14356 7800 14408
rect 8668 14356 8720 14408
rect 9772 14356 9824 14408
rect 11704 14560 11756 14612
rect 12348 14560 12400 14612
rect 13084 14560 13136 14612
rect 16028 14560 16080 14612
rect 16580 14560 16632 14612
rect 11152 14492 11204 14544
rect 10692 14424 10744 14476
rect 10968 14424 11020 14476
rect 12164 14424 12216 14476
rect 13912 14424 13964 14476
rect 15016 14492 15068 14544
rect 17592 14492 17644 14544
rect 10324 14399 10376 14408
rect 10324 14365 10333 14399
rect 10333 14365 10367 14399
rect 10367 14365 10376 14399
rect 10324 14356 10376 14365
rect 10600 14356 10652 14408
rect 11520 14356 11572 14408
rect 6460 14288 6512 14340
rect 6736 14331 6788 14340
rect 6736 14297 6770 14331
rect 6770 14297 6788 14331
rect 6736 14288 6788 14297
rect 9496 14288 9548 14340
rect 11336 14288 11388 14340
rect 11888 14288 11940 14340
rect 12624 14331 12676 14340
rect 12624 14297 12649 14331
rect 12649 14297 12676 14331
rect 12624 14288 12676 14297
rect 13176 14288 13228 14340
rect 14464 14356 14516 14408
rect 14832 14424 14884 14476
rect 18788 14560 18840 14612
rect 19892 14560 19944 14612
rect 17868 14492 17920 14544
rect 18052 14492 18104 14544
rect 19616 14492 19668 14544
rect 15936 14399 15988 14408
rect 15936 14365 15945 14399
rect 15945 14365 15979 14399
rect 15979 14365 15988 14399
rect 15936 14356 15988 14365
rect 16028 14356 16080 14408
rect 17224 14356 17276 14408
rect 17868 14399 17920 14408
rect 17868 14365 17877 14399
rect 17877 14365 17911 14399
rect 17911 14365 17920 14399
rect 17868 14356 17920 14365
rect 15016 14288 15068 14340
rect 15200 14288 15252 14340
rect 15844 14288 15896 14340
rect 16672 14288 16724 14340
rect 19340 14424 19392 14476
rect 19524 14424 19576 14476
rect 18696 14356 18748 14408
rect 18788 14356 18840 14408
rect 19156 14288 19208 14340
rect 19340 14331 19392 14340
rect 19340 14297 19349 14331
rect 19349 14297 19383 14331
rect 19383 14297 19392 14331
rect 19340 14288 19392 14297
rect 2872 14220 2924 14272
rect 5080 14263 5132 14272
rect 5080 14229 5089 14263
rect 5089 14229 5123 14263
rect 5123 14229 5132 14263
rect 5080 14220 5132 14229
rect 5816 14263 5868 14272
rect 5816 14229 5825 14263
rect 5825 14229 5859 14263
rect 5859 14229 5868 14263
rect 5816 14220 5868 14229
rect 7012 14220 7064 14272
rect 8208 14220 8260 14272
rect 10600 14220 10652 14272
rect 13268 14220 13320 14272
rect 15476 14263 15528 14272
rect 15476 14229 15485 14263
rect 15485 14229 15519 14263
rect 15519 14229 15528 14263
rect 15476 14220 15528 14229
rect 17776 14220 17828 14272
rect 18420 14220 18472 14272
rect 18512 14220 18564 14272
rect 21548 14560 21600 14612
rect 22284 14603 22336 14612
rect 22284 14569 22293 14603
rect 22293 14569 22327 14603
rect 22327 14569 22336 14603
rect 22284 14560 22336 14569
rect 23112 14560 23164 14612
rect 21824 14492 21876 14544
rect 21548 14424 21600 14476
rect 23296 14424 23348 14476
rect 23756 14424 23808 14476
rect 21916 14356 21968 14408
rect 24216 14356 24268 14408
rect 25964 14467 26016 14476
rect 25964 14433 25973 14467
rect 25973 14433 26007 14467
rect 26007 14433 26016 14467
rect 25964 14424 26016 14433
rect 22284 14288 22336 14340
rect 23664 14331 23716 14340
rect 23664 14297 23673 14331
rect 23673 14297 23707 14331
rect 23707 14297 23716 14331
rect 23664 14288 23716 14297
rect 21548 14263 21600 14272
rect 21548 14229 21557 14263
rect 21557 14229 21591 14263
rect 21591 14229 21600 14263
rect 21548 14220 21600 14229
rect 22100 14220 22152 14272
rect 22928 14220 22980 14272
rect 24308 14288 24360 14340
rect 24216 14220 24268 14272
rect 25872 14288 25924 14340
rect 9935 14118 9987 14170
rect 9999 14118 10051 14170
rect 10063 14118 10115 14170
rect 10127 14118 10179 14170
rect 10191 14118 10243 14170
rect 18920 14118 18972 14170
rect 18984 14118 19036 14170
rect 19048 14118 19100 14170
rect 19112 14118 19164 14170
rect 19176 14118 19228 14170
rect 1676 14059 1728 14068
rect 1676 14025 1685 14059
rect 1685 14025 1719 14059
rect 1719 14025 1728 14059
rect 1676 14016 1728 14025
rect 3148 14016 3200 14068
rect 3976 14016 4028 14068
rect 6736 14059 6788 14068
rect 6736 14025 6745 14059
rect 6745 14025 6779 14059
rect 6779 14025 6788 14059
rect 6736 14016 6788 14025
rect 8668 14016 8720 14068
rect 1860 13923 1912 13932
rect 1860 13889 1869 13923
rect 1869 13889 1903 13923
rect 1903 13889 1912 13923
rect 1860 13880 1912 13889
rect 4344 13948 4396 14000
rect 5816 13948 5868 14000
rect 8300 13948 8352 14000
rect 8484 13948 8536 14000
rect 2872 13923 2924 13932
rect 2872 13889 2906 13923
rect 2906 13889 2924 13923
rect 1676 13812 1728 13864
rect 2044 13812 2096 13864
rect 2872 13880 2924 13889
rect 7748 13880 7800 13932
rect 8392 13880 8444 13932
rect 4344 13812 4396 13864
rect 10692 14016 10744 14068
rect 10784 14059 10836 14068
rect 10784 14025 10793 14059
rect 10793 14025 10827 14059
rect 10827 14025 10836 14059
rect 10784 14016 10836 14025
rect 11520 14016 11572 14068
rect 12624 14016 12676 14068
rect 12716 14016 12768 14068
rect 12900 14016 12952 14068
rect 14464 14059 14516 14068
rect 14464 14025 14473 14059
rect 14473 14025 14507 14059
rect 14507 14025 14516 14059
rect 14464 14016 14516 14025
rect 15016 14016 15068 14068
rect 15292 14059 15344 14068
rect 15292 14025 15301 14059
rect 15301 14025 15335 14059
rect 15335 14025 15344 14059
rect 15292 14016 15344 14025
rect 15476 14016 15528 14068
rect 18512 14016 18564 14068
rect 13544 13948 13596 14000
rect 14648 13948 14700 14000
rect 15660 13948 15712 14000
rect 16580 13948 16632 14000
rect 18788 14016 18840 14068
rect 19248 14016 19300 14068
rect 20720 14016 20772 14068
rect 10692 13880 10744 13932
rect 11428 13880 11480 13932
rect 11520 13923 11572 13932
rect 11520 13889 11529 13923
rect 11529 13889 11563 13923
rect 11563 13889 11572 13923
rect 11520 13880 11572 13889
rect 11152 13812 11204 13864
rect 11612 13855 11664 13864
rect 11612 13821 11621 13855
rect 11621 13821 11655 13855
rect 11655 13821 11664 13855
rect 11612 13812 11664 13821
rect 11704 13812 11756 13864
rect 8208 13744 8260 13796
rect 9772 13744 9824 13796
rect 10324 13744 10376 13796
rect 10600 13787 10652 13796
rect 10600 13753 10609 13787
rect 10609 13753 10643 13787
rect 10643 13753 10652 13787
rect 10600 13744 10652 13753
rect 2872 13676 2924 13728
rect 3240 13676 3292 13728
rect 4160 13676 4212 13728
rect 5172 13676 5224 13728
rect 5356 13676 5408 13728
rect 8852 13719 8904 13728
rect 8852 13685 8861 13719
rect 8861 13685 8895 13719
rect 8895 13685 8904 13719
rect 8852 13676 8904 13685
rect 9956 13719 10008 13728
rect 9956 13685 9965 13719
rect 9965 13685 9999 13719
rect 9999 13685 10008 13719
rect 9956 13676 10008 13685
rect 10416 13676 10468 13728
rect 11152 13676 11204 13728
rect 12348 13719 12400 13728
rect 12348 13685 12357 13719
rect 12357 13685 12391 13719
rect 12391 13685 12400 13719
rect 12348 13676 12400 13685
rect 18420 13880 18472 13932
rect 18512 13923 18564 13932
rect 18512 13889 18521 13923
rect 18521 13889 18555 13923
rect 18555 13889 18564 13923
rect 19524 13948 19576 14000
rect 19892 13991 19944 14000
rect 19892 13957 19901 13991
rect 19901 13957 19935 13991
rect 19935 13957 19944 13991
rect 19892 13948 19944 13957
rect 21548 13948 21600 14000
rect 18512 13880 18564 13889
rect 14740 13744 14792 13796
rect 16396 13812 16448 13864
rect 16672 13855 16724 13864
rect 16672 13821 16681 13855
rect 16681 13821 16715 13855
rect 16715 13821 16724 13855
rect 16672 13812 16724 13821
rect 15292 13676 15344 13728
rect 15844 13676 15896 13728
rect 17868 13744 17920 13796
rect 17776 13676 17828 13728
rect 17960 13676 18012 13728
rect 18880 13923 18932 13932
rect 18880 13889 18889 13923
rect 18889 13889 18923 13923
rect 18923 13889 18932 13923
rect 18880 13880 18932 13889
rect 19064 13880 19116 13932
rect 19616 13880 19668 13932
rect 19156 13812 19208 13864
rect 20352 13744 20404 13796
rect 20628 13744 20680 13796
rect 21180 13880 21232 13932
rect 21824 13923 21876 13932
rect 21824 13889 21833 13923
rect 21833 13889 21867 13923
rect 21867 13889 21876 13923
rect 21824 13880 21876 13889
rect 21916 13812 21968 13864
rect 22652 13880 22704 13932
rect 23112 13923 23164 13932
rect 23112 13889 23121 13923
rect 23121 13889 23155 13923
rect 23155 13889 23164 13923
rect 23112 13880 23164 13889
rect 23204 13880 23256 13932
rect 25136 14016 25188 14068
rect 26792 14016 26844 14068
rect 24216 13948 24268 14000
rect 24860 13948 24912 14000
rect 25688 13948 25740 14000
rect 24676 13880 24728 13932
rect 25136 13923 25188 13932
rect 25136 13889 25145 13923
rect 25145 13889 25179 13923
rect 25179 13889 25188 13923
rect 25136 13880 25188 13889
rect 25504 13923 25556 13932
rect 25504 13889 25513 13923
rect 25513 13889 25547 13923
rect 25547 13889 25556 13923
rect 25504 13880 25556 13889
rect 26516 13880 26568 13932
rect 22192 13812 22244 13864
rect 23480 13812 23532 13864
rect 21548 13744 21600 13796
rect 21732 13744 21784 13796
rect 23112 13744 23164 13796
rect 24216 13812 24268 13864
rect 25136 13744 25188 13796
rect 25412 13812 25464 13864
rect 25872 13812 25924 13864
rect 26056 13812 26108 13864
rect 19524 13676 19576 13728
rect 20720 13676 20772 13728
rect 22100 13676 22152 13728
rect 26884 13744 26936 13796
rect 26148 13676 26200 13728
rect 5442 13574 5494 13626
rect 5506 13574 5558 13626
rect 5570 13574 5622 13626
rect 5634 13574 5686 13626
rect 5698 13574 5750 13626
rect 14428 13574 14480 13626
rect 14492 13574 14544 13626
rect 14556 13574 14608 13626
rect 14620 13574 14672 13626
rect 14684 13574 14736 13626
rect 23413 13574 23465 13626
rect 23477 13574 23529 13626
rect 23541 13574 23593 13626
rect 23605 13574 23657 13626
rect 23669 13574 23721 13626
rect 5356 13472 5408 13524
rect 3884 13404 3936 13456
rect 8484 13472 8536 13524
rect 10692 13515 10744 13524
rect 4344 13336 4396 13388
rect 5172 13336 5224 13388
rect 1676 13268 1728 13320
rect 8668 13404 8720 13456
rect 10692 13481 10701 13515
rect 10701 13481 10735 13515
rect 10735 13481 10744 13515
rect 10692 13472 10744 13481
rect 14096 13472 14148 13524
rect 15016 13472 15068 13524
rect 16580 13472 16632 13524
rect 17592 13515 17644 13524
rect 17592 13481 17601 13515
rect 17601 13481 17635 13515
rect 17635 13481 17644 13515
rect 17592 13472 17644 13481
rect 11060 13404 11112 13456
rect 11520 13404 11572 13456
rect 18788 13472 18840 13524
rect 19064 13472 19116 13524
rect 20352 13472 20404 13524
rect 20904 13472 20956 13524
rect 21732 13472 21784 13524
rect 22192 13472 22244 13524
rect 23020 13472 23072 13524
rect 26240 13472 26292 13524
rect 26884 13472 26936 13524
rect 7012 13268 7064 13320
rect 2504 13200 2556 13252
rect 4620 13200 4672 13252
rect 5448 13243 5500 13252
rect 4068 13132 4120 13184
rect 5448 13209 5457 13243
rect 5457 13209 5491 13243
rect 5491 13209 5500 13243
rect 5448 13200 5500 13209
rect 7932 13132 7984 13184
rect 8484 13268 8536 13320
rect 10508 13336 10560 13388
rect 11336 13379 11388 13388
rect 11336 13345 11345 13379
rect 11345 13345 11379 13379
rect 11379 13345 11388 13379
rect 11336 13336 11388 13345
rect 15936 13336 15988 13388
rect 22100 13404 22152 13456
rect 23480 13404 23532 13456
rect 9680 13268 9732 13320
rect 12348 13268 12400 13320
rect 13544 13268 13596 13320
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 15384 13268 15436 13320
rect 15660 13311 15712 13320
rect 15660 13277 15670 13311
rect 15670 13277 15704 13311
rect 15704 13277 15712 13311
rect 15660 13268 15712 13277
rect 16948 13311 17000 13320
rect 16948 13277 16957 13311
rect 16957 13277 16991 13311
rect 16991 13277 17000 13311
rect 16948 13268 17000 13277
rect 17132 13311 17184 13320
rect 17132 13277 17139 13311
rect 17139 13277 17184 13311
rect 17132 13268 17184 13277
rect 17776 13268 17828 13320
rect 19892 13336 19944 13388
rect 20720 13336 20772 13388
rect 23572 13336 23624 13388
rect 25412 13336 25464 13388
rect 9036 13200 9088 13252
rect 15844 13243 15896 13252
rect 15844 13209 15853 13243
rect 15853 13209 15887 13243
rect 15887 13209 15896 13243
rect 15844 13200 15896 13209
rect 15936 13243 15988 13252
rect 15936 13209 15945 13243
rect 15945 13209 15979 13243
rect 15979 13209 15988 13243
rect 15936 13200 15988 13209
rect 9772 13132 9824 13184
rect 10784 13132 10836 13184
rect 14096 13132 14148 13184
rect 17960 13200 18012 13252
rect 17868 13132 17920 13184
rect 18052 13132 18104 13184
rect 18788 13268 18840 13320
rect 19156 13200 19208 13252
rect 18420 13132 18472 13184
rect 18512 13132 18564 13184
rect 19524 13243 19576 13252
rect 19524 13209 19533 13243
rect 19533 13209 19567 13243
rect 19567 13209 19576 13243
rect 19524 13200 19576 13209
rect 19616 13277 19633 13298
rect 19633 13277 19667 13298
rect 19667 13277 19668 13298
rect 19616 13246 19668 13277
rect 20076 13268 20128 13320
rect 20628 13311 20680 13320
rect 20628 13277 20637 13311
rect 20637 13277 20671 13311
rect 20671 13277 20680 13311
rect 20628 13268 20680 13277
rect 21824 13268 21876 13320
rect 21916 13268 21968 13320
rect 23756 13268 23808 13320
rect 24676 13268 24728 13320
rect 24952 13311 25004 13320
rect 24952 13277 24961 13311
rect 24961 13277 24995 13311
rect 24995 13277 25004 13311
rect 24952 13268 25004 13277
rect 25596 13268 25648 13320
rect 25964 13311 26016 13320
rect 25964 13277 25973 13311
rect 25973 13277 26007 13311
rect 26007 13277 26016 13311
rect 25964 13268 26016 13277
rect 21180 13200 21232 13252
rect 23296 13200 23348 13252
rect 26424 13200 26476 13252
rect 20076 13132 20128 13184
rect 20720 13132 20772 13184
rect 22100 13132 22152 13184
rect 22284 13132 22336 13184
rect 24032 13132 24084 13184
rect 25412 13132 25464 13184
rect 9935 13030 9987 13082
rect 9999 13030 10051 13082
rect 10063 13030 10115 13082
rect 10127 13030 10179 13082
rect 10191 13030 10243 13082
rect 18920 13030 18972 13082
rect 18984 13030 19036 13082
rect 19048 13030 19100 13082
rect 19112 13030 19164 13082
rect 19176 13030 19228 13082
rect 4252 12928 4304 12980
rect 4620 12928 4672 12980
rect 3608 12860 3660 12912
rect 2044 12792 2096 12844
rect 4344 12860 4396 12912
rect 4712 12860 4764 12912
rect 4896 12860 4948 12912
rect 5540 12860 5592 12912
rect 6368 12860 6420 12912
rect 6920 12860 6972 12912
rect 5080 12792 5132 12844
rect 7012 12792 7064 12844
rect 3424 12724 3476 12776
rect 6368 12724 6420 12776
rect 5080 12656 5132 12708
rect 5448 12656 5500 12708
rect 7472 12928 7524 12980
rect 8484 12928 8536 12980
rect 9312 12860 9364 12912
rect 10324 12928 10376 12980
rect 11152 12928 11204 12980
rect 14004 12928 14056 12980
rect 16672 12928 16724 12980
rect 10784 12860 10836 12912
rect 10968 12860 11020 12912
rect 7932 12835 7984 12844
rect 7932 12801 7941 12835
rect 7941 12801 7975 12835
rect 7975 12801 7984 12835
rect 7932 12792 7984 12801
rect 8392 12792 8444 12844
rect 9128 12792 9180 12844
rect 9220 12792 9272 12844
rect 8852 12767 8904 12776
rect 8852 12733 8861 12767
rect 8861 12733 8895 12767
rect 8895 12733 8904 12767
rect 8852 12724 8904 12733
rect 2688 12588 2740 12640
rect 4160 12588 4212 12640
rect 4344 12588 4396 12640
rect 6644 12588 6696 12640
rect 6828 12588 6880 12640
rect 7380 12588 7432 12640
rect 7840 12588 7892 12640
rect 8024 12588 8076 12640
rect 8392 12588 8444 12640
rect 8668 12588 8720 12640
rect 9772 12792 9824 12844
rect 10048 12835 10100 12844
rect 10048 12801 10057 12835
rect 10057 12801 10091 12835
rect 10091 12801 10100 12835
rect 10048 12792 10100 12801
rect 14280 12860 14332 12912
rect 16028 12860 16080 12912
rect 16396 12860 16448 12912
rect 17868 12928 17920 12980
rect 18420 12928 18472 12980
rect 19524 12928 19576 12980
rect 19616 12928 19668 12980
rect 20076 12928 20128 12980
rect 21364 12928 21416 12980
rect 21824 12928 21876 12980
rect 22008 12928 22060 12980
rect 22376 12928 22428 12980
rect 24676 12928 24728 12980
rect 18144 12860 18196 12912
rect 18328 12860 18380 12912
rect 23480 12860 23532 12912
rect 11520 12835 11572 12844
rect 11520 12801 11529 12835
rect 11529 12801 11563 12835
rect 11563 12801 11572 12835
rect 11520 12792 11572 12801
rect 12256 12835 12308 12844
rect 12256 12801 12265 12835
rect 12265 12801 12299 12835
rect 12299 12801 12308 12835
rect 12256 12792 12308 12801
rect 13268 12835 13320 12844
rect 9496 12656 9548 12708
rect 10600 12724 10652 12776
rect 12164 12724 12216 12776
rect 13268 12801 13277 12835
rect 13277 12801 13311 12835
rect 13311 12801 13320 12835
rect 13268 12792 13320 12801
rect 14832 12792 14884 12844
rect 13544 12767 13596 12776
rect 13544 12733 13553 12767
rect 13553 12733 13587 12767
rect 13587 12733 13596 12767
rect 16580 12792 16632 12844
rect 17132 12835 17184 12844
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 13544 12724 13596 12733
rect 15660 12724 15712 12776
rect 18420 12792 18472 12844
rect 19064 12792 19116 12844
rect 20352 12792 20404 12844
rect 20720 12835 20772 12844
rect 20720 12801 20729 12835
rect 20729 12801 20763 12835
rect 20763 12801 20772 12835
rect 20720 12792 20772 12801
rect 20904 12835 20956 12844
rect 20904 12801 20913 12835
rect 20913 12801 20947 12835
rect 20947 12801 20956 12835
rect 20904 12792 20956 12801
rect 14372 12699 14424 12708
rect 14372 12665 14381 12699
rect 14381 12665 14415 12699
rect 14415 12665 14424 12699
rect 14372 12656 14424 12665
rect 15200 12656 15252 12708
rect 17316 12656 17368 12708
rect 12348 12631 12400 12640
rect 12348 12597 12357 12631
rect 12357 12597 12391 12631
rect 12391 12597 12400 12631
rect 12348 12588 12400 12597
rect 12808 12588 12860 12640
rect 16028 12588 16080 12640
rect 16212 12588 16264 12640
rect 16856 12588 16908 12640
rect 21180 12792 21232 12844
rect 21548 12724 21600 12776
rect 22284 12792 22336 12844
rect 22652 12792 22704 12844
rect 23756 12860 23808 12912
rect 25964 12860 26016 12912
rect 23940 12835 23992 12844
rect 23940 12801 23974 12835
rect 23974 12801 23992 12835
rect 23940 12792 23992 12801
rect 24860 12792 24912 12844
rect 25780 12792 25832 12844
rect 26148 12835 26200 12844
rect 26148 12801 26157 12835
rect 26157 12801 26191 12835
rect 26191 12801 26200 12835
rect 26148 12792 26200 12801
rect 22928 12767 22980 12776
rect 22928 12733 22937 12767
rect 22937 12733 22971 12767
rect 22971 12733 22980 12767
rect 22928 12724 22980 12733
rect 23388 12724 23440 12776
rect 24768 12724 24820 12776
rect 26608 12724 26660 12776
rect 21732 12656 21784 12708
rect 23572 12656 23624 12708
rect 26240 12656 26292 12708
rect 19892 12588 19944 12640
rect 19984 12588 20036 12640
rect 20352 12588 20404 12640
rect 21364 12588 21416 12640
rect 21640 12588 21692 12640
rect 22100 12588 22152 12640
rect 26332 12631 26384 12640
rect 26332 12597 26341 12631
rect 26341 12597 26375 12631
rect 26375 12597 26384 12631
rect 26332 12588 26384 12597
rect 27068 12588 27120 12640
rect 27528 12588 27580 12640
rect 28080 12588 28132 12640
rect 5442 12486 5494 12538
rect 5506 12486 5558 12538
rect 5570 12486 5622 12538
rect 5634 12486 5686 12538
rect 5698 12486 5750 12538
rect 14428 12486 14480 12538
rect 14492 12486 14544 12538
rect 14556 12486 14608 12538
rect 14620 12486 14672 12538
rect 14684 12486 14736 12538
rect 23413 12486 23465 12538
rect 23477 12486 23529 12538
rect 23541 12486 23593 12538
rect 23605 12486 23657 12538
rect 23669 12486 23721 12538
rect 1860 12384 1912 12436
rect 2504 12427 2556 12436
rect 2504 12393 2513 12427
rect 2513 12393 2547 12427
rect 2547 12393 2556 12427
rect 2504 12384 2556 12393
rect 3424 12384 3476 12436
rect 2964 12316 3016 12368
rect 3976 12384 4028 12436
rect 4344 12384 4396 12436
rect 4528 12384 4580 12436
rect 7748 12427 7800 12436
rect 7748 12393 7757 12427
rect 7757 12393 7791 12427
rect 7791 12393 7800 12427
rect 7748 12384 7800 12393
rect 10048 12384 10100 12436
rect 2136 12248 2188 12300
rect 2504 12248 2556 12300
rect 2688 12223 2740 12232
rect 2688 12189 2697 12223
rect 2697 12189 2731 12223
rect 2731 12189 2740 12223
rect 2688 12180 2740 12189
rect 3424 12180 3476 12232
rect 4068 12223 4120 12232
rect 4068 12189 4077 12223
rect 4077 12189 4111 12223
rect 4111 12189 4120 12223
rect 4068 12180 4120 12189
rect 1676 12155 1728 12164
rect 1676 12121 1685 12155
rect 1685 12121 1719 12155
rect 1719 12121 1728 12155
rect 1676 12112 1728 12121
rect 2136 12112 2188 12164
rect 3976 12044 4028 12096
rect 5724 12316 5776 12368
rect 6000 12316 6052 12368
rect 6828 12316 6880 12368
rect 8024 12316 8076 12368
rect 4988 12248 5040 12300
rect 4712 12180 4764 12232
rect 5356 12223 5408 12232
rect 5356 12189 5365 12223
rect 5365 12189 5399 12223
rect 5399 12189 5408 12223
rect 5356 12180 5408 12189
rect 6000 12180 6052 12232
rect 6368 12223 6420 12232
rect 6368 12189 6377 12223
rect 6377 12189 6411 12223
rect 6411 12189 6420 12223
rect 6368 12180 6420 12189
rect 6644 12223 6696 12232
rect 6644 12189 6653 12223
rect 6653 12189 6687 12223
rect 6687 12189 6696 12223
rect 6644 12180 6696 12189
rect 8944 12316 8996 12368
rect 9772 12316 9824 12368
rect 12992 12384 13044 12436
rect 13268 12384 13320 12436
rect 10600 12248 10652 12300
rect 11704 12291 11756 12300
rect 11704 12257 11713 12291
rect 11713 12257 11747 12291
rect 11747 12257 11756 12291
rect 11704 12248 11756 12257
rect 13268 12248 13320 12300
rect 13452 12248 13504 12300
rect 5540 12155 5592 12164
rect 5540 12121 5549 12155
rect 5549 12121 5583 12155
rect 5583 12121 5592 12155
rect 5540 12112 5592 12121
rect 10324 12180 10376 12232
rect 10508 12223 10560 12232
rect 10508 12189 10517 12223
rect 10517 12189 10551 12223
rect 10551 12189 10560 12223
rect 10508 12180 10560 12189
rect 5908 12087 5960 12096
rect 5908 12053 5917 12087
rect 5917 12053 5951 12087
rect 5951 12053 5960 12087
rect 5908 12044 5960 12053
rect 8300 12112 8352 12164
rect 8852 12112 8904 12164
rect 9588 12112 9640 12164
rect 11612 12112 11664 12164
rect 15936 12384 15988 12436
rect 18052 12384 18104 12436
rect 21548 12427 21600 12436
rect 20076 12316 20128 12368
rect 21548 12393 21557 12427
rect 21557 12393 21591 12427
rect 21591 12393 21600 12427
rect 21548 12384 21600 12393
rect 23296 12427 23348 12436
rect 23296 12393 23305 12427
rect 23305 12393 23339 12427
rect 23339 12393 23348 12427
rect 23296 12384 23348 12393
rect 22284 12316 22336 12368
rect 22928 12316 22980 12368
rect 24124 12316 24176 12368
rect 26332 12384 26384 12436
rect 27620 12384 27672 12436
rect 27896 12384 27948 12436
rect 18052 12248 18104 12300
rect 19064 12248 19116 12300
rect 19708 12291 19760 12300
rect 19708 12257 19717 12291
rect 19717 12257 19751 12291
rect 19751 12257 19760 12291
rect 19708 12248 19760 12257
rect 21180 12248 21232 12300
rect 24032 12248 24084 12300
rect 25504 12291 25556 12300
rect 25504 12257 25513 12291
rect 25513 12257 25547 12291
rect 25547 12257 25556 12291
rect 25504 12248 25556 12257
rect 25964 12291 26016 12300
rect 25964 12257 25973 12291
rect 25973 12257 26007 12291
rect 26007 12257 26016 12291
rect 25964 12248 26016 12257
rect 27436 12248 27488 12300
rect 27620 12248 27672 12300
rect 15936 12112 15988 12164
rect 16672 12112 16724 12164
rect 17776 12112 17828 12164
rect 21916 12180 21968 12232
rect 22284 12223 22336 12232
rect 18604 12112 18656 12164
rect 19156 12112 19208 12164
rect 20076 12112 20128 12164
rect 20536 12112 20588 12164
rect 20628 12112 20680 12164
rect 8024 12044 8076 12096
rect 8392 12044 8444 12096
rect 11888 12044 11940 12096
rect 12532 12044 12584 12096
rect 12808 12044 12860 12096
rect 12900 12044 12952 12096
rect 13728 12044 13780 12096
rect 13820 12044 13872 12096
rect 15844 12044 15896 12096
rect 16212 12044 16264 12096
rect 17684 12044 17736 12096
rect 22284 12189 22293 12223
rect 22293 12189 22327 12223
rect 22327 12189 22336 12223
rect 22284 12180 22336 12189
rect 23848 12180 23900 12232
rect 24400 12180 24452 12232
rect 25044 12180 25096 12232
rect 25412 12180 25464 12232
rect 26240 12223 26292 12232
rect 26240 12189 26274 12223
rect 26274 12189 26292 12223
rect 26240 12180 26292 12189
rect 26608 12112 26660 12164
rect 23112 12044 23164 12096
rect 24032 12044 24084 12096
rect 25136 12044 25188 12096
rect 27436 12044 27488 12096
rect 28080 12044 28132 12096
rect 9935 11942 9987 11994
rect 9999 11942 10051 11994
rect 10063 11942 10115 11994
rect 10127 11942 10179 11994
rect 10191 11942 10243 11994
rect 18920 11942 18972 11994
rect 18984 11942 19036 11994
rect 19048 11942 19100 11994
rect 19112 11942 19164 11994
rect 19176 11942 19228 11994
rect 1676 11840 1728 11892
rect 3608 11840 3660 11892
rect 5264 11840 5316 11892
rect 6276 11840 6328 11892
rect 7012 11840 7064 11892
rect 2412 11772 2464 11824
rect 1032 11704 1084 11756
rect 1676 11704 1728 11756
rect 2044 11747 2096 11756
rect 2044 11713 2053 11747
rect 2053 11713 2087 11747
rect 2087 11713 2096 11747
rect 2044 11704 2096 11713
rect 2780 11704 2832 11756
rect 3424 11704 3476 11756
rect 4436 11772 4488 11824
rect 6368 11772 6420 11824
rect 4344 11747 4396 11756
rect 4344 11713 4353 11747
rect 4353 11713 4387 11747
rect 4387 11713 4396 11747
rect 4344 11704 4396 11713
rect 5080 11747 5132 11756
rect 5080 11713 5089 11747
rect 5089 11713 5123 11747
rect 5123 11713 5132 11747
rect 5080 11704 5132 11713
rect 3884 11636 3936 11688
rect 4436 11636 4488 11688
rect 4804 11636 4856 11688
rect 5356 11636 5408 11688
rect 5908 11704 5960 11756
rect 7656 11772 7708 11824
rect 9036 11840 9088 11892
rect 9588 11840 9640 11892
rect 10324 11840 10376 11892
rect 11980 11840 12032 11892
rect 14464 11883 14516 11892
rect 14464 11849 14489 11883
rect 14489 11849 14516 11883
rect 14648 11883 14700 11892
rect 14464 11840 14516 11849
rect 14648 11849 14657 11883
rect 14657 11849 14691 11883
rect 14691 11849 14700 11883
rect 14648 11840 14700 11849
rect 6000 11636 6052 11688
rect 3976 11568 4028 11620
rect 5724 11568 5776 11620
rect 1860 11543 1912 11552
rect 1860 11509 1869 11543
rect 1869 11509 1903 11543
rect 1903 11509 1912 11543
rect 1860 11500 1912 11509
rect 5908 11500 5960 11552
rect 6276 11500 6328 11552
rect 6644 11636 6696 11688
rect 9036 11704 9088 11756
rect 9404 11704 9456 11756
rect 12716 11747 12768 11756
rect 8392 11500 8444 11552
rect 11704 11500 11756 11552
rect 11888 11500 11940 11552
rect 12164 11500 12216 11552
rect 12716 11713 12725 11747
rect 12725 11713 12759 11747
rect 12759 11713 12768 11747
rect 12716 11704 12768 11713
rect 12992 11747 13044 11756
rect 12992 11713 13001 11747
rect 13001 11713 13035 11747
rect 13035 11713 13044 11747
rect 12992 11704 13044 11713
rect 13084 11704 13136 11756
rect 15936 11772 15988 11824
rect 13452 11636 13504 11688
rect 13084 11568 13136 11620
rect 13728 11611 13780 11620
rect 13728 11577 13737 11611
rect 13737 11577 13771 11611
rect 13771 11577 13780 11611
rect 13728 11568 13780 11577
rect 12532 11500 12584 11552
rect 12808 11500 12860 11552
rect 13820 11500 13872 11552
rect 14280 11500 14332 11552
rect 15200 11636 15252 11688
rect 17316 11840 17368 11892
rect 17500 11840 17552 11892
rect 18604 11883 18656 11892
rect 18604 11849 18613 11883
rect 18613 11849 18647 11883
rect 18647 11849 18656 11883
rect 18604 11840 18656 11849
rect 19432 11772 19484 11824
rect 19800 11840 19852 11892
rect 20076 11840 20128 11892
rect 20352 11840 20404 11892
rect 20996 11840 21048 11892
rect 22008 11840 22060 11892
rect 23296 11840 23348 11892
rect 23940 11840 23992 11892
rect 25504 11840 25556 11892
rect 26608 11840 26660 11892
rect 27344 11840 27396 11892
rect 17776 11704 17828 11756
rect 18880 11704 18932 11756
rect 19156 11704 19208 11756
rect 21180 11772 21232 11824
rect 15844 11568 15896 11620
rect 15292 11500 15344 11552
rect 19800 11636 19852 11688
rect 22008 11704 22060 11756
rect 19524 11568 19576 11620
rect 20260 11568 20312 11620
rect 20628 11568 20680 11620
rect 21180 11636 21232 11688
rect 21640 11636 21692 11688
rect 22284 11747 22336 11756
rect 22284 11713 22293 11747
rect 22293 11713 22327 11747
rect 22327 11713 22336 11747
rect 22284 11704 22336 11713
rect 23112 11704 23164 11756
rect 23756 11772 23808 11824
rect 24768 11772 24820 11824
rect 24216 11747 24268 11756
rect 24216 11713 24225 11747
rect 24225 11713 24259 11747
rect 24259 11713 24268 11747
rect 24216 11704 24268 11713
rect 25136 11704 25188 11756
rect 25596 11704 25648 11756
rect 26700 11704 26752 11756
rect 27068 11747 27120 11756
rect 27068 11713 27077 11747
rect 27077 11713 27111 11747
rect 27111 11713 27120 11747
rect 27068 11704 27120 11713
rect 24676 11636 24728 11688
rect 27252 11611 27304 11620
rect 27252 11577 27261 11611
rect 27261 11577 27295 11611
rect 27295 11577 27304 11611
rect 27252 11568 27304 11577
rect 20536 11500 20588 11552
rect 22284 11500 22336 11552
rect 22836 11500 22888 11552
rect 24216 11500 24268 11552
rect 24308 11500 24360 11552
rect 26332 11500 26384 11552
rect 5442 11398 5494 11450
rect 5506 11398 5558 11450
rect 5570 11398 5622 11450
rect 5634 11398 5686 11450
rect 5698 11398 5750 11450
rect 14428 11398 14480 11450
rect 14492 11398 14544 11450
rect 14556 11398 14608 11450
rect 14620 11398 14672 11450
rect 14684 11398 14736 11450
rect 23413 11398 23465 11450
rect 23477 11398 23529 11450
rect 23541 11398 23593 11450
rect 23605 11398 23657 11450
rect 23669 11398 23721 11450
rect 6460 11296 6512 11348
rect 9312 11339 9364 11348
rect 9312 11305 9321 11339
rect 9321 11305 9355 11339
rect 9355 11305 9364 11339
rect 9312 11296 9364 11305
rect 9404 11296 9456 11348
rect 2688 11228 2740 11280
rect 3884 11228 3936 11280
rect 6276 11228 6328 11280
rect 9864 11228 9916 11280
rect 10692 11296 10744 11348
rect 11428 11296 11480 11348
rect 12164 11296 12216 11348
rect 13728 11296 13780 11348
rect 13820 11296 13872 11348
rect 14096 11296 14148 11348
rect 15844 11296 15896 11348
rect 1860 11024 1912 11076
rect 3332 11092 3384 11144
rect 3516 11092 3568 11144
rect 6644 11160 6696 11212
rect 6920 11160 6972 11212
rect 16120 11228 16172 11280
rect 5908 11135 5960 11144
rect 3332 10956 3384 11008
rect 4252 11024 4304 11076
rect 5908 11101 5917 11135
rect 5917 11101 5951 11135
rect 5951 11101 5960 11135
rect 5908 11092 5960 11101
rect 6276 11092 6328 11144
rect 7012 11092 7064 11144
rect 7656 11092 7708 11144
rect 8852 11092 8904 11144
rect 8944 11092 8996 11144
rect 4344 10956 4396 11008
rect 4988 10956 5040 11008
rect 6460 11024 6512 11076
rect 5264 10999 5316 11008
rect 5264 10965 5273 10999
rect 5273 10965 5307 10999
rect 5307 10965 5316 10999
rect 5264 10956 5316 10965
rect 6828 10956 6880 11008
rect 7656 10956 7708 11008
rect 8116 10956 8168 11008
rect 8392 10956 8444 11008
rect 10508 11092 10560 11144
rect 10968 11160 11020 11212
rect 11428 11135 11480 11144
rect 11428 11101 11437 11135
rect 11437 11101 11471 11135
rect 11471 11101 11480 11135
rect 11428 11092 11480 11101
rect 13544 11160 13596 11212
rect 11888 11135 11940 11144
rect 11888 11101 11897 11135
rect 11897 11101 11931 11135
rect 11931 11101 11940 11135
rect 11888 11092 11940 11101
rect 12716 11135 12768 11144
rect 12716 11101 12725 11135
rect 12725 11101 12759 11135
rect 12759 11101 12768 11135
rect 12716 11092 12768 11101
rect 13452 11092 13504 11144
rect 13912 11092 13964 11144
rect 14280 11092 14332 11144
rect 16488 11135 16540 11144
rect 16488 11101 16497 11135
rect 16497 11101 16531 11135
rect 16531 11101 16540 11135
rect 16488 11092 16540 11101
rect 17224 11296 17276 11348
rect 18788 11296 18840 11348
rect 20444 11296 20496 11348
rect 21640 11339 21692 11348
rect 21640 11305 21649 11339
rect 21649 11305 21683 11339
rect 21683 11305 21692 11339
rect 21640 11296 21692 11305
rect 23204 11296 23256 11348
rect 16672 11228 16724 11280
rect 24216 11228 24268 11280
rect 9680 11024 9732 11076
rect 10692 11024 10744 11076
rect 12624 11024 12676 11076
rect 10968 10956 11020 11008
rect 12256 10956 12308 11008
rect 14188 10956 14240 11008
rect 14280 10956 14332 11008
rect 16396 11024 16448 11076
rect 21916 11160 21968 11212
rect 24308 11160 24360 11212
rect 25504 11160 25556 11212
rect 19708 11092 19760 11144
rect 20352 11092 20404 11144
rect 16488 10956 16540 11008
rect 19156 11024 19208 11076
rect 19432 11067 19484 11076
rect 19432 11033 19441 11067
rect 19441 11033 19475 11067
rect 19475 11033 19484 11067
rect 19432 11024 19484 11033
rect 19524 11024 19576 11076
rect 19800 11024 19852 11076
rect 22744 11092 22796 11144
rect 24400 11135 24452 11144
rect 24400 11101 24409 11135
rect 24409 11101 24443 11135
rect 24443 11101 24452 11135
rect 24400 11092 24452 11101
rect 26424 11296 26476 11348
rect 27252 11296 27304 11348
rect 27620 11296 27672 11348
rect 26332 11160 26384 11212
rect 26884 11160 26936 11212
rect 22468 11024 22520 11076
rect 23296 11024 23348 11076
rect 25044 11024 25096 11076
rect 18052 10956 18104 11008
rect 18236 10956 18288 11008
rect 20904 10956 20956 11008
rect 20996 10956 21048 11008
rect 21272 10956 21324 11008
rect 23848 10956 23900 11008
rect 24124 10956 24176 11008
rect 24492 10956 24544 11008
rect 26332 11024 26384 11076
rect 25596 10956 25648 11008
rect 9935 10854 9987 10906
rect 9999 10854 10051 10906
rect 10063 10854 10115 10906
rect 10127 10854 10179 10906
rect 10191 10854 10243 10906
rect 18920 10854 18972 10906
rect 18984 10854 19036 10906
rect 19048 10854 19100 10906
rect 19112 10854 19164 10906
rect 19176 10854 19228 10906
rect 2044 10752 2096 10804
rect 3884 10752 3936 10804
rect 2136 10616 2188 10668
rect 3424 10684 3476 10736
rect 3332 10659 3384 10668
rect 3332 10625 3341 10659
rect 3341 10625 3375 10659
rect 3375 10625 3384 10659
rect 4988 10684 5040 10736
rect 5540 10727 5592 10736
rect 5540 10693 5549 10727
rect 5549 10693 5583 10727
rect 5583 10693 5592 10727
rect 5540 10684 5592 10693
rect 5724 10752 5776 10804
rect 6552 10752 6604 10804
rect 7012 10752 7064 10804
rect 9220 10752 9272 10804
rect 10140 10684 10192 10736
rect 11796 10752 11848 10804
rect 12348 10752 12400 10804
rect 13912 10752 13964 10804
rect 15844 10752 15896 10804
rect 16396 10752 16448 10804
rect 17316 10752 17368 10804
rect 14372 10684 14424 10736
rect 3332 10616 3384 10625
rect 5264 10659 5316 10668
rect 2228 10548 2280 10600
rect 5264 10625 5273 10659
rect 5273 10625 5307 10659
rect 5307 10625 5316 10659
rect 5264 10616 5316 10625
rect 5356 10616 5408 10668
rect 6644 10616 6696 10668
rect 6828 10659 6880 10668
rect 6828 10625 6862 10659
rect 6862 10625 6880 10659
rect 6828 10616 6880 10625
rect 7380 10616 7432 10668
rect 7564 10616 7616 10668
rect 7656 10616 7708 10668
rect 8116 10616 8168 10668
rect 9956 10616 10008 10668
rect 1400 10412 1452 10464
rect 4988 10480 5040 10532
rect 6000 10548 6052 10600
rect 6552 10480 6604 10532
rect 8392 10591 8444 10600
rect 8392 10557 8401 10591
rect 8401 10557 8435 10591
rect 8435 10557 8444 10591
rect 8392 10548 8444 10557
rect 10324 10548 10376 10600
rect 3976 10412 4028 10464
rect 4804 10455 4856 10464
rect 4804 10421 4813 10455
rect 4813 10421 4847 10455
rect 4847 10421 4856 10455
rect 4804 10412 4856 10421
rect 7472 10412 7524 10464
rect 7564 10412 7616 10464
rect 10692 10616 10744 10668
rect 11152 10616 11204 10668
rect 11980 10616 12032 10668
rect 12348 10616 12400 10668
rect 12532 10616 12584 10668
rect 11704 10548 11756 10600
rect 13544 10616 13596 10668
rect 14096 10616 14148 10668
rect 15660 10659 15712 10668
rect 15660 10625 15669 10659
rect 15669 10625 15703 10659
rect 15703 10625 15712 10659
rect 15660 10616 15712 10625
rect 15844 10659 15896 10668
rect 15844 10625 15853 10659
rect 15853 10625 15887 10659
rect 15887 10625 15896 10659
rect 15844 10616 15896 10625
rect 16396 10616 16448 10668
rect 16672 10659 16724 10668
rect 15016 10548 15068 10600
rect 16672 10625 16681 10659
rect 16681 10625 16715 10659
rect 16715 10625 16724 10659
rect 16672 10616 16724 10625
rect 13084 10480 13136 10532
rect 15660 10480 15712 10532
rect 17868 10548 17920 10600
rect 18052 10523 18104 10532
rect 18052 10489 18061 10523
rect 18061 10489 18095 10523
rect 18095 10489 18104 10523
rect 18052 10480 18104 10489
rect 11060 10412 11112 10464
rect 11888 10455 11940 10464
rect 11888 10421 11897 10455
rect 11897 10421 11931 10455
rect 11931 10421 11940 10455
rect 11888 10412 11940 10421
rect 15292 10412 15344 10464
rect 19524 10616 19576 10668
rect 19708 10659 19760 10668
rect 19708 10625 19717 10659
rect 19717 10625 19751 10659
rect 19751 10625 19760 10659
rect 19708 10616 19760 10625
rect 20168 10684 20220 10736
rect 20720 10752 20772 10804
rect 21456 10752 21508 10804
rect 20904 10684 20956 10736
rect 22376 10752 22428 10804
rect 26332 10795 26384 10804
rect 21364 10616 21416 10668
rect 21916 10616 21968 10668
rect 22928 10616 22980 10668
rect 19156 10548 19208 10600
rect 24860 10684 24912 10736
rect 26332 10761 26341 10795
rect 26341 10761 26375 10795
rect 26375 10761 26384 10795
rect 26332 10752 26384 10761
rect 27804 10684 27856 10736
rect 23296 10616 23348 10668
rect 23848 10659 23900 10668
rect 23848 10625 23857 10659
rect 23857 10625 23891 10659
rect 23891 10625 23900 10659
rect 23848 10616 23900 10625
rect 24216 10659 24268 10668
rect 24216 10625 24225 10659
rect 24225 10625 24259 10659
rect 24259 10625 24268 10659
rect 24216 10616 24268 10625
rect 24768 10616 24820 10668
rect 25504 10616 25556 10668
rect 23940 10548 23992 10600
rect 20628 10412 20680 10464
rect 22836 10412 22888 10464
rect 26332 10412 26384 10464
rect 5442 10310 5494 10362
rect 5506 10310 5558 10362
rect 5570 10310 5622 10362
rect 5634 10310 5686 10362
rect 5698 10310 5750 10362
rect 14428 10310 14480 10362
rect 14492 10310 14544 10362
rect 14556 10310 14608 10362
rect 14620 10310 14672 10362
rect 14684 10310 14736 10362
rect 23413 10310 23465 10362
rect 23477 10310 23529 10362
rect 23541 10310 23593 10362
rect 23605 10310 23657 10362
rect 23669 10310 23721 10362
rect 2596 10208 2648 10260
rect 2872 10208 2924 10260
rect 3332 10208 3384 10260
rect 4344 10140 4396 10192
rect 6920 10208 6972 10260
rect 8116 10251 8168 10260
rect 8116 10217 8125 10251
rect 8125 10217 8159 10251
rect 8159 10217 8168 10251
rect 8116 10208 8168 10217
rect 2872 10004 2924 10056
rect 4804 10004 4856 10056
rect 5264 10004 5316 10056
rect 5540 10047 5592 10056
rect 5540 10013 5549 10047
rect 5549 10013 5583 10047
rect 5583 10013 5592 10047
rect 5540 10004 5592 10013
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 2228 9911 2280 9920
rect 2228 9877 2237 9911
rect 2237 9877 2271 9911
rect 2271 9877 2280 9911
rect 2228 9868 2280 9877
rect 3424 9868 3476 9920
rect 4252 9936 4304 9988
rect 4988 9936 5040 9988
rect 5724 9979 5776 9988
rect 5724 9945 5733 9979
rect 5733 9945 5767 9979
rect 5767 9945 5776 9979
rect 5724 9936 5776 9945
rect 4344 9868 4396 9920
rect 5356 9868 5408 9920
rect 6460 10004 6512 10056
rect 6920 10072 6972 10124
rect 8116 10072 8168 10124
rect 11796 10208 11848 10260
rect 11980 10208 12032 10260
rect 14096 10251 14148 10260
rect 10140 10115 10192 10124
rect 7564 10047 7616 10056
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 8300 10004 8352 10056
rect 9220 10047 9272 10056
rect 9220 10013 9229 10047
rect 9229 10013 9263 10047
rect 9263 10013 9272 10047
rect 9220 10004 9272 10013
rect 10140 10081 10149 10115
rect 10149 10081 10183 10115
rect 10183 10081 10192 10115
rect 10140 10072 10192 10081
rect 12164 10072 12216 10124
rect 14096 10217 14105 10251
rect 14105 10217 14139 10251
rect 14139 10217 14148 10251
rect 14096 10208 14148 10217
rect 14188 10208 14240 10260
rect 16396 10251 16448 10260
rect 12716 10140 12768 10192
rect 16396 10217 16405 10251
rect 16405 10217 16439 10251
rect 16439 10217 16448 10251
rect 16396 10208 16448 10217
rect 18236 10208 18288 10260
rect 18420 10208 18472 10260
rect 19524 10208 19576 10260
rect 20444 10208 20496 10260
rect 22468 10208 22520 10260
rect 22928 10208 22980 10260
rect 9680 10004 9732 10056
rect 10968 10004 11020 10056
rect 11336 10004 11388 10056
rect 14648 10072 14700 10124
rect 15016 10115 15068 10124
rect 15016 10081 15025 10115
rect 15025 10081 15059 10115
rect 15059 10081 15068 10115
rect 15016 10072 15068 10081
rect 16120 10072 16172 10124
rect 23664 10140 23716 10192
rect 24768 10140 24820 10192
rect 14280 10004 14332 10056
rect 15292 10047 15344 10056
rect 15292 10013 15326 10047
rect 15326 10013 15344 10047
rect 15292 10004 15344 10013
rect 16488 10004 16540 10056
rect 6552 9868 6604 9920
rect 7012 9868 7064 9920
rect 7564 9868 7616 9920
rect 7840 9979 7892 9988
rect 7840 9945 7849 9979
rect 7849 9945 7883 9979
rect 7883 9945 7892 9979
rect 7840 9936 7892 9945
rect 8484 9868 8536 9920
rect 9496 9868 9548 9920
rect 10968 9868 11020 9920
rect 11888 9868 11940 9920
rect 12256 9936 12308 9988
rect 12532 9868 12584 9920
rect 13084 9936 13136 9988
rect 13912 9868 13964 9920
rect 14188 9868 14240 9920
rect 15660 9936 15712 9988
rect 17316 10004 17368 10056
rect 17592 10004 17644 10056
rect 17684 10004 17736 10056
rect 17868 10047 17920 10056
rect 17868 10013 17877 10047
rect 17877 10013 17911 10047
rect 17911 10013 17920 10047
rect 17868 10004 17920 10013
rect 18604 9936 18656 9988
rect 19340 10004 19392 10056
rect 20904 10004 20956 10056
rect 19432 9979 19484 9988
rect 16396 9868 16448 9920
rect 17592 9868 17644 9920
rect 19432 9945 19441 9979
rect 19441 9945 19475 9979
rect 19475 9945 19484 9979
rect 19432 9936 19484 9945
rect 20996 9936 21048 9988
rect 20720 9868 20772 9920
rect 23112 10004 23164 10056
rect 22744 9979 22796 9988
rect 22744 9945 22753 9979
rect 22753 9945 22787 9979
rect 22787 9945 22796 9979
rect 22744 9936 22796 9945
rect 22652 9868 22704 9920
rect 23296 9868 23348 9920
rect 24216 10004 24268 10056
rect 24676 10004 24728 10056
rect 26700 9936 26752 9988
rect 25780 9868 25832 9920
rect 26884 9868 26936 9920
rect 9935 9766 9987 9818
rect 9999 9766 10051 9818
rect 10063 9766 10115 9818
rect 10127 9766 10179 9818
rect 10191 9766 10243 9818
rect 18920 9766 18972 9818
rect 18984 9766 19036 9818
rect 19048 9766 19100 9818
rect 19112 9766 19164 9818
rect 19176 9766 19228 9818
rect 1584 9664 1636 9716
rect 8116 9664 8168 9716
rect 9036 9664 9088 9716
rect 9496 9664 9548 9716
rect 2228 9596 2280 9648
rect 4344 9596 4396 9648
rect 3332 9528 3384 9580
rect 1584 9460 1636 9512
rect 3792 9460 3844 9512
rect 5540 9392 5592 9444
rect 5724 9596 5776 9648
rect 6644 9596 6696 9648
rect 7564 9596 7616 9648
rect 10968 9596 11020 9648
rect 11888 9664 11940 9716
rect 11796 9596 11848 9648
rect 6552 9528 6604 9580
rect 7840 9528 7892 9580
rect 8484 9528 8536 9580
rect 9404 9528 9456 9580
rect 9496 9528 9548 9580
rect 9864 9528 9916 9580
rect 8300 9503 8352 9512
rect 8300 9469 8309 9503
rect 8309 9469 8343 9503
rect 8343 9469 8352 9503
rect 11060 9528 11112 9580
rect 8300 9460 8352 9469
rect 12164 9460 12216 9512
rect 17040 9664 17092 9716
rect 17684 9664 17736 9716
rect 17776 9664 17828 9716
rect 16672 9596 16724 9648
rect 19524 9664 19576 9716
rect 13176 9503 13228 9512
rect 13176 9469 13185 9503
rect 13185 9469 13219 9503
rect 13219 9469 13228 9503
rect 13176 9460 13228 9469
rect 14648 9528 14700 9580
rect 15844 9571 15896 9580
rect 15844 9537 15853 9571
rect 15853 9537 15887 9571
rect 15887 9537 15896 9571
rect 15844 9528 15896 9537
rect 17040 9528 17092 9580
rect 18236 9528 18288 9580
rect 2964 9324 3016 9376
rect 4252 9324 4304 9376
rect 5816 9324 5868 9376
rect 8392 9392 8444 9444
rect 9036 9324 9088 9376
rect 10232 9392 10284 9444
rect 10508 9392 10560 9444
rect 9956 9324 10008 9376
rect 12256 9392 12308 9444
rect 11152 9324 11204 9376
rect 12532 9392 12584 9444
rect 16672 9460 16724 9512
rect 16948 9460 17000 9512
rect 12900 9324 12952 9376
rect 14832 9324 14884 9376
rect 17776 9392 17828 9444
rect 16948 9324 17000 9376
rect 18052 9324 18104 9376
rect 19340 9596 19392 9648
rect 23296 9664 23348 9716
rect 25228 9596 25280 9648
rect 19524 9528 19576 9580
rect 19800 9571 19852 9580
rect 19800 9537 19809 9571
rect 19809 9537 19843 9571
rect 19843 9537 19852 9571
rect 19800 9528 19852 9537
rect 19892 9528 19944 9580
rect 20720 9528 20772 9580
rect 21272 9571 21324 9580
rect 21272 9537 21281 9571
rect 21281 9537 21315 9571
rect 21315 9537 21324 9571
rect 21272 9528 21324 9537
rect 22100 9571 22152 9580
rect 22100 9537 22134 9571
rect 22134 9537 22152 9571
rect 23664 9571 23716 9580
rect 22100 9528 22152 9537
rect 23664 9537 23673 9571
rect 23673 9537 23707 9571
rect 23707 9537 23716 9571
rect 23664 9528 23716 9537
rect 27344 9664 27396 9716
rect 26424 9596 26476 9648
rect 20812 9460 20864 9512
rect 19708 9324 19760 9376
rect 20444 9367 20496 9376
rect 20444 9333 20453 9367
rect 20453 9333 20487 9367
rect 20487 9333 20496 9367
rect 20444 9324 20496 9333
rect 21364 9324 21416 9376
rect 23664 9392 23716 9444
rect 24860 9392 24912 9444
rect 25320 9392 25372 9444
rect 25780 9528 25832 9580
rect 26056 9528 26108 9580
rect 27160 9460 27212 9512
rect 27068 9392 27120 9444
rect 23848 9324 23900 9376
rect 25504 9367 25556 9376
rect 25504 9333 25513 9367
rect 25513 9333 25547 9367
rect 25547 9333 25556 9367
rect 25504 9324 25556 9333
rect 27620 9324 27672 9376
rect 5442 9222 5494 9274
rect 5506 9222 5558 9274
rect 5570 9222 5622 9274
rect 5634 9222 5686 9274
rect 5698 9222 5750 9274
rect 14428 9222 14480 9274
rect 14492 9222 14544 9274
rect 14556 9222 14608 9274
rect 14620 9222 14672 9274
rect 14684 9222 14736 9274
rect 23413 9222 23465 9274
rect 23477 9222 23529 9274
rect 23541 9222 23593 9274
rect 23605 9222 23657 9274
rect 23669 9222 23721 9274
rect 9956 9120 10008 9172
rect 2596 8984 2648 9036
rect 2688 8984 2740 9036
rect 3976 9052 4028 9104
rect 7564 9052 7616 9104
rect 1768 8916 1820 8968
rect 2964 8959 3016 8968
rect 2964 8925 2973 8959
rect 2973 8925 3007 8959
rect 3007 8925 3016 8959
rect 2964 8916 3016 8925
rect 2320 8848 2372 8900
rect 2596 8780 2648 8832
rect 5908 8984 5960 9036
rect 6644 8984 6696 9036
rect 4344 8916 4396 8968
rect 9404 8984 9456 9036
rect 12348 9120 12400 9172
rect 12532 9163 12584 9172
rect 12532 9129 12541 9163
rect 12541 9129 12575 9163
rect 12575 9129 12584 9163
rect 12532 9120 12584 9129
rect 15844 9120 15896 9172
rect 15936 9120 15988 9172
rect 17316 9120 17368 9172
rect 19800 9163 19852 9172
rect 13176 9052 13228 9104
rect 18696 9052 18748 9104
rect 19800 9129 19809 9163
rect 19809 9129 19843 9163
rect 19843 9129 19852 9163
rect 19800 9120 19852 9129
rect 20444 9120 20496 9172
rect 20260 9052 20312 9104
rect 12532 8984 12584 9036
rect 12808 8984 12860 9036
rect 21548 9120 21600 9172
rect 26056 9120 26108 9172
rect 26700 9163 26752 9172
rect 26700 9129 26709 9163
rect 26709 9129 26743 9163
rect 26743 9129 26752 9163
rect 26700 9120 26752 9129
rect 21640 9052 21692 9104
rect 21916 9052 21968 9104
rect 5908 8848 5960 8900
rect 9220 8916 9272 8968
rect 10508 8959 10560 8968
rect 10508 8925 10517 8959
rect 10517 8925 10551 8959
rect 10551 8925 10560 8959
rect 10508 8916 10560 8925
rect 11060 8916 11112 8968
rect 11704 8916 11756 8968
rect 11888 8916 11940 8968
rect 12900 8916 12952 8968
rect 13176 8959 13228 8968
rect 13176 8925 13185 8959
rect 13185 8925 13219 8959
rect 13219 8925 13228 8959
rect 13176 8916 13228 8925
rect 16948 8959 17000 8968
rect 16948 8925 16982 8959
rect 16982 8925 17000 8959
rect 8392 8848 8444 8900
rect 8484 8848 8536 8900
rect 9588 8848 9640 8900
rect 6644 8780 6696 8832
rect 8300 8823 8352 8832
rect 8300 8789 8309 8823
rect 8309 8789 8343 8823
rect 8343 8789 8352 8823
rect 8300 8780 8352 8789
rect 9036 8780 9088 8832
rect 9220 8780 9272 8832
rect 13636 8848 13688 8900
rect 15108 8848 15160 8900
rect 12164 8780 12216 8832
rect 12532 8780 12584 8832
rect 13360 8780 13412 8832
rect 14832 8780 14884 8832
rect 15476 8780 15528 8832
rect 16948 8916 17000 8925
rect 19248 8959 19300 8968
rect 17316 8780 17368 8832
rect 17776 8780 17828 8832
rect 19248 8925 19257 8959
rect 19257 8925 19291 8959
rect 19291 8925 19300 8959
rect 19248 8916 19300 8925
rect 19432 8959 19484 8968
rect 19432 8925 19441 8959
rect 19441 8925 19475 8959
rect 19475 8925 19484 8959
rect 19432 8916 19484 8925
rect 19340 8848 19392 8900
rect 19892 8916 19944 8968
rect 21088 8916 21140 8968
rect 20076 8848 20128 8900
rect 21548 8848 21600 8900
rect 22376 8916 22428 8968
rect 23204 8959 23256 8968
rect 23204 8925 23213 8959
rect 23213 8925 23247 8959
rect 23247 8925 23256 8959
rect 23204 8916 23256 8925
rect 23388 8848 23440 8900
rect 23848 8984 23900 9036
rect 24216 8916 24268 8968
rect 24768 8984 24820 9036
rect 24860 8848 24912 8900
rect 25504 8916 25556 8968
rect 26700 8916 26752 8968
rect 27344 8984 27396 9036
rect 27160 8959 27212 8968
rect 27160 8925 27169 8959
rect 27169 8925 27203 8959
rect 27203 8925 27212 8959
rect 27160 8916 27212 8925
rect 26608 8848 26660 8900
rect 20904 8780 20956 8832
rect 20996 8780 21048 8832
rect 21916 8780 21968 8832
rect 23940 8780 23992 8832
rect 26424 8780 26476 8832
rect 26884 8780 26936 8832
rect 9935 8678 9987 8730
rect 9999 8678 10051 8730
rect 10063 8678 10115 8730
rect 10127 8678 10179 8730
rect 10191 8678 10243 8730
rect 18920 8678 18972 8730
rect 18984 8678 19036 8730
rect 19048 8678 19100 8730
rect 19112 8678 19164 8730
rect 19176 8678 19228 8730
rect 2872 8576 2924 8628
rect 2596 8551 2648 8560
rect 2596 8517 2605 8551
rect 2605 8517 2639 8551
rect 2639 8517 2648 8551
rect 2596 8508 2648 8517
rect 6552 8576 6604 8628
rect 6644 8576 6696 8628
rect 10508 8576 10560 8628
rect 13176 8619 13228 8628
rect 13176 8585 13185 8619
rect 13185 8585 13219 8619
rect 13219 8585 13228 8619
rect 13176 8576 13228 8585
rect 13636 8619 13688 8628
rect 13636 8585 13645 8619
rect 13645 8585 13679 8619
rect 13679 8585 13688 8619
rect 13636 8576 13688 8585
rect 4620 8551 4672 8560
rect 4620 8517 4629 8551
rect 4629 8517 4663 8551
rect 4663 8517 4672 8551
rect 4620 8508 4672 8517
rect 9496 8551 9548 8560
rect 9496 8517 9505 8551
rect 9505 8517 9539 8551
rect 9539 8517 9548 8551
rect 9496 8508 9548 8517
rect 11612 8508 11664 8560
rect 12716 8508 12768 8560
rect 15200 8508 15252 8560
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 3976 8440 4028 8492
rect 5264 8483 5316 8492
rect 5264 8449 5273 8483
rect 5273 8449 5307 8483
rect 5307 8449 5316 8483
rect 5264 8440 5316 8449
rect 6644 8440 6696 8492
rect 8392 8440 8444 8492
rect 8668 8440 8720 8492
rect 9036 8440 9088 8492
rect 5356 8415 5408 8424
rect 5356 8381 5365 8415
rect 5365 8381 5399 8415
rect 5399 8381 5408 8415
rect 5356 8372 5408 8381
rect 6920 8415 6972 8424
rect 6920 8381 6929 8415
rect 6929 8381 6963 8415
rect 6963 8381 6972 8415
rect 6920 8372 6972 8381
rect 9496 8372 9548 8424
rect 11060 8440 11112 8492
rect 11152 8440 11204 8492
rect 11796 8483 11848 8492
rect 11796 8449 11805 8483
rect 11805 8449 11839 8483
rect 11839 8449 11848 8483
rect 11796 8440 11848 8449
rect 9864 8372 9916 8424
rect 12532 8440 12584 8492
rect 13176 8440 13228 8492
rect 13452 8440 13504 8492
rect 13636 8440 13688 8492
rect 13912 8440 13964 8492
rect 14832 8440 14884 8492
rect 15936 8576 15988 8628
rect 17040 8619 17092 8628
rect 17040 8585 17049 8619
rect 17049 8585 17083 8619
rect 17083 8585 17092 8619
rect 17040 8576 17092 8585
rect 15844 8508 15896 8560
rect 18420 8576 18472 8628
rect 19524 8576 19576 8628
rect 12348 8372 12400 8424
rect 2136 8304 2188 8356
rect 6736 8304 6788 8356
rect 8300 8304 8352 8356
rect 12532 8304 12584 8356
rect 12716 8304 12768 8356
rect 15844 8372 15896 8424
rect 16212 8372 16264 8424
rect 1860 8279 1912 8288
rect 1860 8245 1869 8279
rect 1869 8245 1903 8279
rect 1903 8245 1912 8279
rect 1860 8236 1912 8245
rect 4068 8236 4120 8288
rect 4252 8236 4304 8288
rect 4620 8236 4672 8288
rect 5356 8279 5408 8288
rect 5356 8245 5365 8279
rect 5365 8245 5399 8279
rect 5399 8245 5408 8279
rect 5356 8236 5408 8245
rect 6828 8236 6880 8288
rect 8668 8236 8720 8288
rect 11704 8236 11756 8288
rect 13360 8236 13412 8288
rect 13912 8236 13964 8288
rect 15292 8304 15344 8356
rect 15568 8304 15620 8356
rect 17776 8551 17828 8560
rect 17776 8517 17785 8551
rect 17785 8517 17819 8551
rect 17819 8517 17828 8551
rect 17776 8508 17828 8517
rect 19984 8576 20036 8628
rect 20260 8576 20312 8628
rect 21640 8576 21692 8628
rect 23664 8576 23716 8628
rect 25136 8576 25188 8628
rect 25320 8576 25372 8628
rect 27344 8576 27396 8628
rect 22744 8508 22796 8560
rect 23112 8551 23164 8560
rect 23112 8517 23121 8551
rect 23121 8517 23155 8551
rect 23155 8517 23164 8551
rect 23112 8508 23164 8517
rect 16948 8372 17000 8424
rect 19432 8372 19484 8424
rect 19708 8483 19760 8492
rect 19708 8449 19717 8483
rect 19717 8449 19751 8483
rect 19751 8449 19760 8483
rect 20812 8483 20864 8492
rect 19708 8440 19760 8449
rect 20812 8449 20821 8483
rect 20821 8449 20855 8483
rect 20855 8449 20864 8483
rect 20812 8440 20864 8449
rect 20904 8440 20956 8492
rect 25780 8508 25832 8560
rect 26056 8508 26108 8560
rect 27252 8508 27304 8560
rect 24124 8440 24176 8492
rect 24216 8440 24268 8492
rect 26148 8440 26200 8492
rect 26792 8440 26844 8492
rect 20076 8304 20128 8356
rect 21088 8304 21140 8356
rect 22744 8304 22796 8356
rect 23204 8372 23256 8424
rect 27252 8372 27304 8424
rect 16856 8236 16908 8288
rect 23204 8279 23256 8288
rect 23204 8245 23213 8279
rect 23213 8245 23247 8279
rect 23247 8245 23256 8279
rect 23204 8236 23256 8245
rect 24400 8279 24452 8288
rect 24400 8245 24409 8279
rect 24409 8245 24443 8279
rect 24443 8245 24452 8279
rect 24400 8236 24452 8245
rect 26516 8304 26568 8356
rect 26976 8236 27028 8288
rect 5442 8134 5494 8186
rect 5506 8134 5558 8186
rect 5570 8134 5622 8186
rect 5634 8134 5686 8186
rect 5698 8134 5750 8186
rect 14428 8134 14480 8186
rect 14492 8134 14544 8186
rect 14556 8134 14608 8186
rect 14620 8134 14672 8186
rect 14684 8134 14736 8186
rect 23413 8134 23465 8186
rect 23477 8134 23529 8186
rect 23541 8134 23593 8186
rect 23605 8134 23657 8186
rect 23669 8134 23721 8186
rect 3240 8032 3292 8084
rect 3976 8032 4028 8084
rect 4068 8032 4120 8084
rect 6736 8032 6788 8084
rect 7932 8032 7984 8084
rect 8208 8032 8260 8084
rect 13268 8032 13320 8084
rect 13452 8075 13504 8084
rect 13452 8041 13461 8075
rect 13461 8041 13495 8075
rect 13495 8041 13504 8075
rect 13452 8032 13504 8041
rect 15108 8075 15160 8084
rect 15108 8041 15117 8075
rect 15117 8041 15151 8075
rect 15151 8041 15160 8075
rect 15108 8032 15160 8041
rect 2780 7964 2832 8016
rect 3424 7964 3476 8016
rect 5264 7964 5316 8016
rect 7380 7964 7432 8016
rect 5816 7939 5868 7948
rect 5816 7905 5825 7939
rect 5825 7905 5859 7939
rect 5859 7905 5868 7939
rect 5816 7896 5868 7905
rect 6460 7896 6512 7948
rect 8944 7964 8996 8016
rect 11888 7964 11940 8016
rect 12072 8007 12124 8016
rect 12072 7973 12081 8007
rect 12081 7973 12115 8007
rect 12115 7973 12124 8007
rect 12072 7964 12124 7973
rect 11704 7896 11756 7948
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 3792 7871 3844 7880
rect 1584 7828 1636 7837
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 4620 7828 4672 7880
rect 6644 7871 6696 7880
rect 1860 7803 1912 7812
rect 1860 7769 1894 7803
rect 1894 7769 1912 7803
rect 1860 7760 1912 7769
rect 3424 7760 3476 7812
rect 3240 7692 3292 7744
rect 5264 7692 5316 7744
rect 6644 7837 6653 7871
rect 6653 7837 6687 7871
rect 6687 7837 6696 7871
rect 6644 7828 6696 7837
rect 6736 7828 6788 7880
rect 6368 7760 6420 7812
rect 8116 7828 8168 7880
rect 10048 7828 10100 7880
rect 10508 7828 10560 7880
rect 11060 7828 11112 7880
rect 11980 7828 12032 7880
rect 8944 7803 8996 7812
rect 6736 7692 6788 7744
rect 8944 7769 8953 7803
rect 8953 7769 8987 7803
rect 8987 7769 8996 7803
rect 8944 7760 8996 7769
rect 9496 7760 9548 7812
rect 10140 7760 10192 7812
rect 11336 7760 11388 7812
rect 12348 7760 12400 7812
rect 12716 7760 12768 7812
rect 13544 7964 13596 8016
rect 14188 7964 14240 8016
rect 13360 7896 13412 7948
rect 7932 7692 7984 7744
rect 11060 7692 11112 7744
rect 13544 7828 13596 7880
rect 14372 7871 14424 7880
rect 14372 7837 14381 7871
rect 14381 7837 14415 7871
rect 14415 7837 14424 7871
rect 14372 7828 14424 7837
rect 14832 7964 14884 8016
rect 15292 7871 15344 7880
rect 15292 7837 15301 7871
rect 15301 7837 15335 7871
rect 15335 7837 15344 7871
rect 15292 7828 15344 7837
rect 22008 8032 22060 8084
rect 19248 7964 19300 8016
rect 23112 8032 23164 8084
rect 26148 8032 26200 8084
rect 17316 7939 17368 7948
rect 17316 7905 17325 7939
rect 17325 7905 17359 7939
rect 17359 7905 17368 7939
rect 17316 7896 17368 7905
rect 18604 7896 18656 7948
rect 16212 7871 16264 7880
rect 16212 7837 16221 7871
rect 16221 7837 16255 7871
rect 16255 7837 16264 7871
rect 16212 7828 16264 7837
rect 17592 7871 17644 7880
rect 17592 7837 17626 7871
rect 17626 7837 17644 7871
rect 17592 7828 17644 7837
rect 19892 7828 19944 7880
rect 15568 7760 15620 7812
rect 16304 7760 16356 7812
rect 19248 7803 19300 7812
rect 19248 7769 19257 7803
rect 19257 7769 19291 7803
rect 19291 7769 19300 7803
rect 19248 7760 19300 7769
rect 19340 7760 19392 7812
rect 22192 7828 22244 7880
rect 23204 7828 23256 7880
rect 23296 7760 23348 7812
rect 24308 7828 24360 7880
rect 24584 7828 24636 7880
rect 25044 7828 25096 7880
rect 25964 7828 26016 7880
rect 26700 7828 26752 7880
rect 27160 7828 27212 7880
rect 15476 7692 15528 7744
rect 16948 7692 17000 7744
rect 17684 7692 17736 7744
rect 18144 7692 18196 7744
rect 21548 7735 21600 7744
rect 21548 7701 21557 7735
rect 21557 7701 21591 7735
rect 21591 7701 21600 7735
rect 21548 7692 21600 7701
rect 21916 7692 21968 7744
rect 24216 7760 24268 7812
rect 27988 7760 28040 7812
rect 23756 7692 23808 7744
rect 24584 7692 24636 7744
rect 26976 7692 27028 7744
rect 9935 7590 9987 7642
rect 9999 7590 10051 7642
rect 10063 7590 10115 7642
rect 10127 7590 10179 7642
rect 10191 7590 10243 7642
rect 18920 7590 18972 7642
rect 18984 7590 19036 7642
rect 19048 7590 19100 7642
rect 19112 7590 19164 7642
rect 19176 7590 19228 7642
rect 2044 7488 2096 7540
rect 2688 7488 2740 7540
rect 3792 7488 3844 7540
rect 6276 7488 6328 7540
rect 4252 7420 4304 7472
rect 2136 7352 2188 7404
rect 2780 7352 2832 7404
rect 3240 7395 3292 7404
rect 3240 7361 3249 7395
rect 3249 7361 3283 7395
rect 3283 7361 3292 7395
rect 3240 7352 3292 7361
rect 3700 7352 3752 7404
rect 4344 7395 4396 7404
rect 4344 7361 4353 7395
rect 4353 7361 4387 7395
rect 4387 7361 4396 7395
rect 4344 7352 4396 7361
rect 5264 7395 5316 7404
rect 5264 7361 5273 7395
rect 5273 7361 5307 7395
rect 5307 7361 5316 7395
rect 5264 7352 5316 7361
rect 6828 7420 6880 7472
rect 7748 7420 7800 7472
rect 6460 7395 6512 7404
rect 2596 7284 2648 7336
rect 2872 7284 2924 7336
rect 6460 7361 6469 7395
rect 6469 7361 6503 7395
rect 6503 7361 6512 7395
rect 6460 7352 6512 7361
rect 2780 7216 2832 7268
rect 4068 7216 4120 7268
rect 4252 7148 4304 7200
rect 6368 7284 6420 7336
rect 7840 7352 7892 7404
rect 9864 7352 9916 7404
rect 6920 7284 6972 7336
rect 8208 7327 8260 7336
rect 8208 7293 8217 7327
rect 8217 7293 8251 7327
rect 8251 7293 8260 7327
rect 8208 7284 8260 7293
rect 10600 7488 10652 7540
rect 12532 7488 12584 7540
rect 12624 7463 12676 7472
rect 10232 7352 10284 7404
rect 11520 7284 11572 7336
rect 11796 7395 11848 7404
rect 11796 7361 11805 7395
rect 11805 7361 11839 7395
rect 11839 7361 11848 7395
rect 12624 7429 12633 7463
rect 12633 7429 12667 7463
rect 12667 7429 12676 7463
rect 12624 7420 12676 7429
rect 14188 7420 14240 7472
rect 17868 7488 17920 7540
rect 19248 7488 19300 7540
rect 20628 7488 20680 7540
rect 11796 7352 11848 7361
rect 13544 7352 13596 7404
rect 15200 7352 15252 7404
rect 16120 7395 16172 7404
rect 9404 7216 9456 7268
rect 12348 7284 12400 7336
rect 16120 7361 16129 7395
rect 16129 7361 16163 7395
rect 16163 7361 16172 7395
rect 16120 7352 16172 7361
rect 16580 7420 16632 7472
rect 16764 7395 16816 7404
rect 15660 7284 15712 7336
rect 16764 7361 16773 7395
rect 16773 7361 16807 7395
rect 16807 7361 16816 7395
rect 16764 7352 16816 7361
rect 16948 7395 17000 7404
rect 16948 7361 16957 7395
rect 16957 7361 16991 7395
rect 16991 7361 17000 7395
rect 16948 7352 17000 7361
rect 17592 7395 17644 7404
rect 17592 7361 17601 7395
rect 17601 7361 17635 7395
rect 17635 7361 17644 7395
rect 17592 7352 17644 7361
rect 19064 7395 19116 7404
rect 19064 7361 19073 7395
rect 19073 7361 19107 7395
rect 19107 7361 19116 7395
rect 19064 7352 19116 7361
rect 21548 7420 21600 7472
rect 23664 7488 23716 7540
rect 19432 7395 19484 7404
rect 19432 7361 19441 7395
rect 19441 7361 19475 7395
rect 19475 7361 19484 7395
rect 19432 7352 19484 7361
rect 19616 7352 19668 7404
rect 19340 7284 19392 7336
rect 20168 7352 20220 7404
rect 20444 7352 20496 7404
rect 20904 7395 20956 7404
rect 20904 7361 20913 7395
rect 20913 7361 20947 7395
rect 20947 7361 20956 7395
rect 20904 7352 20956 7361
rect 16304 7216 16356 7268
rect 16764 7216 16816 7268
rect 17868 7216 17920 7268
rect 9588 7191 9640 7200
rect 9588 7157 9597 7191
rect 9597 7157 9631 7191
rect 9631 7157 9640 7191
rect 9588 7148 9640 7157
rect 12532 7148 12584 7200
rect 13912 7191 13964 7200
rect 13912 7157 13921 7191
rect 13921 7157 13955 7191
rect 13955 7157 13964 7191
rect 13912 7148 13964 7157
rect 15292 7148 15344 7200
rect 15476 7148 15528 7200
rect 16396 7148 16448 7200
rect 19064 7148 19116 7200
rect 19340 7191 19392 7200
rect 19340 7157 19349 7191
rect 19349 7157 19383 7191
rect 19383 7157 19392 7191
rect 19340 7148 19392 7157
rect 20444 7148 20496 7200
rect 23756 7463 23808 7472
rect 23756 7429 23765 7463
rect 23765 7429 23799 7463
rect 23799 7429 23808 7463
rect 23756 7420 23808 7429
rect 24216 7488 24268 7540
rect 24308 7420 24360 7472
rect 24584 7463 24636 7472
rect 24584 7429 24593 7463
rect 24593 7429 24627 7463
rect 24627 7429 24636 7463
rect 24584 7420 24636 7429
rect 23112 7395 23164 7404
rect 23112 7361 23121 7395
rect 23121 7361 23155 7395
rect 23155 7361 23164 7395
rect 25964 7488 26016 7540
rect 27160 7531 27212 7540
rect 23112 7352 23164 7361
rect 24308 7284 24360 7336
rect 24952 7352 25004 7404
rect 25504 7352 25556 7404
rect 26148 7420 26200 7472
rect 27160 7497 27195 7531
rect 27195 7497 27212 7531
rect 27160 7488 27212 7497
rect 27528 7488 27580 7540
rect 26884 7420 26936 7472
rect 26700 7352 26752 7404
rect 27344 7352 27396 7404
rect 26148 7284 26200 7336
rect 22468 7216 22520 7268
rect 24216 7216 24268 7268
rect 27068 7216 27120 7268
rect 23204 7148 23256 7200
rect 24860 7148 24912 7200
rect 25044 7148 25096 7200
rect 26240 7191 26292 7200
rect 26240 7157 26249 7191
rect 26249 7157 26283 7191
rect 26283 7157 26292 7191
rect 26240 7148 26292 7157
rect 27436 7148 27488 7200
rect 5442 7046 5494 7098
rect 5506 7046 5558 7098
rect 5570 7046 5622 7098
rect 5634 7046 5686 7098
rect 5698 7046 5750 7098
rect 14428 7046 14480 7098
rect 14492 7046 14544 7098
rect 14556 7046 14608 7098
rect 14620 7046 14672 7098
rect 14684 7046 14736 7098
rect 23413 7046 23465 7098
rect 23477 7046 23529 7098
rect 23541 7046 23593 7098
rect 23605 7046 23657 7098
rect 23669 7046 23721 7098
rect 2596 6944 2648 6996
rect 2964 6944 3016 6996
rect 6368 6944 6420 6996
rect 3608 6808 3660 6860
rect 7012 6876 7064 6928
rect 7748 6808 7800 6860
rect 11060 6944 11112 6996
rect 12716 6987 12768 6996
rect 12716 6953 12725 6987
rect 12725 6953 12759 6987
rect 12759 6953 12768 6987
rect 12716 6944 12768 6953
rect 13544 6944 13596 6996
rect 14924 6944 14976 6996
rect 15752 6944 15804 6996
rect 9220 6876 9272 6928
rect 9496 6876 9548 6928
rect 10232 6876 10284 6928
rect 12992 6876 13044 6928
rect 13360 6876 13412 6928
rect 19340 6876 19392 6928
rect 10416 6851 10468 6860
rect 1952 6715 2004 6724
rect 1952 6681 1961 6715
rect 1961 6681 1995 6715
rect 1995 6681 2004 6715
rect 1952 6672 2004 6681
rect 3608 6672 3660 6724
rect 5080 6715 5132 6724
rect 5080 6681 5089 6715
rect 5089 6681 5123 6715
rect 5123 6681 5132 6715
rect 5080 6672 5132 6681
rect 6552 6672 6604 6724
rect 7012 6672 7064 6724
rect 7840 6783 7892 6792
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 8208 6740 8260 6792
rect 10416 6817 10425 6851
rect 10425 6817 10459 6851
rect 10459 6817 10468 6851
rect 10416 6808 10468 6817
rect 9220 6783 9272 6792
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 12348 6740 12400 6792
rect 12624 6783 12676 6792
rect 12624 6749 12635 6783
rect 12635 6749 12676 6783
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 3332 6604 3384 6656
rect 5908 6647 5960 6656
rect 5908 6613 5917 6647
rect 5917 6613 5951 6647
rect 5951 6613 5960 6647
rect 5908 6604 5960 6613
rect 11704 6672 11756 6724
rect 12624 6740 12676 6749
rect 13728 6808 13780 6860
rect 19616 6808 19668 6860
rect 21180 6944 21232 6996
rect 24400 6944 24452 6996
rect 24676 6944 24728 6996
rect 24860 6944 24912 6996
rect 26240 6944 26292 6996
rect 27344 6987 27396 6996
rect 27344 6953 27353 6987
rect 27353 6953 27387 6987
rect 27387 6953 27396 6987
rect 27344 6944 27396 6953
rect 22652 6876 22704 6928
rect 12900 6740 12952 6792
rect 14924 6740 14976 6792
rect 12716 6672 12768 6724
rect 14280 6672 14332 6724
rect 17316 6740 17368 6792
rect 17500 6783 17552 6792
rect 17500 6749 17534 6783
rect 17534 6749 17552 6783
rect 17500 6740 17552 6749
rect 19064 6740 19116 6792
rect 19708 6740 19760 6792
rect 21640 6808 21692 6860
rect 19892 6740 19944 6792
rect 22192 6740 22244 6792
rect 25504 6808 25556 6860
rect 24032 6740 24084 6792
rect 24216 6740 24268 6792
rect 15292 6715 15344 6724
rect 15292 6681 15326 6715
rect 15326 6681 15344 6715
rect 15292 6672 15344 6681
rect 15568 6672 15620 6724
rect 21824 6672 21876 6724
rect 24400 6715 24452 6724
rect 10600 6604 10652 6656
rect 11796 6647 11848 6656
rect 11796 6613 11805 6647
rect 11805 6613 11839 6647
rect 11839 6613 11848 6647
rect 11796 6604 11848 6613
rect 12440 6604 12492 6656
rect 13268 6647 13320 6656
rect 13268 6613 13277 6647
rect 13277 6613 13311 6647
rect 13311 6613 13320 6647
rect 13268 6604 13320 6613
rect 14924 6604 14976 6656
rect 15936 6604 15988 6656
rect 17868 6604 17920 6656
rect 22008 6604 22060 6656
rect 23020 6647 23072 6656
rect 23020 6613 23029 6647
rect 23029 6613 23063 6647
rect 23063 6613 23072 6647
rect 23020 6604 23072 6613
rect 24032 6604 24084 6656
rect 24400 6681 24409 6715
rect 24409 6681 24443 6715
rect 24443 6681 24452 6715
rect 24400 6672 24452 6681
rect 24768 6604 24820 6656
rect 24952 6604 25004 6656
rect 9935 6502 9987 6554
rect 9999 6502 10051 6554
rect 10063 6502 10115 6554
rect 10127 6502 10179 6554
rect 10191 6502 10243 6554
rect 18920 6502 18972 6554
rect 18984 6502 19036 6554
rect 19048 6502 19100 6554
rect 19112 6502 19164 6554
rect 19176 6502 19228 6554
rect 5356 6400 5408 6452
rect 8944 6400 8996 6452
rect 9680 6400 9732 6452
rect 15292 6400 15344 6452
rect 16672 6400 16724 6452
rect 17592 6400 17644 6452
rect 17868 6400 17920 6452
rect 22560 6400 22612 6452
rect 24308 6443 24360 6452
rect 1400 6196 1452 6248
rect 1584 6264 1636 6316
rect 2320 6264 2372 6316
rect 6276 6264 6328 6316
rect 6920 6332 6972 6384
rect 8484 6375 8536 6384
rect 8484 6341 8493 6375
rect 8493 6341 8527 6375
rect 8527 6341 8536 6375
rect 8484 6332 8536 6341
rect 2688 6196 2740 6248
rect 5816 6196 5868 6248
rect 8944 6264 8996 6316
rect 9220 6264 9272 6316
rect 8484 6196 8536 6248
rect 9588 6264 9640 6316
rect 11060 6332 11112 6384
rect 11520 6332 11572 6384
rect 9864 6264 9916 6316
rect 9496 6128 9548 6180
rect 10416 6264 10468 6316
rect 12532 6332 12584 6384
rect 13268 6332 13320 6384
rect 13360 6332 13412 6384
rect 13912 6332 13964 6384
rect 14832 6307 14884 6316
rect 14832 6273 14841 6307
rect 14841 6273 14875 6307
rect 14875 6273 14884 6307
rect 14832 6264 14884 6273
rect 16212 6332 16264 6384
rect 11520 6239 11572 6248
rect 11520 6205 11529 6239
rect 11529 6205 11563 6239
rect 11563 6205 11572 6239
rect 11520 6196 11572 6205
rect 12716 6196 12768 6248
rect 14740 6196 14792 6248
rect 15292 6196 15344 6248
rect 16396 6264 16448 6316
rect 17960 6332 18012 6384
rect 19708 6332 19760 6384
rect 20168 6375 20220 6384
rect 17592 6264 17644 6316
rect 18420 6264 18472 6316
rect 19432 6307 19484 6316
rect 19432 6273 19441 6307
rect 19441 6273 19475 6307
rect 19475 6273 19484 6307
rect 19432 6264 19484 6273
rect 19892 6307 19944 6316
rect 19892 6273 19901 6307
rect 19901 6273 19935 6307
rect 19935 6273 19944 6307
rect 19892 6264 19944 6273
rect 20168 6341 20202 6375
rect 20202 6341 20220 6375
rect 20168 6332 20220 6341
rect 20720 6332 20772 6384
rect 21640 6332 21692 6384
rect 22008 6264 22060 6316
rect 22192 6264 22244 6316
rect 22652 6264 22704 6316
rect 24308 6409 24317 6443
rect 24317 6409 24351 6443
rect 24351 6409 24360 6443
rect 24308 6400 24360 6409
rect 24768 6400 24820 6452
rect 25228 6400 25280 6452
rect 26240 6400 26292 6452
rect 27160 6443 27212 6452
rect 27160 6409 27185 6443
rect 27185 6409 27212 6443
rect 27344 6443 27396 6452
rect 27160 6400 27212 6409
rect 27344 6409 27353 6443
rect 27353 6409 27387 6443
rect 27387 6409 27396 6443
rect 27344 6400 27396 6409
rect 24216 6332 24268 6384
rect 25044 6375 25096 6384
rect 25044 6341 25078 6375
rect 25078 6341 25096 6375
rect 25044 6332 25096 6341
rect 25964 6332 26016 6384
rect 24768 6307 24820 6316
rect 11980 6128 12032 6180
rect 2780 6060 2832 6112
rect 3056 6060 3108 6112
rect 7012 6060 7064 6112
rect 8208 6060 8260 6112
rect 9404 6060 9456 6112
rect 10968 6060 11020 6112
rect 11704 6060 11756 6112
rect 12164 6060 12216 6112
rect 13544 6060 13596 6112
rect 13728 6060 13780 6112
rect 13912 6060 13964 6112
rect 16396 6060 16448 6112
rect 19340 6196 19392 6248
rect 18236 6128 18288 6180
rect 19708 6128 19760 6180
rect 19892 6128 19944 6180
rect 17592 6060 17644 6112
rect 18604 6103 18656 6112
rect 18604 6069 18613 6103
rect 18613 6069 18647 6103
rect 18647 6069 18656 6103
rect 18604 6060 18656 6069
rect 20812 6060 20864 6112
rect 22100 6060 22152 6112
rect 24768 6273 24777 6307
rect 24777 6273 24811 6307
rect 24811 6273 24820 6307
rect 24768 6264 24820 6273
rect 24676 6128 24728 6180
rect 24308 6060 24360 6112
rect 27896 6128 27948 6180
rect 25964 6060 26016 6112
rect 27436 6060 27488 6112
rect 5442 5958 5494 6010
rect 5506 5958 5558 6010
rect 5570 5958 5622 6010
rect 5634 5958 5686 6010
rect 5698 5958 5750 6010
rect 14428 5958 14480 6010
rect 14492 5958 14544 6010
rect 14556 5958 14608 6010
rect 14620 5958 14672 6010
rect 14684 5958 14736 6010
rect 23413 5958 23465 6010
rect 23477 5958 23529 6010
rect 23541 5958 23593 6010
rect 23605 5958 23657 6010
rect 23669 5958 23721 6010
rect 1952 5856 2004 5908
rect 4252 5856 4304 5908
rect 5080 5899 5132 5908
rect 5080 5865 5089 5899
rect 5089 5865 5123 5899
rect 5123 5865 5132 5899
rect 5080 5856 5132 5865
rect 5908 5856 5960 5908
rect 12992 5856 13044 5908
rect 13728 5856 13780 5908
rect 20812 5899 20864 5908
rect 2872 5788 2924 5840
rect 2964 5788 3016 5840
rect 4068 5788 4120 5840
rect 7288 5788 7340 5840
rect 10232 5788 10284 5840
rect 12716 5788 12768 5840
rect 2780 5652 2832 5704
rect 3056 5720 3108 5772
rect 4896 5720 4948 5772
rect 3240 5695 3292 5704
rect 3240 5661 3249 5695
rect 3249 5661 3283 5695
rect 3283 5661 3292 5695
rect 3240 5652 3292 5661
rect 4252 5652 4304 5704
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 5356 5695 5408 5704
rect 5356 5661 5365 5695
rect 5365 5661 5399 5695
rect 5399 5661 5408 5695
rect 8484 5720 8536 5772
rect 9404 5763 9456 5772
rect 9404 5729 9413 5763
rect 9413 5729 9447 5763
rect 9447 5729 9456 5763
rect 9404 5720 9456 5729
rect 10416 5720 10468 5772
rect 13544 5788 13596 5840
rect 14188 5788 14240 5840
rect 15660 5831 15712 5840
rect 15660 5797 15669 5831
rect 15669 5797 15703 5831
rect 15703 5797 15712 5831
rect 15660 5788 15712 5797
rect 16396 5788 16448 5840
rect 20812 5865 20821 5899
rect 20821 5865 20855 5899
rect 20855 5865 20864 5899
rect 20812 5856 20864 5865
rect 20996 5899 21048 5908
rect 20996 5865 21005 5899
rect 21005 5865 21039 5899
rect 21039 5865 21048 5899
rect 20996 5856 21048 5865
rect 21916 5856 21968 5908
rect 22468 5899 22520 5908
rect 22468 5865 22477 5899
rect 22477 5865 22511 5899
rect 22511 5865 22520 5899
rect 22468 5856 22520 5865
rect 23020 5856 23072 5908
rect 5356 5652 5408 5661
rect 9220 5695 9272 5704
rect 9220 5661 9229 5695
rect 9229 5661 9263 5695
rect 9263 5661 9272 5695
rect 9220 5652 9272 5661
rect 3056 5584 3108 5636
rect 6644 5627 6696 5636
rect 6644 5593 6653 5627
rect 6653 5593 6687 5627
rect 6687 5593 6696 5627
rect 6644 5584 6696 5593
rect 8484 5584 8536 5636
rect 11336 5652 11388 5704
rect 12716 5652 12768 5704
rect 14832 5720 14884 5772
rect 17316 5763 17368 5772
rect 13544 5695 13596 5704
rect 9680 5584 9732 5636
rect 3424 5516 3476 5568
rect 4804 5516 4856 5568
rect 7288 5516 7340 5568
rect 8760 5516 8812 5568
rect 9404 5516 9456 5568
rect 9496 5516 9548 5568
rect 11888 5559 11940 5568
rect 11888 5525 11897 5559
rect 11897 5525 11931 5559
rect 11931 5525 11940 5559
rect 11888 5516 11940 5525
rect 12808 5516 12860 5568
rect 12992 5559 13044 5568
rect 12992 5525 13001 5559
rect 13001 5525 13035 5559
rect 13035 5525 13044 5559
rect 12992 5516 13044 5525
rect 13544 5661 13553 5695
rect 13553 5661 13587 5695
rect 13587 5661 13596 5695
rect 13544 5652 13596 5661
rect 15752 5695 15804 5704
rect 13912 5584 13964 5636
rect 15108 5584 15160 5636
rect 15292 5584 15344 5636
rect 15752 5661 15761 5695
rect 15761 5661 15795 5695
rect 15795 5661 15804 5695
rect 15752 5652 15804 5661
rect 17316 5729 17325 5763
rect 17325 5729 17359 5763
rect 17359 5729 17368 5763
rect 17316 5720 17368 5729
rect 19616 5720 19668 5772
rect 16764 5695 16816 5704
rect 16764 5661 16773 5695
rect 16773 5661 16807 5695
rect 16807 5661 16816 5695
rect 16764 5652 16816 5661
rect 17040 5652 17092 5704
rect 19340 5652 19392 5704
rect 20076 5695 20128 5704
rect 20076 5661 20085 5695
rect 20085 5661 20119 5695
rect 20119 5661 20128 5695
rect 20076 5652 20128 5661
rect 15660 5516 15712 5568
rect 16212 5559 16264 5568
rect 16212 5525 16221 5559
rect 16221 5525 16255 5559
rect 16255 5525 16264 5559
rect 16212 5516 16264 5525
rect 16764 5516 16816 5568
rect 17592 5516 17644 5568
rect 20720 5584 20772 5636
rect 21180 5652 21232 5704
rect 22284 5720 22336 5772
rect 23848 5788 23900 5840
rect 22836 5720 22888 5772
rect 24676 5856 24728 5908
rect 24492 5788 24544 5840
rect 23112 5695 23164 5704
rect 21824 5584 21876 5636
rect 22100 5627 22152 5636
rect 22100 5593 22109 5627
rect 22109 5593 22143 5627
rect 22143 5593 22152 5627
rect 22100 5584 22152 5593
rect 23112 5661 23121 5695
rect 23121 5661 23155 5695
rect 23155 5661 23164 5695
rect 23112 5652 23164 5661
rect 23756 5652 23808 5704
rect 24308 5584 24360 5636
rect 24584 5652 24636 5704
rect 24768 5720 24820 5772
rect 25504 5720 25556 5772
rect 25688 5652 25740 5704
rect 27712 5652 27764 5704
rect 19248 5559 19300 5568
rect 19248 5525 19257 5559
rect 19257 5525 19291 5559
rect 19291 5525 19300 5559
rect 19248 5516 19300 5525
rect 19892 5559 19944 5568
rect 19892 5525 19901 5559
rect 19901 5525 19935 5559
rect 19935 5525 19944 5559
rect 19892 5516 19944 5525
rect 20536 5516 20588 5568
rect 22652 5516 22704 5568
rect 23848 5516 23900 5568
rect 24216 5516 24268 5568
rect 24584 5559 24636 5568
rect 28172 5584 28224 5636
rect 24584 5525 24609 5559
rect 24609 5525 24636 5559
rect 24584 5516 24636 5525
rect 26884 5516 26936 5568
rect 27344 5559 27396 5568
rect 27344 5525 27353 5559
rect 27353 5525 27387 5559
rect 27387 5525 27396 5559
rect 27344 5516 27396 5525
rect 9935 5414 9987 5466
rect 9999 5414 10051 5466
rect 10063 5414 10115 5466
rect 10127 5414 10179 5466
rect 10191 5414 10243 5466
rect 18920 5414 18972 5466
rect 18984 5414 19036 5466
rect 19048 5414 19100 5466
rect 19112 5414 19164 5466
rect 19176 5414 19228 5466
rect 3056 5355 3108 5364
rect 3056 5321 3065 5355
rect 3065 5321 3099 5355
rect 3099 5321 3108 5355
rect 3056 5312 3108 5321
rect 3884 5312 3936 5364
rect 6644 5355 6696 5364
rect 3608 5176 3660 5228
rect 4252 5244 4304 5296
rect 3792 5108 3844 5160
rect 4068 5219 4120 5228
rect 4068 5185 4077 5219
rect 4077 5185 4111 5219
rect 4111 5185 4120 5219
rect 6644 5321 6653 5355
rect 6653 5321 6687 5355
rect 6687 5321 6696 5355
rect 6644 5312 6696 5321
rect 7012 5312 7064 5364
rect 7564 5312 7616 5364
rect 8760 5312 8812 5364
rect 9220 5355 9272 5364
rect 9220 5321 9229 5355
rect 9229 5321 9263 5355
rect 9263 5321 9272 5355
rect 9220 5312 9272 5321
rect 9864 5312 9916 5364
rect 6460 5244 6512 5296
rect 4068 5176 4120 5185
rect 5264 5176 5316 5228
rect 6644 5176 6696 5228
rect 7288 5244 7340 5296
rect 7196 5219 7248 5228
rect 7196 5185 7205 5219
rect 7205 5185 7239 5219
rect 7239 5185 7248 5219
rect 7196 5176 7248 5185
rect 7564 5176 7616 5228
rect 11060 5312 11112 5364
rect 12808 5312 12860 5364
rect 15660 5355 15712 5364
rect 11888 5244 11940 5296
rect 12440 5287 12492 5296
rect 12440 5253 12449 5287
rect 12449 5253 12483 5287
rect 12483 5253 12492 5287
rect 12440 5244 12492 5253
rect 12992 5244 13044 5296
rect 15660 5321 15669 5355
rect 15669 5321 15703 5355
rect 15703 5321 15712 5355
rect 15660 5312 15712 5321
rect 20628 5355 20680 5364
rect 20628 5321 20637 5355
rect 20637 5321 20671 5355
rect 20671 5321 20680 5355
rect 20628 5312 20680 5321
rect 20812 5312 20864 5364
rect 21916 5312 21968 5364
rect 23480 5312 23532 5364
rect 10508 5219 10560 5228
rect 10508 5185 10517 5219
rect 10517 5185 10551 5219
rect 10551 5185 10560 5219
rect 10508 5176 10560 5185
rect 11428 5176 11480 5228
rect 12256 5176 12308 5228
rect 7012 5108 7064 5160
rect 7840 5151 7892 5160
rect 7840 5117 7849 5151
rect 7849 5117 7883 5151
rect 7883 5117 7892 5151
rect 7840 5108 7892 5117
rect 11520 5108 11572 5160
rect 12900 5176 12952 5228
rect 13912 5176 13964 5228
rect 14280 5219 14332 5228
rect 14280 5185 14289 5219
rect 14289 5185 14323 5219
rect 14323 5185 14332 5219
rect 14280 5176 14332 5185
rect 17316 5244 17368 5296
rect 18052 5244 18104 5296
rect 16304 5108 16356 5160
rect 18420 5176 18472 5228
rect 20352 5244 20404 5296
rect 20536 5244 20588 5296
rect 22468 5244 22520 5296
rect 18052 5108 18104 5160
rect 4344 5040 4396 5092
rect 4896 5040 4948 5092
rect 5264 5040 5316 5092
rect 7196 5040 7248 5092
rect 7472 5040 7524 5092
rect 12716 5040 12768 5092
rect 20536 5108 20588 5160
rect 21640 5176 21692 5228
rect 22560 5176 22612 5228
rect 22928 5244 22980 5296
rect 23664 5244 23716 5296
rect 24216 5244 24268 5296
rect 24400 5287 24452 5296
rect 24400 5253 24409 5287
rect 24409 5253 24443 5287
rect 24443 5253 24452 5287
rect 24400 5244 24452 5253
rect 24584 5287 24636 5296
rect 24584 5253 24609 5287
rect 24609 5253 24636 5287
rect 24584 5244 24636 5253
rect 24860 5244 24912 5296
rect 26976 5287 27028 5296
rect 26976 5253 26985 5287
rect 26985 5253 27019 5287
rect 27019 5253 27028 5287
rect 26976 5244 27028 5253
rect 22744 5108 22796 5160
rect 23020 5108 23072 5160
rect 25688 5108 25740 5160
rect 26884 5108 26936 5160
rect 26976 5108 27028 5160
rect 26148 5040 26200 5092
rect 1860 4972 1912 5024
rect 5816 4972 5868 5024
rect 6920 4972 6972 5024
rect 8208 4972 8260 5024
rect 11796 5015 11848 5024
rect 11796 4981 11805 5015
rect 11805 4981 11839 5015
rect 11839 4981 11848 5015
rect 11796 4972 11848 4981
rect 11980 5015 12032 5024
rect 11980 4981 11989 5015
rect 11989 4981 12023 5015
rect 12023 4981 12032 5015
rect 11980 4972 12032 4981
rect 15384 4972 15436 5024
rect 18420 4972 18472 5024
rect 20352 4972 20404 5024
rect 20812 4972 20864 5024
rect 20996 4972 21048 5024
rect 21824 5015 21876 5024
rect 21824 4981 21833 5015
rect 21833 4981 21867 5015
rect 21867 4981 21876 5015
rect 21824 4972 21876 4981
rect 22744 4972 22796 5024
rect 24216 4972 24268 5024
rect 24575 5015 24627 5024
rect 24575 4981 24584 5015
rect 24584 4981 24618 5015
rect 24618 4981 24627 5015
rect 24575 4972 24627 4981
rect 26884 4972 26936 5024
rect 5442 4870 5494 4922
rect 5506 4870 5558 4922
rect 5570 4870 5622 4922
rect 5634 4870 5686 4922
rect 5698 4870 5750 4922
rect 14428 4870 14480 4922
rect 14492 4870 14544 4922
rect 14556 4870 14608 4922
rect 14620 4870 14672 4922
rect 14684 4870 14736 4922
rect 23413 4870 23465 4922
rect 23477 4870 23529 4922
rect 23541 4870 23593 4922
rect 23605 4870 23657 4922
rect 23669 4870 23721 4922
rect 3792 4811 3844 4820
rect 3792 4777 3801 4811
rect 3801 4777 3835 4811
rect 3835 4777 3844 4811
rect 3792 4768 3844 4777
rect 4252 4768 4304 4820
rect 4896 4768 4948 4820
rect 8024 4768 8076 4820
rect 9588 4811 9640 4820
rect 9588 4777 9597 4811
rect 9597 4777 9631 4811
rect 9631 4777 9640 4811
rect 9588 4768 9640 4777
rect 11520 4768 11572 4820
rect 17132 4811 17184 4820
rect 17132 4777 17141 4811
rect 17141 4777 17175 4811
rect 17175 4777 17184 4811
rect 17132 4768 17184 4777
rect 17592 4768 17644 4820
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 2688 4564 2740 4616
rect 4344 4700 4396 4752
rect 6276 4700 6328 4752
rect 8300 4700 8352 4752
rect 8484 4700 8536 4752
rect 10600 4700 10652 4752
rect 11888 4700 11940 4752
rect 20352 4768 20404 4820
rect 20536 4700 20588 4752
rect 22100 4700 22152 4752
rect 6736 4632 6788 4684
rect 7012 4632 7064 4684
rect 7472 4632 7524 4684
rect 1676 4539 1728 4548
rect 1676 4505 1710 4539
rect 1710 4505 1728 4539
rect 4712 4564 4764 4616
rect 5080 4607 5132 4616
rect 5080 4573 5089 4607
rect 5089 4573 5123 4607
rect 5123 4573 5132 4607
rect 5080 4564 5132 4573
rect 6552 4564 6604 4616
rect 11980 4632 12032 4684
rect 1676 4496 1728 4505
rect 4252 4496 4304 4548
rect 5356 4539 5408 4548
rect 5356 4505 5390 4539
rect 5390 4505 5408 4539
rect 9220 4564 9272 4616
rect 9496 4607 9548 4616
rect 9496 4573 9505 4607
rect 9505 4573 9539 4607
rect 9539 4573 9548 4607
rect 9496 4564 9548 4573
rect 9864 4564 9916 4616
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 11704 4607 11756 4616
rect 11704 4573 11713 4607
rect 11713 4573 11747 4607
rect 11747 4573 11756 4607
rect 11704 4564 11756 4573
rect 12808 4564 12860 4616
rect 14096 4564 14148 4616
rect 16396 4632 16448 4684
rect 17316 4632 17368 4684
rect 22836 4700 22888 4752
rect 15476 4607 15528 4616
rect 5356 4496 5408 4505
rect 6736 4428 6788 4480
rect 10784 4496 10836 4548
rect 12532 4496 12584 4548
rect 12716 4496 12768 4548
rect 13176 4496 13228 4548
rect 15476 4573 15485 4607
rect 15485 4573 15519 4607
rect 15519 4573 15528 4607
rect 15476 4564 15528 4573
rect 16212 4564 16264 4616
rect 15292 4496 15344 4548
rect 16672 4496 16724 4548
rect 20536 4564 20588 4616
rect 22284 4632 22336 4684
rect 19064 4496 19116 4548
rect 20260 4496 20312 4548
rect 21824 4496 21876 4548
rect 13268 4428 13320 4480
rect 13820 4428 13872 4480
rect 14832 4428 14884 4480
rect 15200 4428 15252 4480
rect 16580 4428 16632 4480
rect 17960 4428 18012 4480
rect 20628 4471 20680 4480
rect 20628 4437 20637 4471
rect 20637 4437 20671 4471
rect 20671 4437 20680 4471
rect 20628 4428 20680 4437
rect 21548 4428 21600 4480
rect 23020 4564 23072 4616
rect 23296 4700 23348 4752
rect 24308 4768 24360 4820
rect 26148 4768 26200 4820
rect 26884 4811 26936 4820
rect 26884 4777 26893 4811
rect 26893 4777 26927 4811
rect 26927 4777 26936 4811
rect 26884 4768 26936 4777
rect 25780 4700 25832 4752
rect 23388 4607 23440 4616
rect 23388 4573 23397 4607
rect 23397 4573 23431 4607
rect 23431 4573 23440 4607
rect 23388 4564 23440 4573
rect 24308 4564 24360 4616
rect 22560 4496 22612 4548
rect 27160 4564 27212 4616
rect 24860 4539 24912 4548
rect 24860 4505 24894 4539
rect 24894 4505 24912 4539
rect 26700 4539 26752 4548
rect 24860 4496 24912 4505
rect 26700 4505 26709 4539
rect 26709 4505 26743 4539
rect 26743 4505 26752 4539
rect 26700 4496 26752 4505
rect 26976 4496 27028 4548
rect 22468 4471 22520 4480
rect 22468 4437 22477 4471
rect 22477 4437 22511 4471
rect 22511 4437 22520 4471
rect 22468 4428 22520 4437
rect 22928 4471 22980 4480
rect 22928 4437 22937 4471
rect 22937 4437 22971 4471
rect 22971 4437 22980 4471
rect 22928 4428 22980 4437
rect 23480 4428 23532 4480
rect 24400 4428 24452 4480
rect 9935 4326 9987 4378
rect 9999 4326 10051 4378
rect 10063 4326 10115 4378
rect 10127 4326 10179 4378
rect 10191 4326 10243 4378
rect 18920 4326 18972 4378
rect 18984 4326 19036 4378
rect 19048 4326 19100 4378
rect 19112 4326 19164 4378
rect 19176 4326 19228 4378
rect 1676 4267 1728 4276
rect 1676 4233 1685 4267
rect 1685 4233 1719 4267
rect 1719 4233 1728 4267
rect 1676 4224 1728 4233
rect 3424 4224 3476 4276
rect 4344 4224 4396 4276
rect 4896 4267 4948 4276
rect 4896 4233 4905 4267
rect 4905 4233 4939 4267
rect 4939 4233 4948 4267
rect 4896 4224 4948 4233
rect 5356 4267 5408 4276
rect 5356 4233 5365 4267
rect 5365 4233 5399 4267
rect 5399 4233 5408 4267
rect 5356 4224 5408 4233
rect 2964 4156 3016 4208
rect 848 4088 900 4140
rect 1492 4088 1544 4140
rect 1860 4131 1912 4140
rect 1860 4097 1869 4131
rect 1869 4097 1903 4131
rect 1903 4097 1912 4131
rect 1860 4088 1912 4097
rect 2688 4088 2740 4140
rect 2872 4131 2924 4140
rect 2872 4097 2906 4131
rect 2906 4097 2924 4131
rect 4252 4156 4304 4208
rect 2872 4088 2924 4097
rect 3976 4088 4028 4140
rect 4712 4131 4764 4140
rect 4712 4097 4721 4131
rect 4721 4097 4755 4131
rect 4755 4097 4764 4131
rect 4712 4088 4764 4097
rect 4436 4020 4488 4072
rect 4620 4063 4672 4072
rect 4620 4029 4629 4063
rect 4629 4029 4663 4063
rect 4663 4029 4672 4063
rect 4620 4020 4672 4029
rect 6552 4156 6604 4208
rect 4988 4088 5040 4140
rect 5356 4088 5408 4140
rect 5816 4088 5868 4140
rect 6460 4131 6512 4140
rect 6460 4097 6469 4131
rect 6469 4097 6503 4131
rect 6503 4097 6512 4131
rect 6460 4088 6512 4097
rect 6644 4131 6696 4140
rect 6644 4097 6653 4131
rect 6653 4097 6687 4131
rect 6687 4097 6696 4131
rect 6644 4088 6696 4097
rect 6736 4131 6788 4140
rect 6736 4097 6745 4131
rect 6745 4097 6779 4131
rect 6779 4097 6788 4131
rect 7748 4224 7800 4276
rect 8024 4224 8076 4276
rect 8208 4224 8260 4276
rect 6736 4088 6788 4097
rect 5908 4020 5960 4072
rect 6184 4020 6236 4072
rect 6552 4020 6604 4072
rect 6920 4063 6972 4072
rect 6920 4029 6929 4063
rect 6929 4029 6963 4063
rect 6963 4029 6972 4063
rect 6920 4020 6972 4029
rect 7748 4088 7800 4140
rect 7840 4088 7892 4140
rect 8208 4088 8260 4140
rect 10508 4224 10560 4276
rect 10876 4224 10928 4276
rect 11704 4224 11756 4276
rect 13176 4224 13228 4276
rect 10692 4156 10744 4208
rect 17592 4156 17644 4208
rect 19524 4156 19576 4208
rect 9128 4088 9180 4140
rect 10784 4088 10836 4140
rect 11520 4131 11572 4140
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 9404 4020 9456 4072
rect 9956 4020 10008 4072
rect 4252 3952 4304 4004
rect 4804 3952 4856 4004
rect 5264 3952 5316 4004
rect 6644 3952 6696 4004
rect 7196 3952 7248 4004
rect 2872 3884 2924 3936
rect 3332 3884 3384 3936
rect 4068 3884 4120 3936
rect 6368 3884 6420 3936
rect 6828 3884 6880 3936
rect 6920 3884 6972 3936
rect 7564 3884 7616 3936
rect 7840 3952 7892 4004
rect 9496 3952 9548 4004
rect 9220 3884 9272 3936
rect 10876 4020 10928 4072
rect 10324 3952 10376 4004
rect 10692 3952 10744 4004
rect 11244 3952 11296 4004
rect 11704 3952 11756 4004
rect 10416 3884 10468 3936
rect 10968 3884 11020 3936
rect 11980 4088 12032 4140
rect 13820 4088 13872 4140
rect 12440 3952 12492 4004
rect 13268 4020 13320 4072
rect 14924 4088 14976 4140
rect 16764 4088 16816 4140
rect 18144 4088 18196 4140
rect 16212 4020 16264 4072
rect 18052 4020 18104 4072
rect 19340 4088 19392 4140
rect 20444 4088 20496 4140
rect 23480 4224 23532 4276
rect 23756 4224 23808 4276
rect 24400 4224 24452 4276
rect 26148 4224 26200 4276
rect 26884 4224 26936 4276
rect 22100 4156 22152 4208
rect 22928 4156 22980 4208
rect 26240 4199 26292 4208
rect 26240 4165 26249 4199
rect 26249 4165 26283 4199
rect 26283 4165 26292 4199
rect 26240 4156 26292 4165
rect 26792 4156 26844 4208
rect 19432 4020 19484 4072
rect 19524 4020 19576 4072
rect 21732 4088 21784 4140
rect 22376 4088 22428 4140
rect 13360 3952 13412 4004
rect 14096 3952 14148 4004
rect 15752 3952 15804 4004
rect 18604 3952 18656 4004
rect 12992 3884 13044 3936
rect 13636 3884 13688 3936
rect 16212 3884 16264 3936
rect 16396 3884 16448 3936
rect 20444 3952 20496 4004
rect 22100 4020 22152 4072
rect 22284 4020 22336 4072
rect 22560 4088 22612 4140
rect 23020 4088 23072 4140
rect 24584 4131 24636 4140
rect 24584 4097 24593 4131
rect 24593 4097 24627 4131
rect 24627 4097 24636 4131
rect 24584 4088 24636 4097
rect 24768 4088 24820 4140
rect 26332 4088 26384 4140
rect 23756 4020 23808 4072
rect 20260 3884 20312 3936
rect 20536 3884 20588 3936
rect 24860 3952 24912 4004
rect 27528 3952 27580 4004
rect 25412 3884 25464 3936
rect 25872 3884 25924 3936
rect 5442 3782 5494 3834
rect 5506 3782 5558 3834
rect 5570 3782 5622 3834
rect 5634 3782 5686 3834
rect 5698 3782 5750 3834
rect 14428 3782 14480 3834
rect 14492 3782 14544 3834
rect 14556 3782 14608 3834
rect 14620 3782 14672 3834
rect 14684 3782 14736 3834
rect 23413 3782 23465 3834
rect 23477 3782 23529 3834
rect 23541 3782 23593 3834
rect 23605 3782 23657 3834
rect 23669 3782 23721 3834
rect 2964 3680 3016 3732
rect 3240 3680 3292 3732
rect 4344 3680 4396 3732
rect 4436 3680 4488 3732
rect 6920 3680 6972 3732
rect 7288 3723 7340 3732
rect 7288 3689 7297 3723
rect 7297 3689 7331 3723
rect 7331 3689 7340 3723
rect 7288 3680 7340 3689
rect 7472 3723 7524 3732
rect 7472 3689 7481 3723
rect 7481 3689 7515 3723
rect 7515 3689 7524 3723
rect 7472 3680 7524 3689
rect 7748 3680 7800 3732
rect 8484 3612 8536 3664
rect 8760 3612 8812 3664
rect 1216 3544 1268 3596
rect 2964 3544 3016 3596
rect 2780 3476 2832 3528
rect 3700 3408 3752 3460
rect 4252 3519 4304 3528
rect 4252 3485 4261 3519
rect 4261 3485 4295 3519
rect 4295 3485 4304 3519
rect 4252 3476 4304 3485
rect 4804 3544 4856 3596
rect 5540 3587 5592 3596
rect 5540 3553 5549 3587
rect 5549 3553 5583 3587
rect 5583 3553 5592 3587
rect 5540 3544 5592 3553
rect 7840 3544 7892 3596
rect 8024 3544 8076 3596
rect 4896 3521 4948 3528
rect 4896 3487 4905 3521
rect 4905 3487 4939 3521
rect 4939 3487 4948 3521
rect 4896 3476 4948 3487
rect 5816 3476 5868 3528
rect 6920 3476 6972 3528
rect 1768 3383 1820 3392
rect 1768 3349 1777 3383
rect 1777 3349 1811 3383
rect 1811 3349 1820 3383
rect 1768 3340 1820 3349
rect 2504 3340 2556 3392
rect 2872 3340 2924 3392
rect 2964 3340 3016 3392
rect 3424 3340 3476 3392
rect 3976 3340 4028 3392
rect 5264 3408 5316 3460
rect 5908 3383 5960 3392
rect 5908 3349 5917 3383
rect 5917 3349 5951 3383
rect 5951 3349 5960 3383
rect 5908 3340 5960 3349
rect 6460 3340 6512 3392
rect 6736 3408 6788 3460
rect 7288 3519 7340 3528
rect 7288 3485 7297 3519
rect 7297 3485 7331 3519
rect 7331 3485 7340 3519
rect 7288 3476 7340 3485
rect 7564 3408 7616 3460
rect 9496 3476 9548 3528
rect 9956 3612 10008 3664
rect 10968 3680 11020 3732
rect 11428 3680 11480 3732
rect 16120 3680 16172 3732
rect 17500 3680 17552 3732
rect 20904 3680 20956 3732
rect 21088 3723 21140 3732
rect 21088 3689 21097 3723
rect 21097 3689 21131 3723
rect 21131 3689 21140 3723
rect 21088 3680 21140 3689
rect 21272 3723 21324 3732
rect 21272 3689 21281 3723
rect 21281 3689 21315 3723
rect 21315 3689 21324 3723
rect 21272 3680 21324 3689
rect 12808 3655 12860 3664
rect 11612 3544 11664 3596
rect 12808 3621 12817 3655
rect 12817 3621 12851 3655
rect 12851 3621 12860 3655
rect 12808 3612 12860 3621
rect 15108 3612 15160 3664
rect 17040 3612 17092 3664
rect 17132 3612 17184 3664
rect 17960 3612 18012 3664
rect 10600 3476 10652 3528
rect 11336 3476 11388 3528
rect 11428 3519 11480 3528
rect 11428 3485 11437 3519
rect 11437 3485 11471 3519
rect 11471 3485 11480 3519
rect 11428 3476 11480 3485
rect 11888 3476 11940 3528
rect 12440 3519 12492 3528
rect 12440 3485 12449 3519
rect 12449 3485 12483 3519
rect 12483 3485 12492 3519
rect 18144 3544 18196 3596
rect 18604 3544 18656 3596
rect 23112 3680 23164 3732
rect 25872 3680 25924 3732
rect 26148 3723 26200 3732
rect 26148 3689 26157 3723
rect 26157 3689 26191 3723
rect 26191 3689 26200 3723
rect 26148 3680 26200 3689
rect 21456 3612 21508 3664
rect 25596 3612 25648 3664
rect 26608 3612 26660 3664
rect 12440 3476 12492 3485
rect 13268 3519 13320 3528
rect 13268 3485 13277 3519
rect 13277 3485 13311 3519
rect 13311 3485 13320 3519
rect 13268 3476 13320 3485
rect 14188 3476 14240 3528
rect 14372 3519 14424 3528
rect 14372 3485 14406 3519
rect 14406 3485 14424 3519
rect 14372 3476 14424 3485
rect 16488 3476 16540 3528
rect 17408 3476 17460 3528
rect 18696 3476 18748 3528
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 9680 3408 9732 3460
rect 10876 3408 10928 3460
rect 11980 3408 12032 3460
rect 8392 3340 8444 3392
rect 11888 3340 11940 3392
rect 15016 3408 15068 3460
rect 19340 3408 19392 3460
rect 20260 3519 20312 3528
rect 20260 3485 20269 3519
rect 20269 3485 20303 3519
rect 20303 3485 20312 3519
rect 20260 3476 20312 3485
rect 21732 3519 21784 3528
rect 21732 3485 21741 3519
rect 21741 3485 21775 3519
rect 21775 3485 21784 3519
rect 21732 3476 21784 3485
rect 22468 3408 22520 3460
rect 23112 3476 23164 3528
rect 23296 3476 23348 3528
rect 24584 3519 24636 3528
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 24768 3476 24820 3528
rect 27160 3476 27212 3528
rect 28724 3476 28776 3528
rect 25964 3451 26016 3460
rect 25964 3417 25973 3451
rect 25973 3417 26007 3451
rect 26007 3417 26016 3451
rect 25964 3408 26016 3417
rect 26424 3408 26476 3460
rect 13544 3340 13596 3392
rect 15844 3340 15896 3392
rect 16488 3340 16540 3392
rect 17960 3340 18012 3392
rect 18788 3340 18840 3392
rect 20260 3340 20312 3392
rect 20996 3340 21048 3392
rect 22376 3340 22428 3392
rect 23296 3340 23348 3392
rect 24400 3383 24452 3392
rect 24400 3349 24409 3383
rect 24409 3349 24443 3383
rect 24443 3349 24452 3383
rect 24400 3340 24452 3349
rect 24768 3383 24820 3392
rect 24768 3349 24777 3383
rect 24777 3349 24811 3383
rect 24811 3349 24820 3383
rect 24768 3340 24820 3349
rect 25320 3340 25372 3392
rect 26884 3340 26936 3392
rect 9935 3238 9987 3290
rect 9999 3238 10051 3290
rect 10063 3238 10115 3290
rect 10127 3238 10179 3290
rect 10191 3238 10243 3290
rect 18920 3238 18972 3290
rect 18984 3238 19036 3290
rect 19048 3238 19100 3290
rect 19112 3238 19164 3290
rect 19176 3238 19228 3290
rect 4804 3136 4856 3188
rect 5540 3136 5592 3188
rect 6184 3136 6236 3188
rect 2688 3068 2740 3120
rect 1768 3043 1820 3052
rect 1768 3009 1802 3043
rect 1802 3009 1820 3043
rect 1768 3000 1820 3009
rect 2320 3000 2372 3052
rect 3240 3000 3292 3052
rect 5080 3068 5132 3120
rect 5264 3068 5316 3120
rect 5448 3111 5500 3120
rect 5448 3077 5457 3111
rect 5457 3077 5491 3111
rect 5491 3077 5500 3111
rect 5448 3068 5500 3077
rect 3608 3043 3660 3052
rect 3608 3009 3642 3043
rect 3642 3009 3660 3043
rect 3608 3000 3660 3009
rect 2596 2864 2648 2916
rect 3332 2864 3384 2916
rect 4620 3000 4672 3052
rect 6276 3000 6328 3052
rect 5080 2932 5132 2984
rect 6460 3000 6512 3052
rect 6920 3136 6972 3188
rect 7196 3136 7248 3188
rect 7288 3136 7340 3188
rect 7380 3068 7432 3120
rect 7932 3068 7984 3120
rect 8484 3111 8536 3120
rect 8484 3077 8518 3111
rect 8518 3077 8536 3111
rect 8484 3068 8536 3077
rect 8208 3043 8260 3052
rect 8208 3009 8217 3043
rect 8217 3009 8251 3043
rect 8251 3009 8260 3043
rect 8208 3000 8260 3009
rect 9680 3136 9732 3188
rect 10876 3136 10928 3188
rect 10508 3068 10560 3120
rect 10600 3000 10652 3052
rect 12532 3136 12584 3188
rect 13268 3136 13320 3188
rect 14280 3136 14332 3188
rect 15108 3136 15160 3188
rect 15292 3136 15344 3188
rect 10692 2932 10744 2984
rect 12256 3068 12308 3120
rect 12624 3068 12676 3120
rect 15476 3068 15528 3120
rect 12072 3000 12124 3052
rect 13084 3000 13136 3052
rect 16948 3136 17000 3188
rect 18144 3136 18196 3188
rect 18420 3136 18472 3188
rect 20076 3136 20128 3188
rect 16672 3068 16724 3120
rect 20628 3111 20680 3120
rect 20628 3077 20637 3111
rect 20637 3077 20671 3111
rect 20671 3077 20680 3111
rect 20628 3068 20680 3077
rect 20996 3068 21048 3120
rect 16488 3000 16540 3052
rect 13360 2975 13412 2984
rect 13360 2941 13369 2975
rect 13369 2941 13403 2975
rect 13403 2941 13412 2975
rect 13360 2932 13412 2941
rect 15936 2932 15988 2984
rect 17224 3000 17276 3052
rect 18144 2932 18196 2984
rect 18696 3000 18748 3052
rect 19984 3000 20036 3052
rect 21180 3000 21232 3052
rect 20812 2932 20864 2984
rect 21456 2932 21508 2984
rect 4896 2864 4948 2916
rect 10416 2864 10468 2916
rect 11244 2864 11296 2916
rect 12532 2864 12584 2916
rect 15384 2864 15436 2916
rect 19524 2864 19576 2916
rect 19708 2864 19760 2916
rect 20076 2907 20128 2916
rect 20076 2873 20085 2907
rect 20085 2873 20119 2907
rect 20119 2873 20128 2907
rect 20076 2864 20128 2873
rect 4712 2839 4764 2848
rect 4712 2805 4721 2839
rect 4721 2805 4755 2839
rect 4755 2805 4764 2839
rect 4712 2796 4764 2805
rect 7012 2796 7064 2848
rect 7564 2796 7616 2848
rect 9864 2796 9916 2848
rect 13176 2796 13228 2848
rect 20444 2796 20496 2848
rect 20904 2864 20956 2916
rect 21088 2864 21140 2916
rect 21640 3136 21692 3188
rect 24400 3111 24452 3120
rect 22100 3043 22152 3052
rect 22100 3009 22109 3043
rect 22109 3009 22143 3043
rect 22143 3009 22152 3043
rect 22376 3043 22428 3052
rect 22100 3000 22152 3009
rect 22376 3009 22410 3043
rect 22410 3009 22428 3043
rect 22376 3000 22428 3009
rect 23112 3000 23164 3052
rect 23756 3000 23808 3052
rect 24400 3077 24434 3111
rect 24434 3077 24452 3111
rect 24400 3068 24452 3077
rect 24768 3136 24820 3188
rect 26884 3136 26936 3188
rect 27344 3068 27396 3120
rect 21364 2796 21416 2848
rect 27252 2864 27304 2916
rect 22284 2796 22336 2848
rect 23296 2796 23348 2848
rect 24032 2796 24084 2848
rect 25964 2796 26016 2848
rect 26148 2839 26200 2848
rect 26148 2805 26157 2839
rect 26157 2805 26191 2839
rect 26191 2805 26200 2839
rect 26148 2796 26200 2805
rect 5442 2694 5494 2746
rect 5506 2694 5558 2746
rect 5570 2694 5622 2746
rect 5634 2694 5686 2746
rect 5698 2694 5750 2746
rect 14428 2694 14480 2746
rect 14492 2694 14544 2746
rect 14556 2694 14608 2746
rect 14620 2694 14672 2746
rect 14684 2694 14736 2746
rect 23413 2694 23465 2746
rect 23477 2694 23529 2746
rect 23541 2694 23593 2746
rect 23605 2694 23657 2746
rect 23669 2694 23721 2746
rect 3608 2592 3660 2644
rect 5816 2592 5868 2644
rect 7196 2592 7248 2644
rect 8300 2592 8352 2644
rect 10968 2592 11020 2644
rect 11796 2592 11848 2644
rect 12164 2592 12216 2644
rect 13268 2592 13320 2644
rect 13728 2592 13780 2644
rect 14924 2592 14976 2644
rect 15384 2635 15436 2644
rect 15384 2601 15393 2635
rect 15393 2601 15427 2635
rect 15427 2601 15436 2635
rect 15384 2592 15436 2601
rect 15936 2635 15988 2644
rect 15936 2601 15945 2635
rect 15945 2601 15979 2635
rect 15979 2601 15988 2635
rect 15936 2592 15988 2601
rect 3516 2524 3568 2576
rect 4896 2524 4948 2576
rect 3700 2456 3752 2508
rect 2228 2388 2280 2440
rect 4712 2431 4764 2440
rect 296 2320 348 2372
rect 2136 2295 2188 2304
rect 2136 2261 2145 2295
rect 2145 2261 2179 2295
rect 2179 2261 2188 2295
rect 2136 2252 2188 2261
rect 2228 2252 2280 2304
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 6368 2524 6420 2576
rect 7012 2456 7064 2508
rect 10508 2524 10560 2576
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 5264 2320 5316 2372
rect 6920 2363 6972 2372
rect 6920 2329 6929 2363
rect 6929 2329 6963 2363
rect 6963 2329 6972 2363
rect 6920 2320 6972 2329
rect 7012 2363 7064 2372
rect 7012 2329 7021 2363
rect 7021 2329 7055 2363
rect 7055 2329 7064 2363
rect 7012 2320 7064 2329
rect 5908 2252 5960 2304
rect 9864 2388 9916 2440
rect 10600 2388 10652 2440
rect 11152 2524 11204 2576
rect 11336 2524 11388 2576
rect 13360 2456 13412 2508
rect 13912 2456 13964 2508
rect 11888 2388 11940 2440
rect 12440 2388 12492 2440
rect 13268 2388 13320 2440
rect 16120 2431 16172 2440
rect 10968 2320 11020 2372
rect 16120 2397 16129 2431
rect 16129 2397 16163 2431
rect 16163 2397 16172 2431
rect 16120 2388 16172 2397
rect 20076 2592 20128 2644
rect 20904 2592 20956 2644
rect 21732 2592 21784 2644
rect 22192 2635 22244 2644
rect 22192 2601 22201 2635
rect 22201 2601 22235 2635
rect 22235 2601 22244 2635
rect 22192 2592 22244 2601
rect 19248 2524 19300 2576
rect 20628 2524 20680 2576
rect 19892 2456 19944 2508
rect 20076 2456 20128 2508
rect 23020 2524 23072 2576
rect 19616 2388 19668 2440
rect 20812 2388 20864 2440
rect 22652 2431 22704 2440
rect 22652 2397 22661 2431
rect 22661 2397 22695 2431
rect 22695 2397 22704 2431
rect 22652 2388 22704 2397
rect 18236 2320 18288 2372
rect 20720 2320 20772 2372
rect 20996 2320 21048 2372
rect 11060 2252 11112 2304
rect 11888 2295 11940 2304
rect 11888 2261 11897 2295
rect 11897 2261 11931 2295
rect 11931 2261 11940 2295
rect 11888 2252 11940 2261
rect 12164 2252 12216 2304
rect 16764 2252 16816 2304
rect 16856 2295 16908 2304
rect 16856 2261 16865 2295
rect 16865 2261 16899 2295
rect 16899 2261 16908 2295
rect 16856 2252 16908 2261
rect 17316 2252 17368 2304
rect 17868 2252 17920 2304
rect 18420 2252 18472 2304
rect 21272 2295 21324 2304
rect 21272 2261 21281 2295
rect 21281 2261 21315 2295
rect 21315 2261 21324 2295
rect 21272 2252 21324 2261
rect 23296 2456 23348 2508
rect 23940 2456 23992 2508
rect 23204 2388 23256 2440
rect 24308 2388 24360 2440
rect 25136 2431 25188 2440
rect 25136 2397 25145 2431
rect 25145 2397 25179 2431
rect 25179 2397 25188 2431
rect 25136 2388 25188 2397
rect 22192 2252 22244 2304
rect 23388 2252 23440 2304
rect 29000 2320 29052 2372
rect 27252 2295 27304 2304
rect 27252 2261 27261 2295
rect 27261 2261 27295 2295
rect 27295 2261 27304 2295
rect 27252 2252 27304 2261
rect 9935 2150 9987 2202
rect 9999 2150 10051 2202
rect 10063 2150 10115 2202
rect 10127 2150 10179 2202
rect 10191 2150 10243 2202
rect 18920 2150 18972 2202
rect 18984 2150 19036 2202
rect 19048 2150 19100 2202
rect 19112 2150 19164 2202
rect 19176 2150 19228 2202
rect 3148 2048 3200 2100
rect 7012 2048 7064 2100
rect 16764 2048 16816 2100
rect 27252 2048 27304 2100
rect 2136 1980 2188 2032
rect 9036 1980 9088 2032
rect 16856 1980 16908 2032
rect 27068 1980 27120 2032
rect 3792 1912 3844 1964
rect 11888 1912 11940 1964
rect 16764 1912 16816 1964
rect 17132 1912 17184 1964
rect 19524 1912 19576 1964
rect 20352 1912 20404 1964
rect 21272 1912 21324 1964
rect 24124 1912 24176 1964
rect 21088 1436 21140 1488
rect 23388 1436 23440 1488
rect 21640 1368 21692 1420
rect 23020 1368 23072 1420
rect 18788 1028 18840 1080
rect 19248 1028 19300 1080
<< metal2 >>
rect 5442 28860 5750 28880
rect 5442 28858 5448 28860
rect 5504 28858 5528 28860
rect 5584 28858 5608 28860
rect 5664 28858 5688 28860
rect 5744 28858 5750 28860
rect 5504 28806 5506 28858
rect 5686 28806 5688 28858
rect 5442 28804 5448 28806
rect 5504 28804 5528 28806
rect 5584 28804 5608 28806
rect 5664 28804 5688 28806
rect 5744 28804 5750 28806
rect 5442 28784 5750 28804
rect 14428 28860 14736 28880
rect 14428 28858 14434 28860
rect 14490 28858 14514 28860
rect 14570 28858 14594 28860
rect 14650 28858 14674 28860
rect 14730 28858 14736 28860
rect 14490 28806 14492 28858
rect 14672 28806 14674 28858
rect 14428 28804 14434 28806
rect 14490 28804 14514 28806
rect 14570 28804 14594 28806
rect 14650 28804 14674 28806
rect 14730 28804 14736 28806
rect 14428 28784 14736 28804
rect 23413 28860 23721 28880
rect 23413 28858 23419 28860
rect 23475 28858 23499 28860
rect 23555 28858 23579 28860
rect 23635 28858 23659 28860
rect 23715 28858 23721 28860
rect 23475 28806 23477 28858
rect 23657 28806 23659 28858
rect 23413 28804 23419 28806
rect 23475 28804 23499 28806
rect 23555 28804 23579 28806
rect 23635 28804 23659 28806
rect 23715 28804 23721 28806
rect 23413 28784 23721 28804
rect 12808 28756 12860 28762
rect 12808 28698 12860 28704
rect 15752 28756 15804 28762
rect 15752 28698 15804 28704
rect 16672 28756 16724 28762
rect 16672 28698 16724 28704
rect 9128 28688 9180 28694
rect 9128 28630 9180 28636
rect 8300 28552 8352 28558
rect 8300 28494 8352 28500
rect 8392 28552 8444 28558
rect 8392 28494 8444 28500
rect 4344 28416 4396 28422
rect 4344 28358 4396 28364
rect 7104 28416 7156 28422
rect 7104 28358 7156 28364
rect 7472 28416 7524 28422
rect 7472 28358 7524 28364
rect 4356 28218 4384 28358
rect 4344 28212 4396 28218
rect 4344 28154 4396 28160
rect 5908 28212 5960 28218
rect 5908 28154 5960 28160
rect 4252 28144 4304 28150
rect 4252 28086 4304 28092
rect 3884 27872 3936 27878
rect 3884 27814 3936 27820
rect 2596 27464 2648 27470
rect 2596 27406 2648 27412
rect 3700 27464 3752 27470
rect 3700 27406 3752 27412
rect 2504 27328 2556 27334
rect 2504 27270 2556 27276
rect 1400 26988 1452 26994
rect 1400 26930 1452 26936
rect 1412 25922 1440 26930
rect 1860 26920 1912 26926
rect 1860 26862 1912 26868
rect 1676 26784 1728 26790
rect 1676 26726 1728 26732
rect 1584 26512 1636 26518
rect 1584 26454 1636 26460
rect 1320 25894 1440 25922
rect 1320 25702 1348 25894
rect 1400 25832 1452 25838
rect 1596 25786 1624 26454
rect 1400 25774 1452 25780
rect 1308 25696 1360 25702
rect 1308 25638 1360 25644
rect 1308 24744 1360 24750
rect 1308 24686 1360 24692
rect 204 24404 256 24410
rect 204 24346 256 24352
rect 216 22094 244 24346
rect 216 22066 612 22094
rect 110 3496 166 3505
rect 110 3431 166 3440
rect 124 800 152 3431
rect 296 2372 348 2378
rect 296 2314 348 2320
rect 308 800 336 2314
rect 584 800 612 22066
rect 1216 21072 1268 21078
rect 1216 21014 1268 21020
rect 1124 19712 1176 19718
rect 1124 19654 1176 19660
rect 1032 16720 1084 16726
rect 1032 16662 1084 16668
rect 1044 11762 1072 16662
rect 1032 11756 1084 11762
rect 1032 11698 1084 11704
rect 848 4140 900 4146
rect 848 4082 900 4088
rect 860 800 888 4082
rect 1136 3641 1164 19654
rect 1122 3632 1178 3641
rect 1228 3602 1256 21014
rect 1122 3567 1178 3576
rect 1216 3596 1268 3602
rect 1216 3538 1268 3544
rect 1320 2825 1348 24686
rect 1412 24274 1440 25774
rect 1504 25758 1624 25786
rect 1400 24268 1452 24274
rect 1400 24210 1452 24216
rect 1504 20398 1532 25758
rect 1584 25696 1636 25702
rect 1584 25638 1636 25644
rect 1492 20392 1544 20398
rect 1492 20334 1544 20340
rect 1492 20256 1544 20262
rect 1492 20198 1544 20204
rect 1400 18760 1452 18766
rect 1400 18702 1452 18708
rect 1412 16726 1440 18702
rect 1400 16720 1452 16726
rect 1400 16662 1452 16668
rect 1400 16584 1452 16590
rect 1400 16526 1452 16532
rect 1412 15570 1440 16526
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1400 15156 1452 15162
rect 1400 15098 1452 15104
rect 1412 10470 1440 15098
rect 1400 10464 1452 10470
rect 1400 10406 1452 10412
rect 1504 10146 1532 20198
rect 1412 10118 1532 10146
rect 1412 6361 1440 10118
rect 1596 10010 1624 25638
rect 1688 22094 1716 26726
rect 1872 25838 1900 26862
rect 1860 25832 1912 25838
rect 1860 25774 1912 25780
rect 2412 24812 2464 24818
rect 2412 24754 2464 24760
rect 2424 24682 2452 24754
rect 2412 24676 2464 24682
rect 2412 24618 2464 24624
rect 1952 24608 2004 24614
rect 1952 24550 2004 24556
rect 1688 22066 1808 22094
rect 1676 20392 1728 20398
rect 1676 20334 1728 20340
rect 1688 15162 1716 20334
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1676 14340 1728 14346
rect 1676 14282 1728 14288
rect 1688 14074 1716 14282
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1688 13326 1716 13806
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1676 12164 1728 12170
rect 1676 12106 1728 12112
rect 1688 11898 1716 12106
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1504 9982 1624 10010
rect 1398 6352 1454 6361
rect 1398 6287 1454 6296
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1412 4622 1440 6190
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 1504 4146 1532 9982
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1596 9722 1624 9862
rect 1584 9716 1636 9722
rect 1584 9658 1636 9664
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1596 7886 1624 9454
rect 1688 8945 1716 11698
rect 1780 8974 1808 22066
rect 1860 20052 1912 20058
rect 1860 19994 1912 20000
rect 1872 19514 1900 19994
rect 1860 19508 1912 19514
rect 1860 19450 1912 19456
rect 1858 18864 1914 18873
rect 1858 18799 1914 18808
rect 1872 18766 1900 18799
rect 1860 18760 1912 18766
rect 1860 18702 1912 18708
rect 1860 18624 1912 18630
rect 1860 18566 1912 18572
rect 1872 15609 1900 18566
rect 1964 18426 1992 24550
rect 2136 23724 2188 23730
rect 2136 23666 2188 23672
rect 2044 22976 2096 22982
rect 2044 22918 2096 22924
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1952 18216 2004 18222
rect 1952 18158 2004 18164
rect 1964 17678 1992 18158
rect 1952 17672 2004 17678
rect 1952 17614 2004 17620
rect 1964 17134 1992 17614
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 1964 16590 1992 17070
rect 1952 16584 2004 16590
rect 1952 16526 2004 16532
rect 1964 16182 1992 16526
rect 1952 16176 2004 16182
rect 1952 16118 2004 16124
rect 1858 15600 1914 15609
rect 1858 15535 1914 15544
rect 2056 15450 2084 22918
rect 1860 15428 1912 15434
rect 1860 15370 1912 15376
rect 1964 15422 2084 15450
rect 1872 15162 1900 15370
rect 1860 15156 1912 15162
rect 1860 15098 1912 15104
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1872 12442 1900 13874
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1872 11082 1900 11494
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 1768 8968 1820 8974
rect 1674 8936 1730 8945
rect 1768 8910 1820 8916
rect 1674 8871 1730 8880
rect 1860 8288 1912 8294
rect 1860 8230 1912 8236
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1596 6322 1624 7822
rect 1872 7818 1900 8230
rect 1860 7812 1912 7818
rect 1860 7754 1912 7760
rect 1964 7426 1992 15422
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 2056 13870 2084 14350
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 2056 12186 2084 12786
rect 2148 12306 2176 23666
rect 2412 22432 2464 22438
rect 2516 22409 2544 27270
rect 2608 27130 2636 27406
rect 3712 27334 3740 27406
rect 3056 27328 3108 27334
rect 3056 27270 3108 27276
rect 3700 27328 3752 27334
rect 3700 27270 3752 27276
rect 2596 27124 2648 27130
rect 2596 27066 2648 27072
rect 2872 26988 2924 26994
rect 2872 26930 2924 26936
rect 2884 26790 2912 26930
rect 2872 26784 2924 26790
rect 2872 26726 2924 26732
rect 2688 26308 2740 26314
rect 2688 26250 2740 26256
rect 2700 23089 2728 26250
rect 2780 23520 2832 23526
rect 2780 23462 2832 23468
rect 2686 23080 2742 23089
rect 2686 23015 2742 23024
rect 2596 22976 2648 22982
rect 2596 22918 2648 22924
rect 2412 22374 2464 22380
rect 2502 22400 2558 22409
rect 2424 22094 2452 22374
rect 2502 22335 2558 22344
rect 2424 22066 2544 22094
rect 2320 21888 2372 21894
rect 2372 21836 2452 21842
rect 2320 21830 2452 21836
rect 2332 21814 2452 21830
rect 2228 20936 2280 20942
rect 2228 20878 2280 20884
rect 2240 20777 2268 20878
rect 2424 20806 2452 21814
rect 2320 20800 2372 20806
rect 2226 20768 2282 20777
rect 2320 20742 2372 20748
rect 2412 20800 2464 20806
rect 2412 20742 2464 20748
rect 2226 20703 2282 20712
rect 2228 20392 2280 20398
rect 2228 20334 2280 20340
rect 2240 18630 2268 20334
rect 2228 18624 2280 18630
rect 2228 18566 2280 18572
rect 2228 18420 2280 18426
rect 2228 18362 2280 18368
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 2056 12170 2176 12186
rect 2056 12164 2188 12170
rect 2056 12158 2136 12164
rect 2136 12106 2188 12112
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 2056 10810 2084 11698
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 2148 10674 2176 12106
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2056 7546 2084 8434
rect 2148 8362 2176 10610
rect 2240 10606 2268 18362
rect 2332 15450 2360 20742
rect 2516 20074 2544 22066
rect 2608 21865 2636 22918
rect 2688 21888 2740 21894
rect 2594 21856 2650 21865
rect 2688 21830 2740 21836
rect 2594 21791 2650 21800
rect 2596 21344 2648 21350
rect 2596 21286 2648 21292
rect 2608 20233 2636 21286
rect 2700 21049 2728 21830
rect 2686 21040 2742 21049
rect 2686 20975 2742 20984
rect 2688 20460 2740 20466
rect 2688 20402 2740 20408
rect 2594 20224 2650 20233
rect 2594 20159 2650 20168
rect 2516 20046 2636 20074
rect 2412 19984 2464 19990
rect 2412 19926 2464 19932
rect 2502 19952 2558 19961
rect 2424 16266 2452 19926
rect 2502 19887 2558 19896
rect 2516 19378 2544 19887
rect 2504 19372 2556 19378
rect 2504 19314 2556 19320
rect 2608 19281 2636 20046
rect 2700 19417 2728 20402
rect 2686 19408 2742 19417
rect 2686 19343 2742 19352
rect 2594 19272 2650 19281
rect 2594 19207 2650 19216
rect 2688 19236 2740 19242
rect 2688 19178 2740 19184
rect 2596 19168 2648 19174
rect 2700 19145 2728 19178
rect 2596 19110 2648 19116
rect 2686 19136 2742 19145
rect 2504 18284 2556 18290
rect 2504 18226 2556 18232
rect 2516 17338 2544 18226
rect 2608 17882 2636 19110
rect 2686 19071 2742 19080
rect 2688 18760 2740 18766
rect 2686 18728 2688 18737
rect 2740 18728 2742 18737
rect 2686 18663 2742 18672
rect 2596 17876 2648 17882
rect 2596 17818 2648 17824
rect 2504 17332 2556 17338
rect 2504 17274 2556 17280
rect 2792 16289 2820 23462
rect 2884 22094 2912 26726
rect 3068 26353 3096 27270
rect 3424 26512 3476 26518
rect 3424 26454 3476 26460
rect 3054 26344 3110 26353
rect 3054 26279 3110 26288
rect 2964 26240 3016 26246
rect 2964 26182 3016 26188
rect 2976 25498 3004 26182
rect 2964 25492 3016 25498
rect 2964 25434 3016 25440
rect 3240 25288 3292 25294
rect 3240 25230 3292 25236
rect 3056 25152 3108 25158
rect 3056 25094 3108 25100
rect 2964 24608 3016 24614
rect 2964 24550 3016 24556
rect 2976 24342 3004 24550
rect 2964 24336 3016 24342
rect 2964 24278 3016 24284
rect 2964 24064 3016 24070
rect 2964 24006 3016 24012
rect 2976 23118 3004 24006
rect 2964 23112 3016 23118
rect 2964 23054 3016 23060
rect 2964 22976 3016 22982
rect 2964 22918 3016 22924
rect 2976 22778 3004 22918
rect 2964 22772 3016 22778
rect 2964 22714 3016 22720
rect 2884 22066 3004 22094
rect 2870 21992 2926 22001
rect 2870 21927 2926 21936
rect 2884 21690 2912 21927
rect 2872 21684 2924 21690
rect 2872 21626 2924 21632
rect 2872 20868 2924 20874
rect 2872 20810 2924 20816
rect 2884 20505 2912 20810
rect 2870 20496 2926 20505
rect 2870 20431 2926 20440
rect 2872 20256 2924 20262
rect 2872 20198 2924 20204
rect 2884 16658 2912 20198
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2778 16280 2834 16289
rect 2424 16238 2636 16266
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 2424 15745 2452 15846
rect 2410 15736 2466 15745
rect 2410 15671 2466 15680
rect 2516 15570 2544 16050
rect 2504 15564 2556 15570
rect 2504 15506 2556 15512
rect 2332 15422 2544 15450
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2228 10600 2280 10606
rect 2228 10542 2280 10548
rect 2228 9920 2280 9926
rect 2228 9862 2280 9868
rect 2240 9654 2268 9862
rect 2228 9648 2280 9654
rect 2228 9590 2280 9596
rect 2226 8936 2282 8945
rect 2332 8906 2360 15302
rect 2516 15076 2544 15422
rect 2608 15366 2636 16238
rect 2778 16215 2834 16224
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 2792 15706 2820 16050
rect 2872 15904 2924 15910
rect 2872 15846 2924 15852
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2686 15464 2742 15473
rect 2686 15399 2742 15408
rect 2596 15360 2648 15366
rect 2596 15302 2648 15308
rect 2700 15076 2728 15399
rect 2884 15094 2912 15846
rect 2424 15048 2544 15076
rect 2608 15048 2728 15076
rect 2872 15088 2924 15094
rect 2424 11830 2452 15048
rect 2504 13252 2556 13258
rect 2504 13194 2556 13200
rect 2516 12442 2544 13194
rect 2504 12436 2556 12442
rect 2504 12378 2556 12384
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 2412 11824 2464 11830
rect 2412 11766 2464 11772
rect 2516 11676 2544 12242
rect 2424 11648 2544 11676
rect 2226 8871 2282 8880
rect 2320 8900 2372 8906
rect 2136 8356 2188 8362
rect 2136 8298 2188 8304
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 1964 7398 2084 7426
rect 2148 7410 2176 8298
rect 1952 6724 2004 6730
rect 1952 6666 2004 6672
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1964 5914 1992 6666
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1676 4548 1728 4554
rect 1676 4490 1728 4496
rect 1688 4282 1716 4490
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 1872 4146 1900 4966
rect 2056 4321 2084 7398
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 2042 4312 2098 4321
rect 2042 4247 2098 4256
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1768 3392 1820 3398
rect 1768 3334 1820 3340
rect 1780 3058 1808 3334
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 1306 2816 1362 2825
rect 1306 2751 1362 2760
rect 2240 2446 2268 8871
rect 2320 8842 2372 8848
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2332 6322 2360 6598
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2424 6202 2452 11648
rect 2608 10418 2636 15048
rect 2872 15030 2924 15036
rect 2688 14884 2740 14890
rect 2688 14826 2740 14832
rect 2700 12753 2728 14826
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2884 13938 2912 14214
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2872 13728 2924 13734
rect 2976 13705 3004 22066
rect 3068 19802 3096 25094
rect 3148 24676 3200 24682
rect 3148 24618 3200 24624
rect 3160 24274 3188 24618
rect 3252 24410 3280 25230
rect 3332 25220 3384 25226
rect 3332 25162 3384 25168
rect 3240 24404 3292 24410
rect 3240 24346 3292 24352
rect 3148 24268 3200 24274
rect 3148 24210 3200 24216
rect 3240 24132 3292 24138
rect 3240 24074 3292 24080
rect 3252 23594 3280 24074
rect 3240 23588 3292 23594
rect 3240 23530 3292 23536
rect 3148 23112 3200 23118
rect 3148 23054 3200 23060
rect 3160 22166 3188 23054
rect 3148 22160 3200 22166
rect 3148 22102 3200 22108
rect 3160 21622 3188 22102
rect 3240 21888 3292 21894
rect 3240 21830 3292 21836
rect 3252 21690 3280 21830
rect 3240 21684 3292 21690
rect 3240 21626 3292 21632
rect 3148 21616 3200 21622
rect 3148 21558 3200 21564
rect 3238 21584 3294 21593
rect 3238 21519 3294 21528
rect 3252 21418 3280 21519
rect 3240 21412 3292 21418
rect 3240 21354 3292 21360
rect 3148 20936 3200 20942
rect 3146 20904 3148 20913
rect 3200 20904 3202 20913
rect 3146 20839 3202 20848
rect 3240 20800 3292 20806
rect 3238 20768 3240 20777
rect 3292 20768 3294 20777
rect 3238 20703 3294 20712
rect 3068 19774 3280 19802
rect 3056 19712 3108 19718
rect 3056 19654 3108 19660
rect 2872 13670 2924 13676
rect 2962 13696 3018 13705
rect 2686 12744 2742 12753
rect 2686 12679 2742 12688
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2700 12238 2728 12582
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2792 11642 2820 11698
rect 2700 11614 2820 11642
rect 2700 11286 2728 11614
rect 2688 11280 2740 11286
rect 2688 11222 2740 11228
rect 2516 10390 2636 10418
rect 2516 6882 2544 10390
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2608 9042 2636 10202
rect 2700 9042 2728 11222
rect 2884 10266 2912 13670
rect 2962 13631 3018 13640
rect 2964 12368 3016 12374
rect 2964 12310 3016 12316
rect 2976 12073 3004 12310
rect 2962 12064 3018 12073
rect 2962 11999 3018 12008
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 3068 10146 3096 19654
rect 3148 19372 3200 19378
rect 3148 19314 3200 19320
rect 3160 19009 3188 19314
rect 3146 19000 3202 19009
rect 3146 18935 3202 18944
rect 3146 18864 3202 18873
rect 3146 18799 3148 18808
rect 3200 18799 3202 18808
rect 3148 18770 3200 18776
rect 3148 14340 3200 14346
rect 3148 14282 3200 14288
rect 3160 14249 3188 14282
rect 3146 14240 3202 14249
rect 3146 14175 3202 14184
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 2792 10118 3096 10146
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2792 8922 2820 10118
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 3054 10024 3110 10033
rect 2700 8894 2820 8922
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2608 8566 2636 8774
rect 2596 8560 2648 8566
rect 2596 8502 2648 8508
rect 2700 7546 2728 8894
rect 2884 8634 2912 9998
rect 3054 9959 3110 9968
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2976 8974 3004 9318
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2780 8016 2832 8022
rect 2780 7958 2832 7964
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2792 7410 2820 7958
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2608 7002 2636 7278
rect 2780 7268 2832 7274
rect 2780 7210 2832 7216
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 2516 6854 2636 6882
rect 2332 6174 2452 6202
rect 2332 3058 2360 6174
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 2228 2304 2280 2310
rect 2228 2246 2280 2252
rect 2148 2038 2176 2246
rect 2136 2032 2188 2038
rect 2136 1974 2188 1980
rect 2240 800 2268 2246
rect 2516 800 2544 3334
rect 2608 2922 2636 6854
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 2700 4622 2728 6190
rect 2792 6118 2820 7210
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2884 5930 2912 7278
rect 2964 6996 3016 7002
rect 2964 6938 3016 6944
rect 2792 5902 2912 5930
rect 2792 5710 2820 5902
rect 2976 5846 3004 6938
rect 3068 6905 3096 9959
rect 3054 6896 3110 6905
rect 3054 6831 3110 6840
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 2964 5840 3016 5846
rect 2964 5782 3016 5788
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2778 5400 2834 5409
rect 2778 5335 2834 5344
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2700 4146 2728 4558
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2700 3126 2728 4082
rect 2792 3534 2820 5335
rect 2884 4146 2912 5782
rect 3068 5778 3096 6054
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 2962 5672 3018 5681
rect 2962 5607 3018 5616
rect 3056 5636 3108 5642
rect 2976 5250 3004 5607
rect 3056 5578 3108 5584
rect 3068 5370 3096 5578
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 2976 5222 3096 5250
rect 2964 4208 3016 4214
rect 2964 4150 3016 4156
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2884 3398 2912 3878
rect 2976 3738 3004 4150
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 2976 3398 3004 3538
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2870 3224 2926 3233
rect 2870 3159 2926 3168
rect 2688 3120 2740 3126
rect 2688 3062 2740 3068
rect 2596 2916 2648 2922
rect 2596 2858 2648 2864
rect 2884 2774 2912 3159
rect 2792 2746 2912 2774
rect 2792 800 2820 2746
rect 3068 800 3096 5222
rect 3160 2106 3188 14010
rect 3252 13734 3280 19774
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3238 13560 3294 13569
rect 3238 13495 3294 13504
rect 3252 8090 3280 13495
rect 3344 11150 3372 25162
rect 3436 24750 3464 26454
rect 3516 26376 3568 26382
rect 3516 26318 3568 26324
rect 3528 24886 3556 26318
rect 3516 24880 3568 24886
rect 3516 24822 3568 24828
rect 3712 24750 3740 27270
rect 3424 24744 3476 24750
rect 3700 24744 3752 24750
rect 3476 24704 3556 24732
rect 3424 24686 3476 24692
rect 3424 24608 3476 24614
rect 3424 24550 3476 24556
rect 3436 23730 3464 24550
rect 3528 24410 3556 24704
rect 3700 24686 3752 24692
rect 3792 24676 3844 24682
rect 3792 24618 3844 24624
rect 3700 24608 3752 24614
rect 3700 24550 3752 24556
rect 3516 24404 3568 24410
rect 3516 24346 3568 24352
rect 3424 23724 3476 23730
rect 3424 23666 3476 23672
rect 3528 22982 3556 24346
rect 3608 23656 3660 23662
rect 3608 23598 3660 23604
rect 3620 23526 3648 23598
rect 3608 23520 3660 23526
rect 3608 23462 3660 23468
rect 3516 22976 3568 22982
rect 3516 22918 3568 22924
rect 3606 22808 3662 22817
rect 3606 22743 3662 22752
rect 3424 22024 3476 22030
rect 3424 21966 3476 21972
rect 3436 18737 3464 21966
rect 3516 21888 3568 21894
rect 3516 21830 3568 21836
rect 3422 18728 3478 18737
rect 3422 18663 3478 18672
rect 3424 18624 3476 18630
rect 3424 18566 3476 18572
rect 3436 17270 3464 18566
rect 3424 17264 3476 17270
rect 3424 17206 3476 17212
rect 3528 17082 3556 21830
rect 3620 21554 3648 22743
rect 3608 21548 3660 21554
rect 3608 21490 3660 21496
rect 3608 20800 3660 20806
rect 3608 20742 3660 20748
rect 3620 20369 3648 20742
rect 3606 20360 3662 20369
rect 3606 20295 3662 20304
rect 3608 20052 3660 20058
rect 3608 19994 3660 20000
rect 3620 19825 3648 19994
rect 3606 19816 3662 19825
rect 3606 19751 3662 19760
rect 3608 19712 3660 19718
rect 3606 19680 3608 19689
rect 3660 19680 3662 19689
rect 3606 19615 3662 19624
rect 3606 19544 3662 19553
rect 3606 19479 3608 19488
rect 3660 19479 3662 19488
rect 3608 19450 3660 19456
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 3620 18970 3648 19314
rect 3608 18964 3660 18970
rect 3608 18906 3660 18912
rect 3620 18358 3648 18906
rect 3608 18352 3660 18358
rect 3608 18294 3660 18300
rect 3620 17746 3648 18294
rect 3608 17740 3660 17746
rect 3608 17682 3660 17688
rect 3608 17604 3660 17610
rect 3608 17546 3660 17552
rect 3436 17054 3556 17082
rect 3436 12889 3464 17054
rect 3620 16794 3648 17546
rect 3608 16788 3660 16794
rect 3608 16730 3660 16736
rect 3608 16652 3660 16658
rect 3608 16594 3660 16600
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 3422 12880 3478 12889
rect 3422 12815 3478 12824
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 3436 12442 3464 12718
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3436 11762 3464 12174
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3344 10674 3372 10950
rect 3436 10742 3464 11698
rect 3528 11234 3556 16050
rect 3620 13025 3648 16594
rect 3606 13016 3662 13025
rect 3606 12951 3662 12960
rect 3608 12912 3660 12918
rect 3608 12854 3660 12860
rect 3620 11898 3648 12854
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3528 11206 3648 11234
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3424 10736 3476 10742
rect 3424 10678 3476 10684
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 3344 10266 3372 10610
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3436 9926 3464 10678
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3252 7410 3280 7686
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3238 6896 3294 6905
rect 3238 6831 3294 6840
rect 3252 5710 3280 6831
rect 3344 6662 3372 9522
rect 3436 8022 3464 9862
rect 3424 8016 3476 8022
rect 3424 7958 3476 7964
rect 3424 7812 3476 7818
rect 3424 7754 3476 7760
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3330 6488 3386 6497
rect 3330 6423 3386 6432
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 3344 3942 3372 6423
rect 3436 5574 3464 7754
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3424 4276 3476 4282
rect 3424 4218 3476 4224
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3252 3058 3280 3674
rect 3436 3482 3464 4218
rect 3344 3454 3464 3482
rect 3344 3233 3372 3454
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3330 3224 3386 3233
rect 3330 3159 3386 3168
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3332 2916 3384 2922
rect 3332 2858 3384 2864
rect 3148 2100 3200 2106
rect 3148 2042 3200 2048
rect 3344 800 3372 2858
rect 3436 1442 3464 3334
rect 3528 2582 3556 11086
rect 3620 6984 3648 11206
rect 3712 7410 3740 24550
rect 3804 24206 3832 24618
rect 3792 24200 3844 24206
rect 3792 24142 3844 24148
rect 3804 23322 3832 24142
rect 3792 23316 3844 23322
rect 3792 23258 3844 23264
rect 3792 22704 3844 22710
rect 3792 22646 3844 22652
rect 3804 20942 3832 22646
rect 3792 20936 3844 20942
rect 3792 20878 3844 20884
rect 3792 20800 3844 20806
rect 3792 20742 3844 20748
rect 3804 15144 3832 20742
rect 3896 18329 3924 27814
rect 4160 27532 4212 27538
rect 4160 27474 4212 27480
rect 4172 27282 4200 27474
rect 4080 27254 4200 27282
rect 4080 27130 4108 27254
rect 4068 27124 4120 27130
rect 4068 27066 4120 27072
rect 4160 27124 4212 27130
rect 4160 27066 4212 27072
rect 4172 26382 4200 27066
rect 4264 27062 4292 28086
rect 4356 27606 4384 28154
rect 5264 28076 5316 28082
rect 5264 28018 5316 28024
rect 4344 27600 4396 27606
rect 4344 27542 4396 27548
rect 4988 27532 5040 27538
rect 4988 27474 5040 27480
rect 4712 27464 4764 27470
rect 4712 27406 4764 27412
rect 4344 27328 4396 27334
rect 4344 27270 4396 27276
rect 4252 27056 4304 27062
rect 4252 26998 4304 27004
rect 4160 26376 4212 26382
rect 4160 26318 4212 26324
rect 4068 26308 4120 26314
rect 4068 26250 4120 26256
rect 4080 25906 4108 26250
rect 4068 25900 4120 25906
rect 4068 25842 4120 25848
rect 4160 25900 4212 25906
rect 4356 25888 4384 27270
rect 4528 26988 4580 26994
rect 4528 26930 4580 26936
rect 4540 26586 4568 26930
rect 4528 26580 4580 26586
rect 4528 26522 4580 26528
rect 4212 25860 4384 25888
rect 4434 25936 4490 25945
rect 4434 25871 4490 25880
rect 4528 25900 4580 25906
rect 4160 25842 4212 25848
rect 4448 25838 4476 25871
rect 4528 25842 4580 25848
rect 4436 25832 4488 25838
rect 4436 25774 4488 25780
rect 4080 25498 4384 25514
rect 4068 25492 4384 25498
rect 4120 25486 4384 25492
rect 4068 25434 4120 25440
rect 4160 25424 4212 25430
rect 4160 25366 4212 25372
rect 3976 24880 4028 24886
rect 3976 24822 4028 24828
rect 3988 24206 4016 24822
rect 4068 24812 4120 24818
rect 4068 24754 4120 24760
rect 3976 24200 4028 24206
rect 3976 24142 4028 24148
rect 4080 24070 4108 24754
rect 4172 24614 4200 25366
rect 4252 25152 4304 25158
rect 4252 25094 4304 25100
rect 4160 24608 4212 24614
rect 4160 24550 4212 24556
rect 4068 24064 4120 24070
rect 4068 24006 4120 24012
rect 4080 23730 4108 24006
rect 4068 23724 4120 23730
rect 4068 23666 4120 23672
rect 3976 22976 4028 22982
rect 3976 22918 4028 22924
rect 3988 22778 4016 22918
rect 3976 22772 4028 22778
rect 3976 22714 4028 22720
rect 4172 22681 4200 24550
rect 4264 24070 4292 25094
rect 4252 24064 4304 24070
rect 4252 24006 4304 24012
rect 4264 23866 4292 24006
rect 4252 23860 4304 23866
rect 4252 23802 4304 23808
rect 4250 23760 4306 23769
rect 4250 23695 4306 23704
rect 4264 23118 4292 23695
rect 4252 23112 4304 23118
rect 4252 23054 4304 23060
rect 4264 22817 4292 23054
rect 4356 22953 4384 25486
rect 4448 23526 4476 25774
rect 4540 25537 4568 25842
rect 4620 25832 4672 25838
rect 4620 25774 4672 25780
rect 4526 25528 4582 25537
rect 4632 25498 4660 25774
rect 4526 25463 4582 25472
rect 4620 25492 4672 25498
rect 4620 25434 4672 25440
rect 4724 25158 4752 27406
rect 4896 26784 4948 26790
rect 4896 26726 4948 26732
rect 4908 26450 4936 26726
rect 4896 26444 4948 26450
rect 4896 26386 4948 26392
rect 4804 26376 4856 26382
rect 4804 26318 4856 26324
rect 4816 26042 4844 26318
rect 4896 26240 4948 26246
rect 4896 26182 4948 26188
rect 4804 26036 4856 26042
rect 4804 25978 4856 25984
rect 4908 25702 4936 26182
rect 4804 25696 4856 25702
rect 4804 25638 4856 25644
rect 4896 25696 4948 25702
rect 4896 25638 4948 25644
rect 4816 25362 4844 25638
rect 4804 25356 4856 25362
rect 4804 25298 4856 25304
rect 4712 25152 4764 25158
rect 4712 25094 4764 25100
rect 4816 24886 4844 25298
rect 4804 24880 4856 24886
rect 4804 24822 4856 24828
rect 4896 24812 4948 24818
rect 4896 24754 4948 24760
rect 4528 24336 4580 24342
rect 4528 24278 4580 24284
rect 4436 23520 4488 23526
rect 4436 23462 4488 23468
rect 4436 23180 4488 23186
rect 4436 23122 4488 23128
rect 4342 22944 4398 22953
rect 4342 22879 4398 22888
rect 4250 22808 4306 22817
rect 4448 22794 4476 23122
rect 4250 22743 4306 22752
rect 4356 22766 4476 22794
rect 4158 22672 4214 22681
rect 4068 22636 4120 22642
rect 4356 22624 4384 22766
rect 4436 22704 4488 22710
rect 4436 22646 4488 22652
rect 4158 22607 4214 22616
rect 4068 22578 4120 22584
rect 4264 22596 4384 22624
rect 4080 22234 4108 22578
rect 4160 22568 4212 22574
rect 4160 22510 4212 22516
rect 4068 22228 4120 22234
rect 4068 22170 4120 22176
rect 3976 22024 4028 22030
rect 3976 21966 4028 21972
rect 3988 21729 4016 21966
rect 3974 21720 4030 21729
rect 4080 21690 4108 22170
rect 4172 21690 4200 22510
rect 4264 22030 4292 22596
rect 4344 22500 4396 22506
rect 4344 22442 4396 22448
rect 4252 22024 4304 22030
rect 4252 21966 4304 21972
rect 3974 21655 4030 21664
rect 4068 21684 4120 21690
rect 4068 21626 4120 21632
rect 4160 21684 4212 21690
rect 4160 21626 4212 21632
rect 4172 21486 4200 21626
rect 4264 21554 4292 21966
rect 4252 21548 4304 21554
rect 4252 21490 4304 21496
rect 4160 21480 4212 21486
rect 4160 21422 4212 21428
rect 3976 21072 4028 21078
rect 3976 21014 4028 21020
rect 3882 18320 3938 18329
rect 3882 18255 3938 18264
rect 3884 18080 3936 18086
rect 3884 18022 3936 18028
rect 3896 17678 3924 18022
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3896 15337 3924 15846
rect 3882 15328 3938 15337
rect 3882 15263 3938 15272
rect 3804 15116 3924 15144
rect 3792 15020 3844 15026
rect 3792 14962 3844 14968
rect 3804 14618 3832 14962
rect 3792 14612 3844 14618
rect 3792 14554 3844 14560
rect 3896 14498 3924 15116
rect 3804 14470 3924 14498
rect 3804 9602 3832 14470
rect 3882 14376 3938 14385
rect 3882 14311 3938 14320
rect 3896 13954 3924 14311
rect 3988 14074 4016 21014
rect 4160 21004 4212 21010
rect 4160 20946 4212 20952
rect 4172 20369 4200 20946
rect 4158 20360 4214 20369
rect 4158 20295 4214 20304
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 4158 20224 4214 20233
rect 4080 20058 4108 20198
rect 4158 20159 4214 20168
rect 4068 20052 4120 20058
rect 4068 19994 4120 20000
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 4080 18601 4108 19858
rect 4066 18592 4122 18601
rect 4066 18527 4122 18536
rect 4066 18456 4122 18465
rect 4172 18442 4200 20159
rect 4252 19780 4304 19786
rect 4252 19722 4304 19728
rect 4264 18737 4292 19722
rect 4250 18728 4306 18737
rect 4250 18663 4306 18672
rect 4172 18414 4292 18442
rect 4066 18391 4122 18400
rect 4080 16454 4108 18391
rect 4160 18284 4212 18290
rect 4160 18226 4212 18232
rect 4172 17134 4200 18226
rect 4264 18193 4292 18414
rect 4250 18184 4306 18193
rect 4250 18119 4306 18128
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4172 15706 4200 17070
rect 4264 16590 4292 18022
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4356 15552 4384 22442
rect 4448 19990 4476 22646
rect 4540 22506 4568 24278
rect 4712 24268 4764 24274
rect 4712 24210 4764 24216
rect 4620 24132 4672 24138
rect 4620 24074 4672 24080
rect 4528 22500 4580 22506
rect 4528 22442 4580 22448
rect 4526 22400 4582 22409
rect 4526 22335 4582 22344
rect 4540 21672 4568 22335
rect 4632 22030 4660 24074
rect 4620 22024 4672 22030
rect 4620 21966 4672 21972
rect 4540 21644 4660 21672
rect 4528 21548 4580 21554
rect 4528 21490 4580 21496
rect 4540 20330 4568 21490
rect 4528 20324 4580 20330
rect 4528 20266 4580 20272
rect 4632 20210 4660 21644
rect 4724 21026 4752 24210
rect 4908 22545 4936 24754
rect 5000 23746 5028 27474
rect 5172 27396 5224 27402
rect 5172 27338 5224 27344
rect 5080 26784 5132 26790
rect 5080 26726 5132 26732
rect 5092 25888 5120 26726
rect 5184 26518 5212 27338
rect 5276 27130 5304 28018
rect 5816 27872 5868 27878
rect 5816 27814 5868 27820
rect 5442 27772 5750 27792
rect 5442 27770 5448 27772
rect 5504 27770 5528 27772
rect 5584 27770 5608 27772
rect 5664 27770 5688 27772
rect 5744 27770 5750 27772
rect 5504 27718 5506 27770
rect 5686 27718 5688 27770
rect 5442 27716 5448 27718
rect 5504 27716 5528 27718
rect 5584 27716 5608 27718
rect 5664 27716 5688 27718
rect 5744 27716 5750 27718
rect 5442 27696 5750 27716
rect 5828 27606 5856 27814
rect 5448 27600 5500 27606
rect 5448 27542 5500 27548
rect 5540 27600 5592 27606
rect 5540 27542 5592 27548
rect 5816 27600 5868 27606
rect 5816 27542 5868 27548
rect 5264 27124 5316 27130
rect 5264 27066 5316 27072
rect 5460 26897 5488 27542
rect 5552 26994 5580 27542
rect 5816 27124 5868 27130
rect 5816 27066 5868 27072
rect 5540 26988 5592 26994
rect 5540 26930 5592 26936
rect 5446 26888 5502 26897
rect 5446 26823 5502 26832
rect 5356 26784 5408 26790
rect 5356 26726 5408 26732
rect 5172 26512 5224 26518
rect 5172 26454 5224 26460
rect 5184 25956 5212 26454
rect 5368 26450 5396 26726
rect 5442 26684 5750 26704
rect 5442 26682 5448 26684
rect 5504 26682 5528 26684
rect 5584 26682 5608 26684
rect 5664 26682 5688 26684
rect 5744 26682 5750 26684
rect 5504 26630 5506 26682
rect 5686 26630 5688 26682
rect 5442 26628 5448 26630
rect 5504 26628 5528 26630
rect 5584 26628 5608 26630
rect 5664 26628 5688 26630
rect 5744 26628 5750 26630
rect 5442 26608 5750 26628
rect 5828 26586 5856 27066
rect 5816 26580 5868 26586
rect 5816 26522 5868 26528
rect 5356 26444 5408 26450
rect 5356 26386 5408 26392
rect 5448 26444 5500 26450
rect 5448 26386 5500 26392
rect 5264 26376 5316 26382
rect 5264 26318 5316 26324
rect 5276 26081 5304 26318
rect 5262 26072 5318 26081
rect 5262 26007 5318 26016
rect 5264 25968 5316 25974
rect 5184 25928 5264 25956
rect 5264 25910 5316 25916
rect 5092 25860 5212 25888
rect 5078 25528 5134 25537
rect 5184 25498 5212 25860
rect 5078 25463 5134 25472
rect 5172 25492 5224 25498
rect 5092 25294 5120 25463
rect 5172 25434 5224 25440
rect 5080 25288 5132 25294
rect 5080 25230 5132 25236
rect 5092 24138 5120 25230
rect 5080 24132 5132 24138
rect 5080 24074 5132 24080
rect 5184 23905 5212 25434
rect 5276 24410 5304 25910
rect 5460 25906 5488 26386
rect 5632 26376 5684 26382
rect 5920 26330 5948 28154
rect 6552 28008 6604 28014
rect 6552 27950 6604 27956
rect 6182 27568 6238 27577
rect 6182 27503 6238 27512
rect 6000 27464 6052 27470
rect 6000 27406 6052 27412
rect 5632 26318 5684 26324
rect 5644 25945 5672 26318
rect 5828 26302 5948 26330
rect 5630 25936 5686 25945
rect 5448 25900 5500 25906
rect 5368 25860 5448 25888
rect 5368 25158 5396 25860
rect 5630 25871 5686 25880
rect 5448 25842 5500 25848
rect 5442 25596 5750 25616
rect 5442 25594 5448 25596
rect 5504 25594 5528 25596
rect 5584 25594 5608 25596
rect 5664 25594 5688 25596
rect 5744 25594 5750 25596
rect 5504 25542 5506 25594
rect 5686 25542 5688 25594
rect 5442 25540 5448 25542
rect 5504 25540 5528 25542
rect 5584 25540 5608 25542
rect 5664 25540 5688 25542
rect 5744 25540 5750 25542
rect 5442 25520 5750 25540
rect 5724 25288 5776 25294
rect 5724 25230 5776 25236
rect 5356 25152 5408 25158
rect 5356 25094 5408 25100
rect 5736 24818 5764 25230
rect 5828 24954 5856 26302
rect 5908 26240 5960 26246
rect 5908 26182 5960 26188
rect 5920 25537 5948 26182
rect 5906 25528 5962 25537
rect 5906 25463 5962 25472
rect 5908 25356 5960 25362
rect 5908 25298 5960 25304
rect 5816 24948 5868 24954
rect 5816 24890 5868 24896
rect 5920 24818 5948 25298
rect 5540 24812 5592 24818
rect 5540 24754 5592 24760
rect 5724 24812 5776 24818
rect 5724 24754 5776 24760
rect 5908 24812 5960 24818
rect 5908 24754 5960 24760
rect 5552 24721 5580 24754
rect 5632 24744 5684 24750
rect 5538 24712 5594 24721
rect 5684 24692 5856 24698
rect 5632 24686 5856 24692
rect 5644 24670 5856 24686
rect 5538 24647 5594 24656
rect 5442 24508 5750 24528
rect 5442 24506 5448 24508
rect 5504 24506 5528 24508
rect 5584 24506 5608 24508
rect 5664 24506 5688 24508
rect 5744 24506 5750 24508
rect 5504 24454 5506 24506
rect 5686 24454 5688 24506
rect 5442 24452 5448 24454
rect 5504 24452 5528 24454
rect 5584 24452 5608 24454
rect 5664 24452 5688 24454
rect 5744 24452 5750 24454
rect 5442 24432 5750 24452
rect 5264 24404 5316 24410
rect 5264 24346 5316 24352
rect 5828 24342 5856 24670
rect 5920 24410 5948 24754
rect 5908 24404 5960 24410
rect 5908 24346 5960 24352
rect 5816 24336 5868 24342
rect 5816 24278 5868 24284
rect 5356 24268 5408 24274
rect 5356 24210 5408 24216
rect 5170 23896 5226 23905
rect 5368 23866 5396 24210
rect 5908 24064 5960 24070
rect 5908 24006 5960 24012
rect 5170 23831 5226 23840
rect 5356 23860 5408 23866
rect 5356 23802 5408 23808
rect 5000 23718 5212 23746
rect 5080 23112 5132 23118
rect 5080 23054 5132 23060
rect 4988 23044 5040 23050
rect 4988 22986 5040 22992
rect 4894 22536 4950 22545
rect 4894 22471 4950 22480
rect 4804 22432 4856 22438
rect 4804 22374 4856 22380
rect 4896 22432 4948 22438
rect 4896 22374 4948 22380
rect 4816 21554 4844 22374
rect 4908 21690 4936 22374
rect 5000 22234 5028 22986
rect 4988 22228 5040 22234
rect 4988 22170 5040 22176
rect 4988 21956 5040 21962
rect 4988 21898 5040 21904
rect 4896 21684 4948 21690
rect 4896 21626 4948 21632
rect 5000 21622 5028 21898
rect 5092 21894 5120 23054
rect 5080 21888 5132 21894
rect 5080 21830 5132 21836
rect 4988 21616 5040 21622
rect 4988 21558 5040 21564
rect 5092 21554 5120 21830
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 5080 21548 5132 21554
rect 5080 21490 5132 21496
rect 5078 21448 5134 21457
rect 5078 21383 5134 21392
rect 4896 21344 4948 21350
rect 4894 21312 4896 21321
rect 4988 21344 5040 21350
rect 4948 21312 4950 21321
rect 4988 21286 5040 21292
rect 4894 21247 4950 21256
rect 5000 21146 5028 21286
rect 4988 21140 5040 21146
rect 4988 21082 5040 21088
rect 4724 20998 5028 21026
rect 4804 20936 4856 20942
rect 4804 20878 4856 20884
rect 4712 20868 4764 20874
rect 4712 20810 4764 20816
rect 4540 20182 4660 20210
rect 4436 19984 4488 19990
rect 4436 19926 4488 19932
rect 4448 19514 4476 19926
rect 4436 19508 4488 19514
rect 4436 19450 4488 19456
rect 4434 19272 4490 19281
rect 4434 19207 4490 19216
rect 4448 18630 4476 19207
rect 4436 18624 4488 18630
rect 4436 18566 4488 18572
rect 4540 16998 4568 20182
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4632 18601 4660 19110
rect 4618 18592 4674 18601
rect 4618 18527 4674 18536
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 4632 17066 4660 18226
rect 4724 17649 4752 20810
rect 4710 17640 4766 17649
rect 4710 17575 4766 17584
rect 4620 17060 4672 17066
rect 4620 17002 4672 17008
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4356 15524 4568 15552
rect 4436 15428 4488 15434
rect 4436 15370 4488 15376
rect 4448 15094 4476 15370
rect 4436 15088 4488 15094
rect 4436 15030 4488 15036
rect 4160 14884 4212 14890
rect 4160 14826 4212 14832
rect 4172 14414 4200 14826
rect 4344 14816 4396 14822
rect 4344 14758 4396 14764
rect 4356 14482 4384 14758
rect 4344 14476 4396 14482
rect 4344 14418 4396 14424
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4252 14408 4304 14414
rect 4252 14350 4304 14356
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 3896 13926 4016 13954
rect 3882 13832 3938 13841
rect 3882 13767 3938 13776
rect 3896 13462 3924 13767
rect 3884 13456 3936 13462
rect 3884 13398 3936 13404
rect 3896 11694 3924 13398
rect 3988 12442 4016 13926
rect 4160 13728 4212 13734
rect 4160 13670 4212 13676
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 4080 12238 4108 13126
rect 4172 12646 4200 13670
rect 4264 12986 4292 14350
rect 4356 14006 4384 14418
rect 4344 14000 4396 14006
rect 4344 13942 4396 13948
rect 4356 13870 4384 13942
rect 4344 13864 4396 13870
rect 4344 13806 4396 13812
rect 4356 13394 4384 13806
rect 4344 13388 4396 13394
rect 4344 13330 4396 13336
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4356 12918 4384 13330
rect 4344 12912 4396 12918
rect 4264 12860 4344 12866
rect 4264 12854 4396 12860
rect 4264 12838 4384 12854
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4158 12472 4214 12481
rect 4158 12407 4214 12416
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 4066 12064 4122 12073
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 3988 11626 4016 12038
rect 4066 11999 4122 12008
rect 3976 11620 4028 11626
rect 3976 11562 4028 11568
rect 3884 11280 3936 11286
rect 3884 11222 3936 11228
rect 3896 10810 3924 11222
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3988 10470 4016 11562
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3804 9574 3924 9602
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3804 7886 3832 9454
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 3620 6956 3740 6984
rect 3606 6896 3662 6905
rect 3606 6831 3608 6840
rect 3660 6831 3662 6840
rect 3608 6802 3660 6808
rect 3608 6724 3660 6730
rect 3608 6666 3660 6672
rect 3620 5234 3648 6666
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3606 5128 3662 5137
rect 3606 5063 3662 5072
rect 3620 3210 3648 5063
rect 3712 4706 3740 6956
rect 3804 5273 3832 7482
rect 3896 5370 3924 9574
rect 3988 9110 4016 10406
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 3974 8528 4030 8537
rect 3974 8463 3976 8472
rect 4028 8463 4030 8472
rect 3976 8434 4028 8440
rect 4080 8294 4108 11999
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3790 5264 3846 5273
rect 3790 5199 3846 5208
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3804 4826 3832 5102
rect 3988 4842 4016 8026
rect 4080 7274 4108 8026
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 4066 7168 4122 7177
rect 4066 7103 4122 7112
rect 4080 5846 4108 7103
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3896 4814 4016 4842
rect 3712 4678 3832 4706
rect 3698 3768 3754 3777
rect 3698 3703 3754 3712
rect 3712 3466 3740 3703
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 3620 3182 3740 3210
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3620 2650 3648 2994
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 3516 2576 3568 2582
rect 3516 2518 3568 2524
rect 3712 2514 3740 3182
rect 3700 2508 3752 2514
rect 3700 2450 3752 2456
rect 3804 1970 3832 4678
rect 3792 1964 3844 1970
rect 3792 1906 3844 1912
rect 3436 1414 3648 1442
rect 3620 800 3648 1414
rect 3896 800 3924 4814
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3988 3398 4016 4082
rect 4080 3942 4108 5170
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 4172 800 4200 12407
rect 4264 11082 4292 12838
rect 4344 12640 4396 12646
rect 4396 12600 4476 12628
rect 4344 12582 4396 12588
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4356 11762 4384 12378
rect 4448 11830 4476 12600
rect 4540 12442 4568 15524
rect 4620 13252 4672 13258
rect 4620 13194 4672 13200
rect 4632 12986 4660 13194
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4526 12336 4582 12345
rect 4526 12271 4582 12280
rect 4436 11824 4488 11830
rect 4436 11766 4488 11772
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 4436 11688 4488 11694
rect 4436 11630 4488 11636
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4344 11008 4396 11014
rect 4344 10950 4396 10956
rect 4356 10198 4384 10950
rect 4344 10192 4396 10198
rect 4344 10134 4396 10140
rect 4252 9988 4304 9994
rect 4252 9930 4304 9936
rect 4264 9382 4292 9930
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4356 9654 4384 9862
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4356 9058 4384 9590
rect 4264 9030 4384 9058
rect 4264 8401 4292 9030
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4250 8392 4306 8401
rect 4250 8327 4306 8336
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4264 7478 4292 8230
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 4356 7410 4384 8910
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4264 5914 4292 7142
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4264 5794 4292 5850
rect 4264 5766 4384 5794
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4264 5302 4292 5646
rect 4252 5296 4304 5302
rect 4252 5238 4304 5244
rect 4264 4826 4292 5238
rect 4356 5098 4384 5766
rect 4344 5092 4396 5098
rect 4344 5034 4396 5040
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 4356 4758 4384 5034
rect 4344 4752 4396 4758
rect 4344 4694 4396 4700
rect 4448 4570 4476 11630
rect 4252 4548 4304 4554
rect 4252 4490 4304 4496
rect 4356 4542 4476 4570
rect 4264 4214 4292 4490
rect 4356 4282 4384 4542
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4436 4072 4488 4078
rect 4436 4014 4488 4020
rect 4252 4004 4304 4010
rect 4252 3946 4304 3952
rect 4264 3534 4292 3946
rect 4448 3738 4476 4014
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4356 800 4384 3674
rect 4540 2774 4568 12271
rect 4632 8566 4660 12922
rect 4724 12918 4752 16934
rect 4712 12912 4764 12918
rect 4712 12854 4764 12860
rect 4710 12472 4766 12481
rect 4710 12407 4766 12416
rect 4724 12238 4752 12407
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4710 12064 4766 12073
rect 4710 11999 4766 12008
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4632 7886 4660 8230
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4724 4622 4752 11999
rect 4816 11694 4844 20878
rect 4896 20460 4948 20466
rect 4896 20402 4948 20408
rect 4908 19786 4936 20402
rect 4896 19780 4948 19786
rect 4896 19722 4948 19728
rect 4896 19508 4948 19514
rect 4896 19450 4948 19456
rect 4908 18766 4936 19450
rect 4896 18760 4948 18766
rect 4896 18702 4948 18708
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 4908 17746 4936 18158
rect 4896 17740 4948 17746
rect 4896 17682 4948 17688
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 4908 17270 4936 17478
rect 4896 17264 4948 17270
rect 4896 17206 4948 17212
rect 5000 17082 5028 20998
rect 4908 17054 5028 17082
rect 4908 13297 4936 17054
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 5000 16590 5028 16934
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 5000 15706 5028 16186
rect 4988 15700 5040 15706
rect 4988 15642 5040 15648
rect 5092 15450 5120 21383
rect 5184 17218 5212 23718
rect 5264 23724 5316 23730
rect 5264 23666 5316 23672
rect 5276 22545 5304 23666
rect 5356 23656 5408 23662
rect 5356 23598 5408 23604
rect 5368 23254 5396 23598
rect 5442 23420 5750 23440
rect 5442 23418 5448 23420
rect 5504 23418 5528 23420
rect 5584 23418 5608 23420
rect 5664 23418 5688 23420
rect 5744 23418 5750 23420
rect 5504 23366 5506 23418
rect 5686 23366 5688 23418
rect 5442 23364 5448 23366
rect 5504 23364 5528 23366
rect 5584 23364 5608 23366
rect 5664 23364 5688 23366
rect 5744 23364 5750 23366
rect 5442 23344 5750 23364
rect 5920 23322 5948 24006
rect 5908 23316 5960 23322
rect 5908 23258 5960 23264
rect 5356 23248 5408 23254
rect 5356 23190 5408 23196
rect 5814 23080 5870 23089
rect 5356 23044 5408 23050
rect 5814 23015 5870 23024
rect 5356 22986 5408 22992
rect 5368 22778 5396 22986
rect 5446 22808 5502 22817
rect 5356 22772 5408 22778
rect 5446 22743 5502 22752
rect 5356 22714 5408 22720
rect 5460 22642 5488 22743
rect 5448 22636 5500 22642
rect 5448 22578 5500 22584
rect 5262 22536 5318 22545
rect 5262 22471 5318 22480
rect 5368 22506 5488 22522
rect 5368 22500 5500 22506
rect 5368 22494 5448 22500
rect 5264 22432 5316 22438
rect 5264 22374 5316 22380
rect 5276 20058 5304 22374
rect 5368 22094 5396 22494
rect 5448 22442 5500 22448
rect 5442 22332 5750 22352
rect 5442 22330 5448 22332
rect 5504 22330 5528 22332
rect 5584 22330 5608 22332
rect 5664 22330 5688 22332
rect 5744 22330 5750 22332
rect 5504 22278 5506 22330
rect 5686 22278 5688 22330
rect 5442 22276 5448 22278
rect 5504 22276 5528 22278
rect 5584 22276 5608 22278
rect 5664 22276 5688 22278
rect 5744 22276 5750 22278
rect 5442 22256 5750 22276
rect 5540 22160 5592 22166
rect 5540 22102 5592 22108
rect 5368 22066 5488 22094
rect 5368 22030 5396 22066
rect 5356 22024 5408 22030
rect 5356 21966 5408 21972
rect 5460 21842 5488 22066
rect 5552 22030 5580 22102
rect 5540 22024 5592 22030
rect 5540 21966 5592 21972
rect 5368 21814 5488 21842
rect 5368 20806 5396 21814
rect 5552 21554 5580 21966
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5442 21244 5750 21264
rect 5442 21242 5448 21244
rect 5504 21242 5528 21244
rect 5584 21242 5608 21244
rect 5664 21242 5688 21244
rect 5744 21242 5750 21244
rect 5504 21190 5506 21242
rect 5686 21190 5688 21242
rect 5442 21188 5448 21190
rect 5504 21188 5528 21190
rect 5584 21188 5608 21190
rect 5664 21188 5688 21190
rect 5744 21188 5750 21190
rect 5442 21168 5750 21188
rect 5356 20800 5408 20806
rect 5356 20742 5408 20748
rect 5448 20800 5500 20806
rect 5448 20742 5500 20748
rect 5354 20632 5410 20641
rect 5354 20567 5410 20576
rect 5264 20052 5316 20058
rect 5264 19994 5316 20000
rect 5264 19848 5316 19854
rect 5264 19790 5316 19796
rect 5276 19242 5304 19790
rect 5264 19236 5316 19242
rect 5264 19178 5316 19184
rect 5262 19136 5318 19145
rect 5262 19071 5318 19080
rect 5276 17377 5304 19071
rect 5368 18850 5396 20567
rect 5460 20534 5488 20742
rect 5448 20528 5500 20534
rect 5448 20470 5500 20476
rect 5442 20156 5750 20176
rect 5442 20154 5448 20156
rect 5504 20154 5528 20156
rect 5584 20154 5608 20156
rect 5664 20154 5688 20156
rect 5744 20154 5750 20156
rect 5504 20102 5506 20154
rect 5686 20102 5688 20154
rect 5442 20100 5448 20102
rect 5504 20100 5528 20102
rect 5584 20100 5608 20102
rect 5664 20100 5688 20102
rect 5744 20100 5750 20102
rect 5442 20080 5750 20100
rect 5442 19068 5750 19088
rect 5442 19066 5448 19068
rect 5504 19066 5528 19068
rect 5584 19066 5608 19068
rect 5664 19066 5688 19068
rect 5744 19066 5750 19068
rect 5504 19014 5506 19066
rect 5686 19014 5688 19066
rect 5442 19012 5448 19014
rect 5504 19012 5528 19014
rect 5584 19012 5608 19014
rect 5664 19012 5688 19014
rect 5744 19012 5750 19014
rect 5442 18992 5750 19012
rect 5368 18822 5488 18850
rect 5356 18760 5408 18766
rect 5356 18702 5408 18708
rect 5368 18426 5396 18702
rect 5356 18420 5408 18426
rect 5356 18362 5408 18368
rect 5356 18284 5408 18290
rect 5356 18226 5408 18232
rect 5368 17610 5396 18226
rect 5460 18193 5488 18822
rect 5540 18692 5592 18698
rect 5592 18652 5764 18680
rect 5540 18634 5592 18640
rect 5540 18352 5592 18358
rect 5538 18320 5540 18329
rect 5592 18320 5594 18329
rect 5736 18290 5764 18652
rect 5538 18255 5594 18264
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5446 18184 5502 18193
rect 5446 18119 5502 18128
rect 5442 17980 5750 18000
rect 5442 17978 5448 17980
rect 5504 17978 5528 17980
rect 5584 17978 5608 17980
rect 5664 17978 5688 17980
rect 5744 17978 5750 17980
rect 5504 17926 5506 17978
rect 5686 17926 5688 17978
rect 5442 17924 5448 17926
rect 5504 17924 5528 17926
rect 5584 17924 5608 17926
rect 5664 17924 5688 17926
rect 5744 17924 5750 17926
rect 5442 17904 5750 17924
rect 5632 17740 5684 17746
rect 5632 17682 5684 17688
rect 5356 17604 5408 17610
rect 5356 17546 5408 17552
rect 5262 17368 5318 17377
rect 5262 17303 5318 17312
rect 5184 17190 5304 17218
rect 5368 17202 5396 17546
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5552 17270 5580 17478
rect 5540 17264 5592 17270
rect 5540 17206 5592 17212
rect 5644 17202 5672 17682
rect 5724 17536 5776 17542
rect 5724 17478 5776 17484
rect 5736 17338 5764 17478
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5828 17218 5856 23015
rect 5908 22976 5960 22982
rect 5908 22918 5960 22924
rect 5920 21962 5948 22918
rect 5908 21956 5960 21962
rect 5908 21898 5960 21904
rect 5906 20360 5962 20369
rect 5906 20295 5962 20304
rect 5920 18358 5948 20295
rect 5908 18352 5960 18358
rect 5908 18294 5960 18300
rect 5908 18148 5960 18154
rect 5908 18090 5960 18096
rect 5920 17678 5948 18090
rect 5908 17672 5960 17678
rect 5908 17614 5960 17620
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 5184 15706 5212 16526
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5000 15422 5120 15450
rect 4894 13288 4950 13297
rect 4894 13223 4950 13232
rect 4896 12912 4948 12918
rect 4896 12854 4948 12860
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4816 10062 4844 10406
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4802 9888 4858 9897
rect 4802 9823 4858 9832
rect 4816 5658 4844 9823
rect 4908 5778 4936 12854
rect 5000 12306 5028 15422
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 5184 15162 5212 15302
rect 5172 15156 5224 15162
rect 5172 15098 5224 15104
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 5092 12850 5120 14214
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5184 13394 5212 13670
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5170 13288 5226 13297
rect 5170 13223 5226 13232
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 5080 12708 5132 12714
rect 5080 12650 5132 12656
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 5092 11762 5120 12650
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 5078 11656 5134 11665
rect 5078 11591 5134 11600
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 5000 10742 5028 10950
rect 4988 10736 5040 10742
rect 4988 10678 5040 10684
rect 4988 10532 5040 10538
rect 4988 10474 5040 10480
rect 5000 9994 5028 10474
rect 4988 9988 5040 9994
rect 4988 9930 5040 9936
rect 5092 9874 5120 11591
rect 5000 9846 5120 9874
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4816 5630 4936 5658
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4620 4072 4672 4078
rect 4620 4014 4672 4020
rect 4632 3058 4660 4014
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4724 2854 4752 4082
rect 4816 4010 4844 5510
rect 4908 5098 4936 5630
rect 4896 5092 4948 5098
rect 4896 5034 4948 5040
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4908 4282 4936 4762
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 5000 4146 5028 9846
rect 5078 9752 5134 9761
rect 5078 9687 5134 9696
rect 5092 6905 5120 9687
rect 5078 6896 5134 6905
rect 5078 6831 5134 6840
rect 5080 6724 5132 6730
rect 5080 6666 5132 6672
rect 5092 5914 5120 6666
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4804 4004 4856 4010
rect 4804 3946 4856 3952
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 4816 3194 4844 3538
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4908 2922 4936 3470
rect 5092 3126 5120 4558
rect 5080 3120 5132 3126
rect 5080 3062 5132 3068
rect 5092 2990 5120 3062
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4540 2746 4660 2774
rect 4632 800 4660 2746
rect 4724 2446 4752 2790
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 4908 800 4936 2518
rect 5184 800 5212 13223
rect 5276 12617 5304 17190
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 5632 17196 5684 17202
rect 5828 17190 5948 17218
rect 5632 17138 5684 17144
rect 5816 17128 5868 17134
rect 5816 17070 5868 17076
rect 5442 16892 5750 16912
rect 5442 16890 5448 16892
rect 5504 16890 5528 16892
rect 5584 16890 5608 16892
rect 5664 16890 5688 16892
rect 5744 16890 5750 16892
rect 5504 16838 5506 16890
rect 5686 16838 5688 16890
rect 5442 16836 5448 16838
rect 5504 16836 5528 16838
rect 5584 16836 5608 16838
rect 5664 16836 5688 16838
rect 5744 16836 5750 16838
rect 5442 16816 5750 16836
rect 5828 16658 5856 17070
rect 5816 16652 5868 16658
rect 5816 16594 5868 16600
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5460 16114 5488 16390
rect 5828 16182 5856 16594
rect 5816 16176 5868 16182
rect 5816 16118 5868 16124
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5442 15804 5750 15824
rect 5442 15802 5448 15804
rect 5504 15802 5528 15804
rect 5584 15802 5608 15804
rect 5664 15802 5688 15804
rect 5744 15802 5750 15804
rect 5504 15750 5506 15802
rect 5686 15750 5688 15802
rect 5442 15748 5448 15750
rect 5504 15748 5528 15750
rect 5584 15748 5608 15750
rect 5664 15748 5688 15750
rect 5744 15748 5750 15750
rect 5442 15728 5750 15748
rect 5828 15706 5856 16118
rect 5816 15700 5868 15706
rect 5816 15642 5868 15648
rect 5442 14716 5750 14736
rect 5442 14714 5448 14716
rect 5504 14714 5528 14716
rect 5584 14714 5608 14716
rect 5664 14714 5688 14716
rect 5744 14714 5750 14716
rect 5504 14662 5506 14714
rect 5686 14662 5688 14714
rect 5442 14660 5448 14662
rect 5504 14660 5528 14662
rect 5584 14660 5608 14662
rect 5664 14660 5688 14662
rect 5744 14660 5750 14662
rect 5442 14640 5750 14660
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5828 14006 5856 14214
rect 5816 14000 5868 14006
rect 5816 13942 5868 13948
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 5368 13530 5396 13670
rect 5442 13628 5750 13648
rect 5442 13626 5448 13628
rect 5504 13626 5528 13628
rect 5584 13626 5608 13628
rect 5664 13626 5688 13628
rect 5744 13626 5750 13628
rect 5504 13574 5506 13626
rect 5686 13574 5688 13626
rect 5442 13572 5448 13574
rect 5504 13572 5528 13574
rect 5584 13572 5608 13574
rect 5664 13572 5688 13574
rect 5744 13572 5750 13574
rect 5442 13552 5750 13572
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5262 12608 5318 12617
rect 5262 12543 5318 12552
rect 5262 12472 5318 12481
rect 5262 12407 5318 12416
rect 5276 11898 5304 12407
rect 5368 12238 5396 13466
rect 5448 13252 5500 13258
rect 5448 13194 5500 13200
rect 5460 12714 5488 13194
rect 5540 12912 5592 12918
rect 5538 12880 5540 12889
rect 5592 12880 5594 12889
rect 5538 12815 5594 12824
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5442 12540 5750 12560
rect 5442 12538 5448 12540
rect 5504 12538 5528 12540
rect 5584 12538 5608 12540
rect 5664 12538 5688 12540
rect 5744 12538 5750 12540
rect 5504 12486 5506 12538
rect 5686 12486 5688 12538
rect 5442 12484 5448 12486
rect 5504 12484 5528 12486
rect 5584 12484 5608 12486
rect 5664 12484 5688 12486
rect 5744 12484 5750 12486
rect 5442 12464 5750 12484
rect 5920 12458 5948 17190
rect 5828 12406 5948 12458
rect 5724 12368 5776 12374
rect 5724 12310 5776 12316
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5356 11688 5408 11694
rect 5552 11676 5580 12106
rect 5408 11648 5580 11676
rect 5356 11630 5408 11636
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 5276 10674 5304 10950
rect 5368 10674 5396 11630
rect 5736 11626 5764 12310
rect 5920 12220 5948 12406
rect 6012 12374 6040 27406
rect 6090 27024 6146 27033
rect 6090 26959 6092 26968
rect 6144 26959 6146 26968
rect 6092 26930 6144 26936
rect 6196 26926 6224 27503
rect 6460 27464 6512 27470
rect 6564 27452 6592 27950
rect 6828 27940 6880 27946
rect 6828 27882 6880 27888
rect 6644 27668 6696 27674
rect 6644 27610 6696 27616
rect 6512 27424 6592 27452
rect 6460 27406 6512 27412
rect 6368 27396 6420 27402
rect 6368 27338 6420 27344
rect 6380 27130 6408 27338
rect 6368 27124 6420 27130
rect 6368 27066 6420 27072
rect 6184 26920 6236 26926
rect 6184 26862 6236 26868
rect 6092 26376 6144 26382
rect 6092 26318 6144 26324
rect 6184 26376 6236 26382
rect 6184 26318 6236 26324
rect 6104 25294 6132 26318
rect 6092 25288 6144 25294
rect 6092 25230 6144 25236
rect 6104 24682 6132 25230
rect 6196 24750 6224 26318
rect 6460 26240 6512 26246
rect 6460 26182 6512 26188
rect 6366 26072 6422 26081
rect 6366 26007 6422 26016
rect 6276 25696 6328 25702
rect 6276 25638 6328 25644
rect 6184 24744 6236 24750
rect 6184 24686 6236 24692
rect 6092 24676 6144 24682
rect 6092 24618 6144 24624
rect 6104 23866 6132 24618
rect 6184 24608 6236 24614
rect 6182 24576 6184 24585
rect 6236 24576 6238 24585
rect 6182 24511 6238 24520
rect 6184 24336 6236 24342
rect 6184 24278 6236 24284
rect 6092 23860 6144 23866
rect 6092 23802 6144 23808
rect 6196 22930 6224 24278
rect 6288 23066 6316 25638
rect 6380 25226 6408 26007
rect 6472 25702 6500 26182
rect 6460 25696 6512 25702
rect 6460 25638 6512 25644
rect 6458 25528 6514 25537
rect 6458 25463 6514 25472
rect 6368 25220 6420 25226
rect 6368 25162 6420 25168
rect 6472 24954 6500 25463
rect 6460 24948 6512 24954
rect 6380 24908 6460 24936
rect 6380 24206 6408 24908
rect 6460 24890 6512 24896
rect 6460 24744 6512 24750
rect 6460 24686 6512 24692
rect 6368 24200 6420 24206
rect 6368 24142 6420 24148
rect 6368 24064 6420 24070
rect 6368 24006 6420 24012
rect 6380 23322 6408 24006
rect 6368 23316 6420 23322
rect 6368 23258 6420 23264
rect 6472 23254 6500 24686
rect 6460 23248 6512 23254
rect 6460 23190 6512 23196
rect 6288 23038 6500 23066
rect 6196 22902 6408 22930
rect 6276 22772 6328 22778
rect 6276 22714 6328 22720
rect 6092 22568 6144 22574
rect 6092 22510 6144 22516
rect 6104 22098 6132 22510
rect 6092 22092 6144 22098
rect 6092 22034 6144 22040
rect 6184 21004 6236 21010
rect 6184 20946 6236 20952
rect 6196 20641 6224 20946
rect 6182 20632 6238 20641
rect 6182 20567 6238 20576
rect 6092 20460 6144 20466
rect 6092 20402 6144 20408
rect 6104 19854 6132 20402
rect 6184 20392 6236 20398
rect 6184 20334 6236 20340
rect 6196 19922 6224 20334
rect 6184 19916 6236 19922
rect 6184 19858 6236 19864
rect 6092 19848 6144 19854
rect 6092 19790 6144 19796
rect 6104 19514 6132 19790
rect 6092 19508 6144 19514
rect 6092 19450 6144 19456
rect 6104 19378 6132 19450
rect 6092 19372 6144 19378
rect 6288 19334 6316 22714
rect 6092 19314 6144 19320
rect 6196 19306 6316 19334
rect 6092 18624 6144 18630
rect 6092 18566 6144 18572
rect 6000 12368 6052 12374
rect 6000 12310 6052 12316
rect 5828 12192 5948 12220
rect 6000 12232 6052 12238
rect 5724 11620 5776 11626
rect 5724 11562 5776 11568
rect 5442 11452 5750 11472
rect 5442 11450 5448 11452
rect 5504 11450 5528 11452
rect 5584 11450 5608 11452
rect 5664 11450 5688 11452
rect 5744 11450 5750 11452
rect 5504 11398 5506 11450
rect 5686 11398 5688 11450
rect 5442 11396 5448 11398
rect 5504 11396 5528 11398
rect 5584 11396 5608 11398
rect 5664 11396 5688 11398
rect 5744 11396 5750 11398
rect 5442 11376 5750 11396
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5540 10736 5592 10742
rect 5736 10690 5764 10746
rect 5592 10684 5764 10690
rect 5540 10678 5764 10684
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5356 10668 5408 10674
rect 5552 10662 5764 10678
rect 5356 10610 5408 10616
rect 5276 10062 5304 10610
rect 5368 10248 5396 10610
rect 5442 10364 5750 10384
rect 5442 10362 5448 10364
rect 5504 10362 5528 10364
rect 5584 10362 5608 10364
rect 5664 10362 5688 10364
rect 5744 10362 5750 10364
rect 5504 10310 5506 10362
rect 5686 10310 5688 10362
rect 5442 10308 5448 10310
rect 5504 10308 5528 10310
rect 5584 10308 5608 10310
rect 5664 10308 5688 10310
rect 5744 10308 5750 10310
rect 5442 10288 5750 10308
rect 5368 10220 5764 10248
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5276 8022 5304 8434
rect 5368 8430 5396 9862
rect 5552 9450 5580 9998
rect 5736 9994 5764 10220
rect 5724 9988 5776 9994
rect 5724 9930 5776 9936
rect 5736 9654 5764 9930
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 5828 9602 5856 12192
rect 6000 12174 6052 12180
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 5920 11762 5948 12038
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 6012 11694 6040 12174
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5920 11150 5948 11494
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 6012 10606 6040 11630
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 5828 9574 6040 9602
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5442 9276 5750 9296
rect 5442 9274 5448 9276
rect 5504 9274 5528 9276
rect 5584 9274 5608 9276
rect 5664 9274 5688 9276
rect 5744 9274 5750 9276
rect 5504 9222 5506 9274
rect 5686 9222 5688 9274
rect 5442 9220 5448 9222
rect 5504 9220 5528 9222
rect 5584 9220 5608 9222
rect 5664 9220 5688 9222
rect 5744 9220 5750 9222
rect 5442 9200 5750 9220
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5276 7410 5304 7686
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5368 6458 5396 8230
rect 5442 8188 5750 8208
rect 5442 8186 5448 8188
rect 5504 8186 5528 8188
rect 5584 8186 5608 8188
rect 5664 8186 5688 8188
rect 5744 8186 5750 8188
rect 5504 8134 5506 8186
rect 5686 8134 5688 8186
rect 5442 8132 5448 8134
rect 5504 8132 5528 8134
rect 5584 8132 5608 8134
rect 5664 8132 5688 8134
rect 5744 8132 5750 8134
rect 5442 8112 5750 8132
rect 5828 7954 5856 9318
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 5920 8906 5948 8978
rect 5908 8900 5960 8906
rect 5908 8842 5960 8848
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5442 7100 5750 7120
rect 5442 7098 5448 7100
rect 5504 7098 5528 7100
rect 5584 7098 5608 7100
rect 5664 7098 5688 7100
rect 5744 7098 5750 7100
rect 5504 7046 5506 7098
rect 5686 7046 5688 7098
rect 5442 7044 5448 7046
rect 5504 7044 5528 7046
rect 5584 7044 5608 7046
rect 5664 7044 5688 7046
rect 5744 7044 5750 7046
rect 5442 7024 5750 7044
rect 5920 6769 5948 8842
rect 5906 6760 5962 6769
rect 5906 6695 5962 6704
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5368 5710 5396 6394
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5442 6012 5750 6032
rect 5442 6010 5448 6012
rect 5504 6010 5528 6012
rect 5584 6010 5608 6012
rect 5664 6010 5688 6012
rect 5744 6010 5750 6012
rect 5504 5958 5506 6010
rect 5686 5958 5688 6010
rect 5442 5956 5448 5958
rect 5504 5956 5528 5958
rect 5584 5956 5608 5958
rect 5664 5956 5688 5958
rect 5744 5956 5750 5958
rect 5442 5936 5750 5956
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5276 5234 5304 5646
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5828 5114 5856 6190
rect 5920 5914 5948 6598
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 5264 5092 5316 5098
rect 5828 5086 5948 5114
rect 5264 5034 5316 5040
rect 5276 4010 5304 5034
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5442 4924 5750 4944
rect 5442 4922 5448 4924
rect 5504 4922 5528 4924
rect 5584 4922 5608 4924
rect 5664 4922 5688 4924
rect 5744 4922 5750 4924
rect 5504 4870 5506 4922
rect 5686 4870 5688 4922
rect 5442 4868 5448 4870
rect 5504 4868 5528 4870
rect 5584 4868 5608 4870
rect 5664 4868 5688 4870
rect 5744 4868 5750 4870
rect 5442 4848 5750 4868
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5368 4282 5396 4490
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5828 4146 5856 4966
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 5262 3768 5318 3777
rect 5262 3703 5318 3712
rect 5276 3466 5304 3703
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5262 3224 5318 3233
rect 5262 3159 5318 3168
rect 5276 3126 5304 3159
rect 5264 3120 5316 3126
rect 5264 3062 5316 3068
rect 5276 2378 5304 3062
rect 5264 2372 5316 2378
rect 5264 2314 5316 2320
rect 5368 1442 5396 4082
rect 5920 4078 5948 5086
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 5442 3836 5750 3856
rect 5442 3834 5448 3836
rect 5504 3834 5528 3836
rect 5584 3834 5608 3836
rect 5664 3834 5688 3836
rect 5744 3834 5750 3836
rect 5504 3782 5506 3834
rect 5686 3782 5688 3834
rect 5442 3780 5448 3782
rect 5504 3780 5528 3782
rect 5584 3780 5608 3782
rect 5664 3780 5688 3782
rect 5744 3780 5750 3782
rect 5442 3760 5750 3780
rect 5446 3632 5502 3641
rect 5446 3567 5502 3576
rect 5540 3596 5592 3602
rect 5460 3126 5488 3567
rect 5540 3538 5592 3544
rect 5552 3194 5580 3538
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5442 2748 5750 2768
rect 5442 2746 5448 2748
rect 5504 2746 5528 2748
rect 5584 2746 5608 2748
rect 5664 2746 5688 2748
rect 5744 2746 5750 2748
rect 5504 2694 5506 2746
rect 5686 2694 5688 2746
rect 5442 2692 5448 2694
rect 5504 2692 5528 2694
rect 5584 2692 5608 2694
rect 5664 2692 5688 2694
rect 5744 2692 5750 2694
rect 5442 2672 5750 2692
rect 5828 2650 5856 3470
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 5722 2544 5778 2553
rect 5722 2479 5778 2488
rect 5368 1414 5488 1442
rect 5460 800 5488 1414
rect 5736 800 5764 2479
rect 5920 2310 5948 3334
rect 5908 2304 5960 2310
rect 5908 2246 5960 2252
rect 6012 800 6040 9574
rect 6104 2774 6132 18566
rect 6196 4078 6224 19306
rect 6380 18630 6408 22902
rect 6368 18624 6420 18630
rect 6368 18566 6420 18572
rect 6472 18442 6500 23038
rect 6564 22438 6592 27424
rect 6656 24138 6684 27610
rect 6840 27418 6868 27882
rect 6840 27390 6960 27418
rect 6828 27328 6880 27334
rect 6748 27288 6828 27316
rect 6644 24132 6696 24138
rect 6644 24074 6696 24080
rect 6656 22574 6684 24074
rect 6644 22568 6696 22574
rect 6644 22510 6696 22516
rect 6552 22432 6604 22438
rect 6552 22374 6604 22380
rect 6564 18766 6592 22374
rect 6644 21888 6696 21894
rect 6644 21830 6696 21836
rect 6656 21622 6684 21830
rect 6644 21616 6696 21622
rect 6644 21558 6696 21564
rect 6644 21480 6696 21486
rect 6642 21448 6644 21457
rect 6696 21448 6698 21457
rect 6642 21383 6698 21392
rect 6644 21140 6696 21146
rect 6644 21082 6696 21088
rect 6656 20262 6684 21082
rect 6748 20890 6776 27288
rect 6828 27270 6880 27276
rect 6932 27146 6960 27390
rect 6840 27118 6960 27146
rect 7012 27124 7064 27130
rect 6840 25888 6868 27118
rect 7012 27066 7064 27072
rect 6840 25860 6960 25888
rect 6828 25764 6880 25770
rect 6828 25706 6880 25712
rect 6840 25294 6868 25706
rect 6828 25288 6880 25294
rect 6828 25230 6880 25236
rect 6932 25106 6960 25860
rect 6840 25078 6960 25106
rect 6840 22778 6868 25078
rect 6920 24744 6972 24750
rect 6918 24712 6920 24721
rect 6972 24712 6974 24721
rect 6918 24647 6974 24656
rect 6920 24608 6972 24614
rect 6918 24576 6920 24585
rect 6972 24576 6974 24585
rect 6918 24511 6974 24520
rect 6920 24268 6972 24274
rect 6920 24210 6972 24216
rect 6932 23662 6960 24210
rect 7024 23866 7052 27066
rect 7012 23860 7064 23866
rect 7012 23802 7064 23808
rect 6920 23656 6972 23662
rect 6920 23598 6972 23604
rect 6932 23322 6960 23598
rect 6920 23316 6972 23322
rect 6920 23258 6972 23264
rect 6828 22772 6880 22778
rect 6828 22714 6880 22720
rect 7024 22710 7052 23802
rect 7012 22704 7064 22710
rect 7012 22646 7064 22652
rect 6920 22568 6972 22574
rect 6920 22510 6972 22516
rect 6932 22030 6960 22510
rect 7012 22432 7064 22438
rect 7012 22374 7064 22380
rect 6920 22024 6972 22030
rect 6920 21966 6972 21972
rect 6828 21888 6880 21894
rect 6828 21830 6880 21836
rect 6840 21554 6868 21830
rect 6828 21548 6880 21554
rect 6828 21490 6880 21496
rect 6932 21486 6960 21966
rect 7024 21554 7052 22374
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 6920 21480 6972 21486
rect 6920 21422 6972 21428
rect 6748 20862 6868 20890
rect 6736 20800 6788 20806
rect 6736 20742 6788 20748
rect 6748 20466 6776 20742
rect 6736 20460 6788 20466
rect 6736 20402 6788 20408
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 6656 19854 6684 20198
rect 6840 20074 6868 20862
rect 6932 20602 6960 21422
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 6748 20046 6868 20074
rect 6644 19848 6696 19854
rect 6644 19790 6696 19796
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 6472 18414 6592 18442
rect 6460 18284 6512 18290
rect 6460 18226 6512 18232
rect 6368 18216 6420 18222
rect 6368 18158 6420 18164
rect 6276 17196 6328 17202
rect 6276 17138 6328 17144
rect 6288 16794 6316 17138
rect 6380 17134 6408 18158
rect 6472 17882 6500 18226
rect 6460 17876 6512 17882
rect 6460 17818 6512 17824
rect 6368 17128 6420 17134
rect 6368 17070 6420 17076
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 6276 16448 6328 16454
rect 6276 16390 6328 16396
rect 6288 14498 6316 16390
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6380 15502 6408 15846
rect 6368 15496 6420 15502
rect 6368 15438 6420 15444
rect 6460 15496 6512 15502
rect 6460 15438 6512 15444
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6380 14822 6408 15302
rect 6472 15162 6500 15438
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6288 14470 6408 14498
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 6288 11898 6316 14350
rect 6380 12918 6408 14470
rect 6460 14340 6512 14346
rect 6460 14282 6512 14288
rect 6368 12912 6420 12918
rect 6368 12854 6420 12860
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6380 12238 6408 12718
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6366 11928 6422 11937
rect 6276 11892 6328 11898
rect 6366 11863 6422 11872
rect 6276 11834 6328 11840
rect 6380 11830 6408 11863
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 6276 11552 6328 11558
rect 6328 11512 6408 11540
rect 6276 11494 6328 11500
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 6288 11150 6316 11222
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6274 10024 6330 10033
rect 6274 9959 6330 9968
rect 6288 7546 6316 9959
rect 6380 8537 6408 11512
rect 6472 11354 6500 14282
rect 6564 12617 6592 18414
rect 6644 17672 6696 17678
rect 6644 17614 6696 17620
rect 6656 13954 6684 17614
rect 6748 16454 6776 20046
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6840 18902 6868 19858
rect 6920 19780 6972 19786
rect 6920 19722 6972 19728
rect 6932 19174 6960 19722
rect 7024 19417 7052 20198
rect 7010 19408 7066 19417
rect 7010 19343 7066 19352
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 6828 18896 6880 18902
rect 6920 18896 6972 18902
rect 6828 18838 6880 18844
rect 6918 18864 6920 18873
rect 6972 18864 6974 18873
rect 6918 18799 6974 18808
rect 7024 18766 7052 19110
rect 7012 18760 7064 18766
rect 6918 18728 6974 18737
rect 7012 18702 7064 18708
rect 6918 18663 6920 18672
rect 6972 18663 6974 18672
rect 6920 18634 6972 18640
rect 6828 18352 6880 18358
rect 6828 18294 6880 18300
rect 6736 16448 6788 16454
rect 6736 16390 6788 16396
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 6748 15162 6776 16050
rect 6840 15609 6868 18294
rect 6826 15600 6882 15609
rect 6826 15535 6882 15544
rect 6828 15428 6880 15434
rect 6828 15370 6880 15376
rect 6840 15162 6868 15370
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6736 14340 6788 14346
rect 6736 14282 6788 14288
rect 6748 14074 6776 14282
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6826 13968 6882 13977
rect 6656 13926 6776 13954
rect 6644 12640 6696 12646
rect 6550 12608 6606 12617
rect 6644 12582 6696 12588
rect 6550 12543 6606 12552
rect 6550 12336 6606 12345
rect 6550 12271 6606 12280
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 6472 10062 6500 11018
rect 6564 10810 6592 12271
rect 6656 12238 6684 12582
rect 6748 12345 6776 13926
rect 6826 13903 6882 13912
rect 6840 12646 6868 13903
rect 6932 12918 6960 18634
rect 7010 18456 7066 18465
rect 7010 18391 7066 18400
rect 7024 15570 7052 18391
rect 7012 15564 7064 15570
rect 7012 15506 7064 15512
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 7024 13326 7052 14214
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6828 12368 6880 12374
rect 6734 12336 6790 12345
rect 6828 12310 6880 12316
rect 6734 12271 6790 12280
rect 6644 12232 6696 12238
rect 6840 12220 6868 12310
rect 6644 12174 6696 12180
rect 6748 12192 6868 12220
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6656 11218 6684 11630
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6656 10674 6684 11154
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6552 10532 6604 10538
rect 6552 10474 6604 10480
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6366 8528 6422 8537
rect 6366 8463 6422 8472
rect 6472 7954 6500 9998
rect 6564 9926 6592 10474
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6564 9586 6592 9862
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6656 9042 6684 9590
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6644 8832 6696 8838
rect 6564 8792 6644 8820
rect 6564 8634 6592 8792
rect 6644 8774 6696 8780
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6550 8528 6606 8537
rect 6656 8498 6684 8570
rect 6550 8463 6606 8472
rect 6644 8492 6696 8498
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 6380 7342 6408 7754
rect 6472 7410 6500 7890
rect 6564 7698 6592 8463
rect 6644 8434 6696 8440
rect 6656 7886 6684 8434
rect 6748 8362 6776 12192
rect 6826 12064 6882 12073
rect 6826 11999 6882 12008
rect 6840 11098 6868 11999
rect 6932 11218 6960 12854
rect 7024 12850 7052 13262
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 7010 12472 7066 12481
rect 7010 12407 7066 12416
rect 7024 11898 7052 12407
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 7012 11144 7064 11150
rect 6840 11070 6960 11098
rect 7012 11086 7064 11092
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6840 10674 6868 10950
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6932 10554 6960 11070
rect 7024 10810 7052 11086
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6840 10526 6960 10554
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 6840 8294 6868 10526
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6932 10130 6960 10202
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6918 10024 6974 10033
rect 6918 9959 6974 9968
rect 6932 8537 6960 9959
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 6918 8528 6974 8537
rect 6918 8463 6974 8472
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6748 7886 6776 8026
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6736 7744 6788 7750
rect 6564 7670 6684 7698
rect 6736 7686 6788 7692
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6380 7002 6408 7278
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6288 4758 6316 6258
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 6380 4128 6408 6938
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6472 4146 6500 5238
rect 6564 4622 6592 6666
rect 6656 5930 6684 7670
rect 6748 7460 6776 7686
rect 6828 7472 6880 7478
rect 6748 7432 6828 7460
rect 6828 7414 6880 7420
rect 6656 5902 6776 5930
rect 6644 5636 6696 5642
rect 6644 5578 6696 5584
rect 6656 5370 6684 5578
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6550 4448 6606 4457
rect 6550 4383 6606 4392
rect 6564 4214 6592 4383
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6656 4146 6684 5170
rect 6748 4690 6776 5902
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6748 4146 6776 4422
rect 6288 4100 6408 4128
rect 6460 4140 6512 4146
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6182 3904 6238 3913
rect 6182 3839 6238 3848
rect 6196 3194 6224 3839
rect 6288 3233 6316 4100
rect 6460 4082 6512 4088
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6274 3224 6330 3233
rect 6184 3188 6236 3194
rect 6274 3159 6330 3168
rect 6184 3130 6236 3136
rect 6276 3052 6328 3058
rect 6380 3040 6408 3878
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6472 3058 6500 3334
rect 6328 3012 6408 3040
rect 6276 2994 6328 3000
rect 6104 2746 6316 2774
rect 6288 800 6316 2746
rect 6380 2582 6408 3012
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6368 2576 6420 2582
rect 6368 2518 6420 2524
rect 6564 800 6592 4014
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6656 2774 6684 3946
rect 6748 3466 6776 4082
rect 6840 3942 6868 7414
rect 6932 7342 6960 8366
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6932 6390 6960 7278
rect 7024 6934 7052 9862
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 7010 6760 7066 6769
rect 7010 6695 7012 6704
rect 7064 6695 7066 6704
rect 7012 6666 7064 6672
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 6932 5250 6960 6326
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 7024 5370 7052 6054
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6932 5222 7052 5250
rect 7024 5166 7052 5222
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6932 4078 6960 4966
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6932 3738 6960 3878
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6736 3460 6788 3466
rect 6736 3402 6788 3408
rect 6826 3224 6882 3233
rect 6932 3194 6960 3470
rect 6826 3159 6882 3168
rect 6920 3188 6972 3194
rect 6840 3074 6868 3159
rect 6920 3130 6972 3136
rect 6840 3046 6960 3074
rect 6656 2746 6868 2774
rect 6840 800 6868 2746
rect 6932 2378 6960 3046
rect 7024 2961 7052 4626
rect 7010 2952 7066 2961
rect 7010 2887 7066 2896
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 7024 2514 7052 2790
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 6920 2372 6972 2378
rect 6920 2314 6972 2320
rect 7012 2372 7064 2378
rect 7012 2314 7064 2320
rect 7024 2106 7052 2314
rect 7012 2100 7064 2106
rect 7012 2042 7064 2048
rect 7116 800 7144 28358
rect 7484 27577 7512 28358
rect 7470 27568 7526 27577
rect 7470 27503 7526 27512
rect 7288 27056 7340 27062
rect 7194 27024 7250 27033
rect 7288 26998 7340 27004
rect 7194 26959 7196 26968
rect 7248 26959 7250 26968
rect 7196 26930 7248 26936
rect 7196 26240 7248 26246
rect 7196 26182 7248 26188
rect 7208 26042 7236 26182
rect 7196 26036 7248 26042
rect 7196 25978 7248 25984
rect 7300 25702 7328 26998
rect 7484 26926 7512 27503
rect 8116 27464 8168 27470
rect 8116 27406 8168 27412
rect 7840 27328 7892 27334
rect 7840 27270 7892 27276
rect 8024 27328 8076 27334
rect 8024 27270 8076 27276
rect 7564 27056 7616 27062
rect 7564 26998 7616 27004
rect 7472 26920 7524 26926
rect 7472 26862 7524 26868
rect 7576 26858 7604 26998
rect 7852 26926 7880 27270
rect 7840 26920 7892 26926
rect 7840 26862 7892 26868
rect 7564 26852 7616 26858
rect 7564 26794 7616 26800
rect 7472 26580 7524 26586
rect 7472 26522 7524 26528
rect 7484 26382 7512 26522
rect 8036 26450 8064 27270
rect 8128 26926 8156 27406
rect 8116 26920 8168 26926
rect 8116 26862 8168 26868
rect 8312 26586 8340 28494
rect 8208 26580 8260 26586
rect 8208 26522 8260 26528
rect 8300 26580 8352 26586
rect 8300 26522 8352 26528
rect 8220 26466 8248 26522
rect 8404 26518 8432 28494
rect 8576 28484 8628 28490
rect 8576 28426 8628 28432
rect 8760 28484 8812 28490
rect 8760 28426 8812 28432
rect 8588 27878 8616 28426
rect 8576 27872 8628 27878
rect 8576 27814 8628 27820
rect 8666 27432 8722 27441
rect 8666 27367 8722 27376
rect 8576 26988 8628 26994
rect 8576 26930 8628 26936
rect 8392 26512 8444 26518
rect 8024 26444 8076 26450
rect 8220 26438 8340 26466
rect 8392 26454 8444 26460
rect 8024 26386 8076 26392
rect 7472 26376 7524 26382
rect 7472 26318 7524 26324
rect 7472 26240 7524 26246
rect 7472 26182 7524 26188
rect 7484 25974 7512 26182
rect 7840 26036 7892 26042
rect 7840 25978 7892 25984
rect 7472 25968 7524 25974
rect 7472 25910 7524 25916
rect 7288 25696 7340 25702
rect 7288 25638 7340 25644
rect 7484 25430 7512 25910
rect 7564 25900 7616 25906
rect 7564 25842 7616 25848
rect 7472 25424 7524 25430
rect 7472 25366 7524 25372
rect 7484 24886 7512 25366
rect 7576 25226 7604 25842
rect 7564 25220 7616 25226
rect 7564 25162 7616 25168
rect 7472 24880 7524 24886
rect 7472 24822 7524 24828
rect 7576 23730 7604 25162
rect 7656 24812 7708 24818
rect 7656 24754 7708 24760
rect 7748 24812 7800 24818
rect 7748 24754 7800 24760
rect 7668 24342 7696 24754
rect 7760 24410 7788 24754
rect 7852 24682 7880 25978
rect 8036 25430 8064 26386
rect 8024 25424 8076 25430
rect 8024 25366 8076 25372
rect 7840 24676 7892 24682
rect 7840 24618 7892 24624
rect 7748 24404 7800 24410
rect 7748 24346 7800 24352
rect 7656 24336 7708 24342
rect 7656 24278 7708 24284
rect 7668 23866 7696 24278
rect 8036 24206 8064 25366
rect 8312 24410 8340 26438
rect 8484 24744 8536 24750
rect 8484 24686 8536 24692
rect 8300 24404 8352 24410
rect 8300 24346 8352 24352
rect 8496 24274 8524 24686
rect 8116 24268 8168 24274
rect 8116 24210 8168 24216
rect 8484 24268 8536 24274
rect 8484 24210 8536 24216
rect 7932 24200 7984 24206
rect 7932 24142 7984 24148
rect 8024 24200 8076 24206
rect 8024 24142 8076 24148
rect 7840 24064 7892 24070
rect 7840 24006 7892 24012
rect 7852 23866 7880 24006
rect 7656 23860 7708 23866
rect 7656 23802 7708 23808
rect 7840 23860 7892 23866
rect 7840 23802 7892 23808
rect 7288 23724 7340 23730
rect 7288 23666 7340 23672
rect 7564 23724 7616 23730
rect 7564 23666 7616 23672
rect 7196 23112 7248 23118
rect 7196 23054 7248 23060
rect 7208 22642 7236 23054
rect 7300 22778 7328 23666
rect 7656 23656 7708 23662
rect 7656 23598 7708 23604
rect 7564 23248 7616 23254
rect 7564 23190 7616 23196
rect 7576 23050 7604 23190
rect 7668 23118 7696 23598
rect 7852 23186 7880 23802
rect 7944 23662 7972 24142
rect 7932 23656 7984 23662
rect 7932 23598 7984 23604
rect 7944 23254 7972 23598
rect 8024 23588 8076 23594
rect 8024 23530 8076 23536
rect 7932 23248 7984 23254
rect 7932 23190 7984 23196
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7656 23112 7708 23118
rect 7656 23054 7708 23060
rect 7564 23044 7616 23050
rect 7564 22986 7616 22992
rect 7288 22772 7340 22778
rect 7288 22714 7340 22720
rect 7196 22636 7248 22642
rect 7472 22636 7524 22642
rect 7248 22596 7328 22624
rect 7196 22578 7248 22584
rect 7300 21962 7328 22596
rect 7472 22578 7524 22584
rect 7484 22438 7512 22578
rect 7472 22432 7524 22438
rect 7472 22374 7524 22380
rect 7484 22166 7512 22374
rect 7472 22160 7524 22166
rect 7472 22102 7524 22108
rect 7380 22092 7432 22098
rect 7380 22034 7432 22040
rect 7288 21956 7340 21962
rect 7288 21898 7340 21904
rect 7196 21548 7248 21554
rect 7196 21490 7248 21496
rect 7208 21350 7236 21490
rect 7196 21344 7248 21350
rect 7196 21286 7248 21292
rect 7300 21162 7328 21898
rect 7392 21690 7420 22034
rect 7576 21865 7604 22986
rect 7668 22982 7696 23054
rect 7656 22976 7708 22982
rect 7656 22918 7708 22924
rect 7852 22488 7880 23122
rect 8036 23118 8064 23530
rect 8128 23118 8156 24210
rect 8300 24064 8352 24070
rect 8300 24006 8352 24012
rect 8208 23792 8260 23798
rect 8208 23734 8260 23740
rect 8024 23112 8076 23118
rect 8024 23054 8076 23060
rect 8116 23112 8168 23118
rect 8116 23054 8168 23060
rect 8024 22772 8076 22778
rect 8024 22714 8076 22720
rect 7932 22500 7984 22506
rect 7852 22460 7932 22488
rect 7932 22442 7984 22448
rect 7944 22080 7972 22442
rect 7852 22052 7972 22080
rect 7656 22024 7708 22030
rect 7656 21966 7708 21972
rect 7562 21856 7618 21865
rect 7562 21791 7618 21800
rect 7562 21720 7618 21729
rect 7380 21684 7432 21690
rect 7668 21690 7696 21966
rect 7562 21655 7618 21664
rect 7656 21684 7708 21690
rect 7380 21626 7432 21632
rect 7472 21616 7524 21622
rect 7470 21584 7472 21593
rect 7524 21584 7526 21593
rect 7470 21519 7526 21528
rect 7472 21480 7524 21486
rect 7472 21422 7524 21428
rect 7380 21344 7432 21350
rect 7380 21286 7432 21292
rect 7208 21134 7328 21162
rect 7208 20806 7236 21134
rect 7288 21004 7340 21010
rect 7288 20946 7340 20952
rect 7196 20800 7248 20806
rect 7196 20742 7248 20748
rect 7194 20632 7250 20641
rect 7194 20567 7250 20576
rect 7208 14498 7236 20567
rect 7300 20369 7328 20946
rect 7286 20360 7342 20369
rect 7286 20295 7342 20304
rect 7300 19514 7328 20295
rect 7392 19786 7420 21286
rect 7484 20942 7512 21422
rect 7472 20936 7524 20942
rect 7472 20878 7524 20884
rect 7484 20330 7512 20878
rect 7576 20806 7604 21655
rect 7656 21626 7708 21632
rect 7852 21554 7880 22052
rect 7930 21856 7986 21865
rect 7930 21791 7986 21800
rect 7748 21548 7800 21554
rect 7748 21490 7800 21496
rect 7840 21548 7892 21554
rect 7840 21490 7892 21496
rect 7656 21140 7708 21146
rect 7656 21082 7708 21088
rect 7564 20800 7616 20806
rect 7564 20742 7616 20748
rect 7668 20466 7696 21082
rect 7564 20460 7616 20466
rect 7564 20402 7616 20408
rect 7656 20460 7708 20466
rect 7656 20402 7708 20408
rect 7472 20324 7524 20330
rect 7472 20266 7524 20272
rect 7380 19780 7432 19786
rect 7380 19722 7432 19728
rect 7472 19712 7524 19718
rect 7378 19680 7434 19689
rect 7472 19654 7524 19660
rect 7378 19615 7434 19624
rect 7288 19508 7340 19514
rect 7288 19450 7340 19456
rect 7288 19236 7340 19242
rect 7288 19178 7340 19184
rect 7300 19145 7328 19178
rect 7286 19136 7342 19145
rect 7286 19071 7342 19080
rect 7288 18760 7340 18766
rect 7288 18702 7340 18708
rect 7300 18426 7328 18702
rect 7288 18420 7340 18426
rect 7288 18362 7340 18368
rect 7392 17105 7420 19615
rect 7378 17096 7434 17105
rect 7378 17031 7434 17040
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7392 15910 7420 16934
rect 7484 16130 7512 19654
rect 7576 19310 7604 20402
rect 7668 20058 7696 20402
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7656 19916 7708 19922
rect 7656 19858 7708 19864
rect 7564 19304 7616 19310
rect 7564 19246 7616 19252
rect 7576 18834 7604 19246
rect 7564 18828 7616 18834
rect 7564 18770 7616 18776
rect 7564 16584 7616 16590
rect 7564 16526 7616 16532
rect 7576 16250 7604 16526
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7484 16102 7604 16130
rect 7380 15904 7432 15910
rect 7380 15846 7432 15852
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 7208 14470 7328 14498
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7208 12345 7236 14350
rect 7194 12336 7250 12345
rect 7194 12271 7250 12280
rect 7194 12064 7250 12073
rect 7194 11999 7250 12008
rect 7208 5234 7236 11999
rect 7300 7562 7328 14470
rect 7392 12730 7420 15642
rect 7472 15632 7524 15638
rect 7472 15574 7524 15580
rect 7484 12986 7512 15574
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7392 12702 7512 12730
rect 7380 12640 7432 12646
rect 7378 12608 7380 12617
rect 7432 12608 7434 12617
rect 7378 12543 7434 12552
rect 7378 12472 7434 12481
rect 7378 12407 7434 12416
rect 7392 12345 7420 12407
rect 7378 12336 7434 12345
rect 7378 12271 7434 12280
rect 7380 10668 7432 10674
rect 7380 10610 7432 10616
rect 7392 8022 7420 10610
rect 7484 10554 7512 12702
rect 7576 10674 7604 16102
rect 7668 15638 7696 19858
rect 7656 15632 7708 15638
rect 7656 15574 7708 15580
rect 7760 14414 7788 21490
rect 7852 20466 7880 21490
rect 7944 20942 7972 21791
rect 7932 20936 7984 20942
rect 7932 20878 7984 20884
rect 7840 20460 7892 20466
rect 7840 20402 7892 20408
rect 7944 19961 7972 20878
rect 8036 20874 8064 22714
rect 8220 22574 8248 23734
rect 8312 22778 8340 24006
rect 8392 23792 8444 23798
rect 8392 23734 8444 23740
rect 8300 22772 8352 22778
rect 8300 22714 8352 22720
rect 8208 22568 8260 22574
rect 8208 22510 8260 22516
rect 8116 22432 8168 22438
rect 8116 22374 8168 22380
rect 8128 21554 8156 22374
rect 8404 22250 8432 23734
rect 8496 23526 8524 24210
rect 8484 23520 8536 23526
rect 8484 23462 8536 23468
rect 8484 23248 8536 23254
rect 8484 23190 8536 23196
rect 8220 22234 8432 22250
rect 8208 22228 8432 22234
rect 8260 22222 8432 22228
rect 8208 22170 8260 22176
rect 8300 22024 8352 22030
rect 8300 21966 8352 21972
rect 8312 21865 8340 21966
rect 8298 21856 8354 21865
rect 8298 21791 8354 21800
rect 8116 21548 8168 21554
rect 8116 21490 8168 21496
rect 8404 21146 8432 22222
rect 8496 21894 8524 23190
rect 8588 23050 8616 26930
rect 8680 26790 8708 27367
rect 8668 26784 8720 26790
rect 8668 26726 8720 26732
rect 8668 26308 8720 26314
rect 8668 26250 8720 26256
rect 8680 26042 8708 26250
rect 8668 26036 8720 26042
rect 8668 25978 8720 25984
rect 8772 24818 8800 28426
rect 9140 27402 9168 28630
rect 10508 28552 10560 28558
rect 10508 28494 10560 28500
rect 11336 28552 11388 28558
rect 11336 28494 11388 28500
rect 10416 28416 10468 28422
rect 10416 28358 10468 28364
rect 9935 28316 10243 28336
rect 9935 28314 9941 28316
rect 9997 28314 10021 28316
rect 10077 28314 10101 28316
rect 10157 28314 10181 28316
rect 10237 28314 10243 28316
rect 9997 28262 9999 28314
rect 10179 28262 10181 28314
rect 9935 28260 9941 28262
rect 9997 28260 10021 28262
rect 10077 28260 10101 28262
rect 10157 28260 10181 28262
rect 10237 28260 10243 28262
rect 9935 28240 10243 28260
rect 9680 28144 9732 28150
rect 9680 28086 9732 28092
rect 9220 27872 9272 27878
rect 9220 27814 9272 27820
rect 9128 27396 9180 27402
rect 9128 27338 9180 27344
rect 9232 26994 9260 27814
rect 9692 27674 9720 28086
rect 9864 28076 9916 28082
rect 9864 28018 9916 28024
rect 9680 27668 9732 27674
rect 9680 27610 9732 27616
rect 9220 26988 9272 26994
rect 9220 26930 9272 26936
rect 9404 26988 9456 26994
rect 9404 26930 9456 26936
rect 8852 25900 8904 25906
rect 8852 25842 8904 25848
rect 8864 25770 8892 25842
rect 8852 25764 8904 25770
rect 8852 25706 8904 25712
rect 9416 25294 9444 26930
rect 9680 26784 9732 26790
rect 9680 26726 9732 26732
rect 9692 25906 9720 26726
rect 9876 26586 9904 28018
rect 10324 27328 10376 27334
rect 10324 27270 10376 27276
rect 9935 27228 10243 27248
rect 9935 27226 9941 27228
rect 9997 27226 10021 27228
rect 10077 27226 10101 27228
rect 10157 27226 10181 27228
rect 10237 27226 10243 27228
rect 9997 27174 9999 27226
rect 10179 27174 10181 27226
rect 9935 27172 9941 27174
rect 9997 27172 10021 27174
rect 10077 27172 10101 27174
rect 10157 27172 10181 27174
rect 10237 27172 10243 27174
rect 9935 27152 10243 27172
rect 9864 26580 9916 26586
rect 9864 26522 9916 26528
rect 10048 26580 10100 26586
rect 10048 26522 10100 26528
rect 10060 26450 10088 26522
rect 10336 26518 10364 27270
rect 10324 26512 10376 26518
rect 10324 26454 10376 26460
rect 10048 26444 10100 26450
rect 10048 26386 10100 26392
rect 9772 26240 9824 26246
rect 9772 26182 9824 26188
rect 9588 25900 9640 25906
rect 9588 25842 9640 25848
rect 9680 25900 9732 25906
rect 9680 25842 9732 25848
rect 9600 25498 9628 25842
rect 9588 25492 9640 25498
rect 9588 25434 9640 25440
rect 9404 25288 9456 25294
rect 9404 25230 9456 25236
rect 9312 24948 9364 24954
rect 9312 24890 9364 24896
rect 8760 24812 8812 24818
rect 8812 24772 8892 24800
rect 8760 24754 8812 24760
rect 8864 23254 8892 24772
rect 9036 24200 9088 24206
rect 9036 24142 9088 24148
rect 8944 23860 8996 23866
rect 8944 23802 8996 23808
rect 8956 23662 8984 23802
rect 9048 23798 9076 24142
rect 9220 23860 9272 23866
rect 9220 23802 9272 23808
rect 9036 23792 9088 23798
rect 9036 23734 9088 23740
rect 9128 23792 9180 23798
rect 9128 23734 9180 23740
rect 9140 23662 9168 23734
rect 8944 23656 8996 23662
rect 8944 23598 8996 23604
rect 9128 23656 9180 23662
rect 9128 23598 9180 23604
rect 9036 23520 9088 23526
rect 9036 23462 9088 23468
rect 8852 23248 8904 23254
rect 8852 23190 8904 23196
rect 9048 23050 9076 23462
rect 9232 23186 9260 23802
rect 9324 23662 9352 24890
rect 9312 23656 9364 23662
rect 9312 23598 9364 23604
rect 9220 23180 9272 23186
rect 9220 23122 9272 23128
rect 8576 23044 8628 23050
rect 8576 22986 8628 22992
rect 8852 23044 8904 23050
rect 8852 22986 8904 22992
rect 9036 23044 9088 23050
rect 9036 22986 9088 22992
rect 8576 22568 8628 22574
rect 8576 22510 8628 22516
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8496 21554 8524 21830
rect 8588 21622 8616 22510
rect 8668 22432 8720 22438
rect 8668 22374 8720 22380
rect 8680 22234 8708 22374
rect 8668 22228 8720 22234
rect 8668 22170 8720 22176
rect 8668 21956 8720 21962
rect 8668 21898 8720 21904
rect 8576 21616 8628 21622
rect 8576 21558 8628 21564
rect 8484 21548 8536 21554
rect 8484 21490 8536 21496
rect 8680 21418 8708 21898
rect 8668 21412 8720 21418
rect 8668 21354 8720 21360
rect 8392 21140 8444 21146
rect 8392 21082 8444 21088
rect 8024 20868 8076 20874
rect 8024 20810 8076 20816
rect 8036 20534 8064 20810
rect 8666 20632 8722 20641
rect 8864 20602 8892 22986
rect 8944 22024 8996 22030
rect 8944 21966 8996 21972
rect 8956 21865 8984 21966
rect 8942 21856 8998 21865
rect 8942 21791 8998 21800
rect 8956 21622 8984 21791
rect 8944 21616 8996 21622
rect 8944 21558 8996 21564
rect 8944 20936 8996 20942
rect 8944 20878 8996 20884
rect 8666 20567 8722 20576
rect 8852 20596 8904 20602
rect 8024 20528 8076 20534
rect 8024 20470 8076 20476
rect 8116 20052 8168 20058
rect 8116 19994 8168 20000
rect 8128 19961 8156 19994
rect 8484 19984 8536 19990
rect 7930 19952 7986 19961
rect 7930 19887 7986 19896
rect 8114 19952 8170 19961
rect 8484 19926 8536 19932
rect 8114 19887 8170 19896
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8300 19508 8352 19514
rect 7852 19468 8300 19496
rect 7852 19378 7880 19468
rect 8300 19450 8352 19456
rect 8114 19408 8170 19417
rect 7840 19372 7892 19378
rect 8404 19394 8432 19654
rect 8114 19343 8116 19352
rect 7840 19314 7892 19320
rect 8168 19343 8170 19352
rect 8220 19366 8432 19394
rect 8116 19314 8168 19320
rect 8220 19258 8248 19366
rect 8392 19304 8444 19310
rect 8128 19230 8248 19258
rect 8312 19264 8392 19292
rect 8128 19174 8156 19230
rect 8116 19168 8168 19174
rect 8116 19110 8168 19116
rect 7838 19000 7894 19009
rect 7838 18935 7894 18944
rect 7852 15706 7880 18935
rect 8206 18592 8262 18601
rect 8206 18527 8262 18536
rect 7930 18456 7986 18465
rect 7930 18391 7932 18400
rect 7984 18391 7986 18400
rect 7932 18362 7984 18368
rect 8022 18320 8078 18329
rect 8022 18255 8078 18264
rect 7932 16176 7984 16182
rect 7932 16118 7984 16124
rect 7944 15706 7972 16118
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7840 15564 7892 15570
rect 7840 15506 7892 15512
rect 7852 14906 7880 15506
rect 7930 15056 7986 15065
rect 7930 14991 7932 15000
rect 7984 14991 7986 15000
rect 7932 14962 7984 14968
rect 7852 14878 7972 14906
rect 7840 14816 7892 14822
rect 7840 14758 7892 14764
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7654 12472 7710 12481
rect 7760 12442 7788 13874
rect 7852 12753 7880 14758
rect 7944 13297 7972 14878
rect 7930 13288 7986 13297
rect 7930 13223 7986 13232
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 7944 12850 7972 13126
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7838 12744 7894 12753
rect 8036 12730 8064 18255
rect 8220 16538 8248 18527
rect 8312 17882 8340 19264
rect 8496 19292 8524 19926
rect 8576 19916 8628 19922
rect 8576 19858 8628 19864
rect 8444 19264 8524 19292
rect 8392 19246 8444 19252
rect 8588 19242 8616 19858
rect 8680 19553 8708 20567
rect 8852 20538 8904 20544
rect 8852 20324 8904 20330
rect 8852 20266 8904 20272
rect 8666 19544 8722 19553
rect 8666 19479 8722 19488
rect 8576 19236 8628 19242
rect 8576 19178 8628 19184
rect 8482 19136 8538 19145
rect 8482 19071 8538 19080
rect 8496 18970 8524 19071
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8312 17202 8340 17682
rect 8588 17610 8616 19178
rect 8680 17678 8708 19479
rect 8758 19272 8814 19281
rect 8758 19207 8814 19216
rect 8772 18086 8800 19207
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8576 17604 8628 17610
rect 8576 17546 8628 17552
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 8588 17134 8616 17546
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 7838 12679 7894 12688
rect 7944 12702 8064 12730
rect 8128 16510 8248 16538
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7654 12407 7710 12416
rect 7748 12436 7800 12442
rect 7668 11830 7696 12407
rect 7748 12378 7800 12384
rect 7746 12336 7802 12345
rect 7746 12271 7802 12280
rect 7656 11824 7708 11830
rect 7656 11766 7708 11772
rect 7656 11144 7708 11150
rect 7654 11112 7656 11121
rect 7708 11112 7710 11121
rect 7654 11047 7710 11056
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7668 10674 7696 10950
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 7484 10526 7696 10554
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7380 8016 7432 8022
rect 7380 7958 7432 7964
rect 7300 7534 7420 7562
rect 7286 7440 7342 7449
rect 7286 7375 7342 7384
rect 7300 5846 7328 7375
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7300 5409 7328 5510
rect 7286 5400 7342 5409
rect 7286 5335 7342 5344
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 7208 4010 7236 5034
rect 7196 4004 7248 4010
rect 7196 3946 7248 3952
rect 7300 3738 7328 5238
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7300 3194 7328 3470
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7208 2650 7236 3130
rect 7392 3126 7420 7534
rect 7484 5098 7512 10406
rect 7576 10062 7604 10406
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7576 9654 7604 9862
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 7576 9110 7604 9590
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7562 8528 7618 8537
rect 7562 8463 7618 8472
rect 7576 5370 7604 8463
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7472 5092 7524 5098
rect 7472 5034 7524 5040
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7484 3738 7512 4626
rect 7576 3942 7604 5170
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7564 3460 7616 3466
rect 7564 3402 7616 3408
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7378 2952 7434 2961
rect 7378 2887 7434 2896
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7392 800 7420 2887
rect 7576 2854 7604 3402
rect 7564 2848 7616 2854
rect 7564 2790 7616 2796
rect 7668 800 7696 10526
rect 7760 7478 7788 12271
rect 7852 9994 7880 12582
rect 7840 9988 7892 9994
rect 7840 9930 7892 9936
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 7852 7410 7880 9522
rect 7944 8090 7972 12702
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 8036 12374 8064 12582
rect 8024 12368 8076 12374
rect 8024 12310 8076 12316
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7746 7304 7802 7313
rect 7746 7239 7802 7248
rect 7760 6866 7788 7239
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7852 5250 7880 6734
rect 7760 5222 7880 5250
rect 7760 4282 7788 5222
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7852 4146 7880 5102
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 7760 3738 7788 4082
rect 7840 4004 7892 4010
rect 7840 3946 7892 3952
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7852 3602 7880 3946
rect 7840 3596 7892 3602
rect 7944 3584 7972 7686
rect 8036 4826 8064 12038
rect 8128 11014 8156 16510
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 8220 15910 8248 16390
rect 8404 16250 8432 16526
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8680 16182 8708 17614
rect 8668 16176 8720 16182
rect 8668 16118 8720 16124
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8312 15162 8340 15302
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8496 15116 8708 15144
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 8220 14278 8248 14962
rect 8312 14958 8340 15098
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8312 14006 8340 14894
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 8404 13938 8432 14418
rect 8496 14006 8524 15116
rect 8574 15056 8630 15065
rect 8680 15026 8708 15116
rect 8574 14991 8630 15000
rect 8668 15020 8720 15026
rect 8484 14000 8536 14006
rect 8484 13942 8536 13948
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 8220 12152 8248 13738
rect 8404 12850 8432 13874
rect 8496 13530 8524 13942
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8496 12986 8524 13262
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8588 12889 8616 14991
rect 8668 14962 8720 14968
rect 8864 14793 8892 20266
rect 8956 19922 8984 20878
rect 9036 20800 9088 20806
rect 9088 20760 9168 20788
rect 9036 20742 9088 20748
rect 9036 20528 9088 20534
rect 9036 20470 9088 20476
rect 8944 19916 8996 19922
rect 8944 19858 8996 19864
rect 9048 19786 9076 20470
rect 9036 19780 9088 19786
rect 8956 19740 9036 19768
rect 8956 18850 8984 19740
rect 9036 19722 9088 19728
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 9048 18970 9076 19314
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 8956 18822 9076 18850
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 8956 16658 8984 17614
rect 8944 16652 8996 16658
rect 8944 16594 8996 16600
rect 8956 16114 8984 16594
rect 8944 16108 8996 16114
rect 8944 16050 8996 16056
rect 8850 14784 8906 14793
rect 8850 14719 8906 14728
rect 9048 14618 9076 18822
rect 9140 18306 9168 20760
rect 9232 20466 9260 23122
rect 9324 23118 9352 23598
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 9220 20460 9272 20466
rect 9220 20402 9272 20408
rect 9324 20262 9352 23054
rect 9416 22642 9444 25230
rect 9600 24818 9628 25434
rect 9588 24812 9640 24818
rect 9588 24754 9640 24760
rect 9692 24750 9720 25842
rect 9784 24954 9812 26182
rect 9935 26140 10243 26160
rect 9935 26138 9941 26140
rect 9997 26138 10021 26140
rect 10077 26138 10101 26140
rect 10157 26138 10181 26140
rect 10237 26138 10243 26140
rect 9997 26086 9999 26138
rect 10179 26086 10181 26138
rect 9935 26084 9941 26086
rect 9997 26084 10021 26086
rect 10077 26084 10101 26086
rect 10157 26084 10181 26086
rect 10237 26084 10243 26086
rect 9935 26064 10243 26084
rect 9864 25696 9916 25702
rect 9864 25638 9916 25644
rect 9772 24948 9824 24954
rect 9772 24890 9824 24896
rect 9680 24744 9732 24750
rect 9680 24686 9732 24692
rect 9588 24064 9640 24070
rect 9588 24006 9640 24012
rect 9600 23730 9628 24006
rect 9588 23724 9640 23730
rect 9588 23666 9640 23672
rect 9600 23118 9628 23666
rect 9784 23168 9812 24890
rect 9876 24682 9904 25638
rect 10336 25430 10364 26454
rect 10428 26382 10456 28358
rect 10416 26376 10468 26382
rect 10416 26318 10468 26324
rect 10416 26240 10468 26246
rect 10416 26182 10468 26188
rect 10324 25424 10376 25430
rect 10324 25366 10376 25372
rect 9935 25052 10243 25072
rect 9935 25050 9941 25052
rect 9997 25050 10021 25052
rect 10077 25050 10101 25052
rect 10157 25050 10181 25052
rect 10237 25050 10243 25052
rect 9997 24998 9999 25050
rect 10179 24998 10181 25050
rect 9935 24996 9941 24998
rect 9997 24996 10021 24998
rect 10077 24996 10101 24998
rect 10157 24996 10181 24998
rect 10237 24996 10243 24998
rect 9935 24976 10243 24996
rect 10336 24818 10364 25366
rect 10324 24812 10376 24818
rect 10324 24754 10376 24760
rect 9864 24676 9916 24682
rect 9864 24618 9916 24624
rect 9864 24268 9916 24274
rect 9864 24210 9916 24216
rect 9692 23140 9812 23168
rect 9588 23112 9640 23118
rect 9588 23054 9640 23060
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9496 22500 9548 22506
rect 9496 22442 9548 22448
rect 9402 22128 9458 22137
rect 9402 22063 9458 22072
rect 9416 21554 9444 22063
rect 9404 21548 9456 21554
rect 9404 21490 9456 21496
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 9508 19854 9536 22442
rect 9692 22030 9720 23140
rect 9876 23118 9904 24210
rect 10428 24206 10456 26182
rect 9956 24200 10008 24206
rect 10140 24200 10192 24206
rect 10008 24160 10140 24188
rect 9956 24142 10008 24148
rect 10140 24142 10192 24148
rect 10416 24200 10468 24206
rect 10416 24142 10468 24148
rect 9935 23964 10243 23984
rect 9935 23962 9941 23964
rect 9997 23962 10021 23964
rect 10077 23962 10101 23964
rect 10157 23962 10181 23964
rect 10237 23962 10243 23964
rect 9997 23910 9999 23962
rect 10179 23910 10181 23962
rect 9935 23908 9941 23910
rect 9997 23908 10021 23910
rect 10077 23908 10101 23910
rect 10157 23908 10181 23910
rect 10237 23908 10243 23910
rect 9935 23888 10243 23908
rect 10416 23792 10468 23798
rect 10416 23734 10468 23740
rect 10232 23656 10284 23662
rect 10284 23616 10364 23644
rect 10232 23598 10284 23604
rect 9864 23112 9916 23118
rect 9864 23054 9916 23060
rect 9935 22876 10243 22896
rect 9935 22874 9941 22876
rect 9997 22874 10021 22876
rect 10077 22874 10101 22876
rect 10157 22874 10181 22876
rect 10237 22874 10243 22876
rect 9997 22822 9999 22874
rect 10179 22822 10181 22874
rect 9935 22820 9941 22822
rect 9997 22820 10021 22822
rect 10077 22820 10101 22822
rect 10157 22820 10181 22822
rect 10237 22820 10243 22822
rect 9935 22800 10243 22820
rect 9864 22772 9916 22778
rect 10336 22760 10364 23616
rect 9864 22714 9916 22720
rect 10152 22732 10364 22760
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 9784 22098 9812 22578
rect 9772 22092 9824 22098
rect 9772 22034 9824 22040
rect 9680 22024 9732 22030
rect 9680 21966 9732 21972
rect 9588 21616 9640 21622
rect 9588 21558 9640 21564
rect 9600 21486 9628 21558
rect 9692 21486 9720 21966
rect 9588 21480 9640 21486
rect 9588 21422 9640 21428
rect 9680 21480 9732 21486
rect 9784 21457 9812 22034
rect 9876 21554 9904 22714
rect 10152 22166 10180 22732
rect 10324 22636 10376 22642
rect 10324 22578 10376 22584
rect 10232 22568 10284 22574
rect 10232 22510 10284 22516
rect 10140 22160 10192 22166
rect 10140 22102 10192 22108
rect 10244 22030 10272 22510
rect 10336 22098 10364 22578
rect 10428 22574 10456 23734
rect 10520 23474 10548 28494
rect 10968 28416 11020 28422
rect 11152 28416 11204 28422
rect 11020 28376 11100 28404
rect 10968 28358 11020 28364
rect 10968 28008 11020 28014
rect 10968 27950 11020 27956
rect 10692 27872 10744 27878
rect 10692 27814 10744 27820
rect 10704 26994 10732 27814
rect 10980 27674 11008 27950
rect 10968 27668 11020 27674
rect 10968 27610 11020 27616
rect 10980 27470 11008 27610
rect 10968 27464 11020 27470
rect 10968 27406 11020 27412
rect 10876 27056 10928 27062
rect 10876 26998 10928 27004
rect 10692 26988 10744 26994
rect 10692 26930 10744 26936
rect 10600 26920 10652 26926
rect 10600 26862 10652 26868
rect 10612 26382 10640 26862
rect 10888 26489 10916 26998
rect 10874 26480 10930 26489
rect 10874 26415 10930 26424
rect 10600 26376 10652 26382
rect 10600 26318 10652 26324
rect 10876 26376 10928 26382
rect 10876 26318 10928 26324
rect 10612 23662 10640 26318
rect 10784 26240 10836 26246
rect 10784 26182 10836 26188
rect 10796 25974 10824 26182
rect 10888 26042 10916 26318
rect 10876 26036 10928 26042
rect 10876 25978 10928 25984
rect 10784 25968 10836 25974
rect 10784 25910 10836 25916
rect 10980 25294 11008 27406
rect 10968 25288 11020 25294
rect 10968 25230 11020 25236
rect 10876 25220 10928 25226
rect 10876 25162 10928 25168
rect 10888 24954 10916 25162
rect 10968 25152 11020 25158
rect 10968 25094 11020 25100
rect 10876 24948 10928 24954
rect 10876 24890 10928 24896
rect 10784 24812 10836 24818
rect 10784 24754 10836 24760
rect 10876 24812 10928 24818
rect 10876 24754 10928 24760
rect 10692 24744 10744 24750
rect 10692 24686 10744 24692
rect 10600 23656 10652 23662
rect 10600 23598 10652 23604
rect 10520 23446 10640 23474
rect 10508 23180 10560 23186
rect 10508 23122 10560 23128
rect 10416 22568 10468 22574
rect 10416 22510 10468 22516
rect 10414 22128 10470 22137
rect 10324 22092 10376 22098
rect 10414 22063 10416 22072
rect 10324 22034 10376 22040
rect 10468 22063 10470 22072
rect 10416 22034 10468 22040
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 9935 21788 10243 21808
rect 9935 21786 9941 21788
rect 9997 21786 10021 21788
rect 10077 21786 10101 21788
rect 10157 21786 10181 21788
rect 10237 21786 10243 21788
rect 9997 21734 9999 21786
rect 10179 21734 10181 21786
rect 9935 21732 9941 21734
rect 9997 21732 10021 21734
rect 10077 21732 10101 21734
rect 10157 21732 10181 21734
rect 10237 21732 10243 21734
rect 9935 21712 10243 21732
rect 10336 21570 10364 22034
rect 10416 21684 10468 21690
rect 10416 21626 10468 21632
rect 9864 21548 9916 21554
rect 9864 21490 9916 21496
rect 10152 21542 10364 21570
rect 9680 21422 9732 21428
rect 9770 21448 9826 21457
rect 9770 21383 9826 21392
rect 9680 21344 9732 21350
rect 9680 21286 9732 21292
rect 9864 21344 9916 21350
rect 9864 21286 9916 21292
rect 9692 20942 9720 21286
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 9680 20936 9732 20942
rect 9876 20890 9904 21286
rect 10152 21078 10180 21542
rect 10322 21448 10378 21457
rect 10322 21383 10378 21392
rect 10336 21078 10364 21383
rect 10140 21072 10192 21078
rect 10140 21014 10192 21020
rect 10324 21072 10376 21078
rect 10324 21014 10376 21020
rect 9956 20936 10008 20942
rect 9680 20878 9732 20884
rect 9600 20534 9628 20878
rect 9784 20862 9904 20890
rect 9954 20904 9956 20913
rect 10008 20904 10010 20913
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9588 20528 9640 20534
rect 9588 20470 9640 20476
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 9600 19446 9628 19790
rect 9588 19440 9640 19446
rect 9588 19382 9640 19388
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 9140 18278 9444 18306
rect 9508 18290 9536 18566
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 9232 17202 9260 18158
rect 9416 18034 9444 18278
rect 9496 18284 9548 18290
rect 9496 18226 9548 18232
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9416 18006 9536 18034
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9128 15904 9180 15910
rect 9128 15846 9180 15852
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8680 14074 8708 14350
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8680 13462 8708 14010
rect 8864 13734 8892 14554
rect 8852 13728 8904 13734
rect 8852 13670 8904 13676
rect 8668 13456 8720 13462
rect 8668 13398 8720 13404
rect 8574 12880 8630 12889
rect 8392 12844 8444 12850
rect 8574 12815 8630 12824
rect 8392 12786 8444 12792
rect 8404 12646 8432 12786
rect 8680 12646 8708 13398
rect 8864 12782 8892 13670
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 9048 12832 9076 13194
rect 9140 13161 9168 15846
rect 9232 15638 9260 17138
rect 9416 16182 9444 17818
rect 9404 16176 9456 16182
rect 9404 16118 9456 16124
rect 9220 15632 9272 15638
rect 9220 15574 9272 15580
rect 9232 15162 9260 15574
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9508 14498 9536 18006
rect 9600 17785 9628 18226
rect 9586 17776 9642 17785
rect 9586 17711 9642 17720
rect 9588 17604 9640 17610
rect 9588 17546 9640 17552
rect 9600 17338 9628 17546
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9692 16998 9720 20742
rect 9784 20641 9812 20862
rect 9954 20839 10010 20848
rect 9935 20700 10243 20720
rect 9935 20698 9941 20700
rect 9997 20698 10021 20700
rect 10077 20698 10101 20700
rect 10157 20698 10181 20700
rect 10237 20698 10243 20700
rect 9997 20646 9999 20698
rect 10179 20646 10181 20698
rect 9935 20644 9941 20646
rect 9997 20644 10021 20646
rect 10077 20644 10101 20646
rect 10157 20644 10181 20646
rect 10237 20644 10243 20646
rect 9770 20632 9826 20641
rect 9935 20624 10243 20644
rect 9770 20567 9826 20576
rect 9772 20460 9824 20466
rect 9772 20402 9824 20408
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9588 16516 9640 16522
rect 9588 16458 9640 16464
rect 9600 15502 9628 16458
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9692 15144 9720 16526
rect 9416 14470 9536 14498
rect 9600 15116 9720 15144
rect 9126 13152 9182 13161
rect 9126 13087 9182 13096
rect 9218 13016 9274 13025
rect 9218 12951 9274 12960
rect 9232 12850 9260 12951
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 9128 12844 9180 12850
rect 9048 12804 9128 12832
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8392 12640 8444 12646
rect 8392 12582 8444 12588
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8850 12608 8906 12617
rect 8300 12164 8352 12170
rect 8220 12124 8300 12152
rect 8300 12106 8352 12112
rect 8404 12102 8432 12582
rect 8850 12543 8906 12552
rect 8666 12472 8722 12481
rect 8588 12416 8666 12434
rect 8864 12434 8892 12543
rect 9048 12458 9076 12804
rect 9128 12786 9180 12792
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 8588 12407 8722 12416
rect 8588 12406 8708 12407
rect 8772 12406 8892 12434
rect 9039 12430 9076 12458
rect 8392 12096 8444 12102
rect 8206 12064 8262 12073
rect 8392 12038 8444 12044
rect 8206 11999 8262 12008
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 8128 10266 8156 10610
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 8128 9897 8156 10066
rect 8114 9888 8170 9897
rect 8114 9823 8170 9832
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8128 7970 8156 9658
rect 8220 8090 8248 11999
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8404 11014 8432 11494
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8404 10606 8432 10950
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8312 9518 8340 9998
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8496 9586 8524 9862
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8392 9444 8444 9450
rect 8392 9386 8444 9392
rect 8404 8906 8432 9386
rect 8496 8906 8524 9522
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8312 8362 8340 8774
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 8128 7942 8248 7970
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 8022 4720 8078 4729
rect 8022 4655 8078 4664
rect 8036 4282 8064 4655
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 8024 3596 8076 3602
rect 7944 3556 8024 3584
rect 7840 3538 7892 3544
rect 8024 3538 8076 3544
rect 7852 2446 7880 3538
rect 7932 3120 7984 3126
rect 7932 3062 7984 3068
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 7944 800 7972 3062
rect 8128 2774 8156 7822
rect 8220 7426 8248 7942
rect 8220 7398 8340 7426
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8220 6798 8248 7278
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8220 5030 8248 6054
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 8312 4842 8340 7398
rect 8220 4814 8340 4842
rect 8220 4282 8248 4814
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8220 3058 8248 4082
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8128 2746 8248 2774
rect 8220 800 8248 2746
rect 8312 2650 8340 4694
rect 8404 3398 8432 8434
rect 8496 6390 8524 8842
rect 8484 6384 8536 6390
rect 8484 6326 8536 6332
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8496 5778 8524 6190
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8484 5636 8536 5642
rect 8484 5578 8536 5584
rect 8496 4758 8524 5578
rect 8484 4752 8536 4758
rect 8484 4694 8536 4700
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 8496 3126 8524 3606
rect 8484 3120 8536 3126
rect 8484 3062 8536 3068
rect 8588 2774 8616 12406
rect 8666 12336 8722 12345
rect 8666 12271 8722 12280
rect 8680 8498 8708 12271
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8404 2746 8616 2774
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8404 800 8432 2746
rect 8680 800 8708 8230
rect 8772 5574 8800 12406
rect 8944 12368 8996 12374
rect 9039 12356 9067 12430
rect 9039 12328 9076 12356
rect 8944 12310 8996 12316
rect 8852 12164 8904 12170
rect 8852 12106 8904 12112
rect 8864 11150 8892 12106
rect 8956 11150 8984 12310
rect 9048 11898 9076 12328
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 9048 11098 9076 11698
rect 9324 11354 9352 12854
rect 9416 12617 9444 14470
rect 9496 14340 9548 14346
rect 9496 14282 9548 14288
rect 9508 12714 9536 14282
rect 9496 12708 9548 12714
rect 9496 12650 9548 12656
rect 9402 12608 9458 12617
rect 9402 12543 9458 12552
rect 9402 12472 9458 12481
rect 9402 12407 9458 12416
rect 9416 11762 9444 12407
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9508 11370 9536 12650
rect 9600 12345 9628 15116
rect 9784 15094 9812 20402
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 9864 19780 9916 19786
rect 9864 19722 9916 19728
rect 9772 15088 9824 15094
rect 9772 15030 9824 15036
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9692 14822 9720 14962
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9692 13326 9720 14758
rect 9784 14618 9812 15030
rect 9876 14890 9904 19722
rect 9935 19612 10243 19632
rect 9935 19610 9941 19612
rect 9997 19610 10021 19612
rect 10077 19610 10101 19612
rect 10157 19610 10181 19612
rect 10237 19610 10243 19612
rect 9997 19558 9999 19610
rect 10179 19558 10181 19610
rect 9935 19556 9941 19558
rect 9997 19556 10021 19558
rect 10077 19556 10101 19558
rect 10157 19556 10181 19558
rect 10237 19556 10243 19558
rect 9935 19536 10243 19556
rect 10232 19372 10284 19378
rect 10336 19360 10364 19790
rect 10284 19332 10364 19360
rect 10232 19314 10284 19320
rect 10244 19174 10272 19314
rect 10324 19236 10376 19242
rect 10324 19178 10376 19184
rect 9956 19168 10008 19174
rect 9956 19110 10008 19116
rect 10232 19168 10284 19174
rect 10232 19110 10284 19116
rect 9968 18766 9996 19110
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9935 18524 10243 18544
rect 9935 18522 9941 18524
rect 9997 18522 10021 18524
rect 10077 18522 10101 18524
rect 10157 18522 10181 18524
rect 10237 18522 10243 18524
rect 9997 18470 9999 18522
rect 10179 18470 10181 18522
rect 9935 18468 9941 18470
rect 9997 18468 10021 18470
rect 10077 18468 10101 18470
rect 10157 18468 10181 18470
rect 10237 18468 10243 18470
rect 9935 18448 10243 18468
rect 10336 18426 10364 19178
rect 10428 18465 10456 21626
rect 10414 18456 10470 18465
rect 10324 18420 10376 18426
rect 10414 18391 10470 18400
rect 10324 18362 10376 18368
rect 10140 18284 10192 18290
rect 10520 18272 10548 23122
rect 10612 22094 10640 23446
rect 10704 23254 10732 24686
rect 10796 24410 10824 24754
rect 10784 24404 10836 24410
rect 10784 24346 10836 24352
rect 10784 23724 10836 23730
rect 10784 23666 10836 23672
rect 10796 23322 10824 23666
rect 10784 23316 10836 23322
rect 10784 23258 10836 23264
rect 10692 23248 10744 23254
rect 10692 23190 10744 23196
rect 10888 23186 10916 24754
rect 10980 24274 11008 25094
rect 10968 24268 11020 24274
rect 10968 24210 11020 24216
rect 11072 23202 11100 28376
rect 11152 28358 11204 28364
rect 11164 27470 11192 28358
rect 11152 27464 11204 27470
rect 11152 27406 11204 27412
rect 11348 27130 11376 28494
rect 11980 28416 12032 28422
rect 11980 28358 12032 28364
rect 12164 28416 12216 28422
rect 12164 28358 12216 28364
rect 11336 27124 11388 27130
rect 11336 27066 11388 27072
rect 11520 26988 11572 26994
rect 11520 26930 11572 26936
rect 11428 26920 11480 26926
rect 11428 26862 11480 26868
rect 11152 26784 11204 26790
rect 11152 26726 11204 26732
rect 11164 24818 11192 26726
rect 11440 26586 11468 26862
rect 11428 26580 11480 26586
rect 11428 26522 11480 26528
rect 11440 26372 11468 26522
rect 11428 26366 11480 26372
rect 11256 26314 11428 26330
rect 11256 26308 11480 26314
rect 11256 26302 11468 26308
rect 11152 24812 11204 24818
rect 11152 24754 11204 24760
rect 11152 24200 11204 24206
rect 11152 24142 11204 24148
rect 11164 23798 11192 24142
rect 11152 23792 11204 23798
rect 11152 23734 11204 23740
rect 10876 23180 10928 23186
rect 11072 23174 11192 23202
rect 10876 23122 10928 23128
rect 11060 23112 11112 23118
rect 11060 23054 11112 23060
rect 11072 22778 11100 23054
rect 11060 22772 11112 22778
rect 11060 22714 11112 22720
rect 10876 22568 10928 22574
rect 10876 22510 10928 22516
rect 10612 22066 10824 22094
rect 10600 22024 10652 22030
rect 10600 21966 10652 21972
rect 10612 21690 10640 21966
rect 10600 21684 10652 21690
rect 10652 21644 10732 21672
rect 10600 21626 10652 21632
rect 10598 21584 10654 21593
rect 10598 21519 10600 21528
rect 10652 21519 10654 21528
rect 10600 21490 10652 21496
rect 10704 21418 10732 21644
rect 10692 21412 10744 21418
rect 10692 21354 10744 21360
rect 10692 21140 10744 21146
rect 10692 21082 10744 21088
rect 10600 20936 10652 20942
rect 10600 20878 10652 20884
rect 10612 20534 10640 20878
rect 10600 20528 10652 20534
rect 10600 20470 10652 20476
rect 10600 20392 10652 20398
rect 10704 20369 10732 21082
rect 10600 20334 10652 20340
rect 10690 20360 10746 20369
rect 10612 18873 10640 20334
rect 10690 20295 10746 20304
rect 10692 19440 10744 19446
rect 10692 19382 10744 19388
rect 10704 18902 10732 19382
rect 10796 19281 10824 22066
rect 10888 21350 10916 22510
rect 11164 22409 11192 23174
rect 11150 22400 11206 22409
rect 11150 22335 11206 22344
rect 11256 22094 11284 26302
rect 11428 26240 11480 26246
rect 11428 26182 11480 26188
rect 11336 22636 11388 22642
rect 11336 22578 11388 22584
rect 11072 22066 11284 22094
rect 10968 21956 11020 21962
rect 10968 21898 11020 21904
rect 10876 21344 10928 21350
rect 10876 21286 10928 21292
rect 10876 20936 10928 20942
rect 10874 20904 10876 20913
rect 10928 20904 10930 20913
rect 10874 20839 10930 20848
rect 10876 19780 10928 19786
rect 10876 19722 10928 19728
rect 10782 19272 10838 19281
rect 10782 19207 10838 19216
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10692 18896 10744 18902
rect 10598 18864 10654 18873
rect 10692 18838 10744 18844
rect 10598 18799 10654 18808
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 10600 18692 10652 18698
rect 10600 18634 10652 18640
rect 10140 18226 10192 18232
rect 10336 18244 10548 18272
rect 10152 18193 10180 18226
rect 10138 18184 10194 18193
rect 10048 18148 10100 18154
rect 10138 18119 10194 18128
rect 10048 18090 10100 18096
rect 10060 17921 10088 18090
rect 10140 18080 10192 18086
rect 10138 18048 10140 18057
rect 10192 18048 10194 18057
rect 10138 17983 10194 17992
rect 10046 17912 10102 17921
rect 10046 17847 10102 17856
rect 9935 17436 10243 17456
rect 9935 17434 9941 17436
rect 9997 17434 10021 17436
rect 10077 17434 10101 17436
rect 10157 17434 10181 17436
rect 10237 17434 10243 17436
rect 9997 17382 9999 17434
rect 10179 17382 10181 17434
rect 9935 17380 9941 17382
rect 9997 17380 10021 17382
rect 10077 17380 10101 17382
rect 10157 17380 10181 17382
rect 10237 17380 10243 17382
rect 9935 17360 10243 17380
rect 9935 16348 10243 16368
rect 9935 16346 9941 16348
rect 9997 16346 10021 16348
rect 10077 16346 10101 16348
rect 10157 16346 10181 16348
rect 10237 16346 10243 16348
rect 9997 16294 9999 16346
rect 10179 16294 10181 16346
rect 9935 16292 9941 16294
rect 9997 16292 10021 16294
rect 10077 16292 10101 16294
rect 10157 16292 10181 16294
rect 10237 16292 10243 16294
rect 9935 16272 10243 16292
rect 10336 15994 10364 18244
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10520 17202 10548 17478
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10140 15972 10192 15978
rect 10336 15966 10456 15994
rect 10140 15914 10192 15920
rect 10152 15706 10180 15914
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10336 15502 10364 15846
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 9935 15260 10243 15280
rect 9935 15258 9941 15260
rect 9997 15258 10021 15260
rect 10077 15258 10101 15260
rect 10157 15258 10181 15260
rect 10237 15258 10243 15260
rect 9997 15206 9999 15258
rect 10179 15206 10181 15258
rect 9935 15204 9941 15206
rect 9997 15204 10021 15206
rect 10077 15204 10101 15206
rect 10157 15204 10181 15206
rect 10237 15204 10243 15206
rect 9935 15184 10243 15204
rect 10428 14906 10456 15966
rect 10520 15638 10548 17138
rect 10612 15706 10640 18634
rect 10704 18601 10732 18702
rect 10690 18592 10746 18601
rect 10690 18527 10746 18536
rect 10796 17678 10824 19110
rect 10888 18902 10916 19722
rect 10980 19446 11008 21898
rect 10968 19440 11020 19446
rect 10968 19382 11020 19388
rect 10876 18896 10928 18902
rect 10876 18838 10928 18844
rect 10966 18864 11022 18873
rect 10966 18799 11022 18808
rect 10874 18728 10930 18737
rect 10874 18663 10876 18672
rect 10928 18663 10930 18672
rect 10876 18634 10928 18640
rect 10980 18601 11008 18799
rect 10966 18592 11022 18601
rect 10966 18527 11022 18536
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10888 18290 10916 18362
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 10888 17542 10916 18226
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10690 17232 10746 17241
rect 10690 17167 10746 17176
rect 10704 16522 10732 17167
rect 10980 17134 11008 18527
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 10968 16992 11020 16998
rect 10968 16934 11020 16940
rect 10980 16522 11008 16934
rect 10692 16516 10744 16522
rect 10692 16458 10744 16464
rect 10968 16516 11020 16522
rect 10968 16458 11020 16464
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 10508 15632 10560 15638
rect 10508 15574 10560 15580
rect 10600 15564 10652 15570
rect 10600 15506 10652 15512
rect 10612 15026 10640 15506
rect 10600 15020 10652 15026
rect 10600 14962 10652 14968
rect 9864 14884 9916 14890
rect 10428 14878 10640 14906
rect 9864 14826 9916 14832
rect 9862 14648 9918 14657
rect 9772 14612 9824 14618
rect 9862 14583 9918 14592
rect 9772 14554 9824 14560
rect 9876 14550 9904 14583
rect 9864 14544 9916 14550
rect 10612 14498 10640 14878
rect 9864 14486 9916 14492
rect 10428 14470 10640 14498
rect 10704 14482 10732 16458
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10796 15570 10824 16050
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10784 14884 10836 14890
rect 10784 14826 10836 14832
rect 10692 14476 10744 14482
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 9784 13802 9812 14350
rect 9935 14172 10243 14192
rect 9935 14170 9941 14172
rect 9997 14170 10021 14172
rect 10077 14170 10101 14172
rect 10157 14170 10181 14172
rect 10237 14170 10243 14172
rect 9997 14118 9999 14170
rect 10179 14118 10181 14170
rect 9935 14116 9941 14118
rect 9997 14116 10021 14118
rect 10077 14116 10101 14118
rect 10157 14116 10181 14118
rect 10237 14116 10243 14118
rect 9935 14096 10243 14116
rect 10336 13802 10364 14350
rect 9772 13796 9824 13802
rect 9772 13738 9824 13744
rect 10324 13796 10376 13802
rect 10324 13738 10376 13744
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9784 13190 9812 13738
rect 9956 13728 10008 13734
rect 9876 13688 9956 13716
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9784 12374 9812 12786
rect 9772 12368 9824 12374
rect 9586 12336 9642 12345
rect 9772 12310 9824 12316
rect 9586 12271 9642 12280
rect 9588 12164 9640 12170
rect 9876 12152 9904 13688
rect 9956 13670 10008 13676
rect 9935 13084 10243 13104
rect 9935 13082 9941 13084
rect 9997 13082 10021 13084
rect 10077 13082 10101 13084
rect 10157 13082 10181 13084
rect 10237 13082 10243 13084
rect 9997 13030 9999 13082
rect 10179 13030 10181 13082
rect 9935 13028 9941 13030
rect 9997 13028 10021 13030
rect 10077 13028 10101 13030
rect 10157 13028 10181 13030
rect 10237 13028 10243 13030
rect 9935 13008 10243 13028
rect 10336 12986 10364 13738
rect 10428 13734 10456 14470
rect 10692 14418 10744 14424
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 10690 14376 10746 14385
rect 10612 14278 10640 14350
rect 10690 14311 10746 14320
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10612 13802 10640 14214
rect 10704 14074 10732 14311
rect 10796 14074 10824 14826
rect 10888 14113 10916 14894
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 10874 14104 10930 14113
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10784 14068 10836 14074
rect 10874 14039 10930 14048
rect 10784 14010 10836 14016
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10704 13530 10732 13874
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10060 12442 10088 12786
rect 10414 12744 10470 12753
rect 10414 12679 10470 12688
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 9588 12106 9640 12112
rect 9784 12124 9904 12152
rect 9600 11898 9628 12106
rect 9784 12050 9812 12124
rect 9692 12022 9812 12050
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9586 11792 9642 11801
rect 9586 11727 9642 11736
rect 9416 11354 9536 11370
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9404 11348 9536 11354
rect 9456 11342 9536 11348
rect 9404 11290 9456 11296
rect 9310 11248 9366 11257
rect 9310 11183 9366 11192
rect 9048 11070 9168 11098
rect 8942 10976 8998 10985
rect 8942 10911 8998 10920
rect 8850 10840 8906 10849
rect 8850 10775 8906 10784
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8772 3670 8800 5306
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 8864 2774 8892 10775
rect 8956 8022 8984 10911
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 9048 9382 9076 9658
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9048 8838 9076 9318
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 8944 8016 8996 8022
rect 8944 7958 8996 7964
rect 8944 7812 8996 7818
rect 8944 7754 8996 7760
rect 8956 6458 8984 7754
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8942 6352 8998 6361
rect 8942 6287 8944 6296
rect 8996 6287 8998 6296
rect 8944 6258 8996 6264
rect 8864 2746 8984 2774
rect 8956 800 8984 2746
rect 9048 2038 9076 8434
rect 9140 4146 9168 11070
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 9232 10062 9260 10746
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9232 8974 9260 9998
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 9232 6934 9260 8774
rect 9220 6928 9272 6934
rect 9220 6870 9272 6876
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9232 6322 9260 6734
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9232 5370 9260 5646
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9232 4622 9260 5306
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9036 2032 9088 2038
rect 9036 1974 9088 1980
rect 9232 800 9260 3878
rect 9324 2774 9352 11183
rect 9416 9586 9444 11290
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9508 9722 9536 9862
rect 9600 9738 9628 11727
rect 9692 11082 9720 12022
rect 9935 11996 10243 12016
rect 9935 11994 9941 11996
rect 9997 11994 10021 11996
rect 10077 11994 10101 11996
rect 10157 11994 10181 11996
rect 10237 11994 10243 11996
rect 9997 11942 9999 11994
rect 10179 11942 10181 11994
rect 9935 11940 9941 11942
rect 9997 11940 10021 11942
rect 10077 11940 10101 11942
rect 10157 11940 10181 11942
rect 10237 11940 10243 11942
rect 9935 11920 10243 11940
rect 10336 11898 10364 12174
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 9770 11792 9826 11801
rect 9770 11727 9826 11736
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9692 10062 9720 11018
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9784 9874 9812 11727
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 9876 9874 9904 11222
rect 9935 10908 10243 10928
rect 9935 10906 9941 10908
rect 9997 10906 10021 10908
rect 10077 10906 10101 10908
rect 10157 10906 10181 10908
rect 10237 10906 10243 10908
rect 9997 10854 9999 10906
rect 10179 10854 10181 10906
rect 9935 10852 9941 10854
rect 9997 10852 10021 10854
rect 10077 10852 10101 10854
rect 10157 10852 10181 10854
rect 10237 10852 10243 10854
rect 9935 10832 10243 10852
rect 10140 10736 10192 10742
rect 9954 10704 10010 10713
rect 10140 10678 10192 10684
rect 9954 10639 9956 10648
rect 10008 10639 10010 10648
rect 9956 10610 10008 10616
rect 10152 10441 10180 10678
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10138 10432 10194 10441
rect 10138 10367 10194 10376
rect 10138 10160 10194 10169
rect 10138 10095 10140 10104
rect 10192 10095 10194 10104
rect 10140 10066 10192 10072
rect 10336 9897 10364 10542
rect 10428 10010 10456 12679
rect 10520 12238 10548 13330
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10612 12306 10640 12718
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10598 12200 10654 12209
rect 10598 12135 10654 12144
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10428 9982 10468 10010
rect 9753 9846 9812 9874
rect 9856 9846 9904 9874
rect 10322 9888 10378 9897
rect 9496 9716 9548 9722
rect 9600 9710 9720 9738
rect 9496 9658 9548 9664
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9416 7274 9444 8978
rect 9508 8566 9536 9522
rect 9586 8936 9642 8945
rect 9586 8871 9588 8880
rect 9640 8871 9642 8880
rect 9588 8842 9640 8848
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9496 8424 9548 8430
rect 9494 8392 9496 8401
rect 9548 8392 9550 8401
rect 9494 8327 9550 8336
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9404 7268 9456 7274
rect 9404 7210 9456 7216
rect 9508 6934 9536 7754
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9496 6928 9548 6934
rect 9496 6870 9548 6876
rect 9508 6186 9536 6870
rect 9600 6322 9628 7142
rect 9692 6458 9720 9710
rect 9753 9674 9781 9846
rect 9856 9674 9884 9846
rect 9935 9820 10243 9840
rect 10322 9823 10378 9832
rect 9935 9818 9941 9820
rect 9997 9818 10021 9820
rect 10077 9818 10101 9820
rect 10157 9818 10181 9820
rect 10237 9818 10243 9820
rect 9997 9766 9999 9818
rect 10179 9766 10181 9818
rect 9935 9764 9941 9766
rect 9997 9764 10021 9766
rect 10077 9764 10101 9766
rect 10157 9764 10181 9766
rect 10237 9764 10243 9766
rect 9935 9744 10243 9764
rect 10322 9752 10378 9761
rect 10322 9687 10378 9696
rect 9753 9646 9812 9674
rect 9856 9646 9904 9674
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9496 6180 9548 6186
rect 9496 6122 9548 6128
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9416 5778 9444 6054
rect 9404 5772 9456 5778
rect 9404 5714 9456 5720
rect 9508 5574 9536 6122
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9416 4078 9444 5510
rect 9600 4826 9628 6258
rect 9678 5672 9734 5681
rect 9678 5607 9680 5616
rect 9732 5607 9734 5616
rect 9680 5578 9732 5584
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9508 4010 9536 4558
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 9508 3534 9536 3946
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9692 3194 9720 3402
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9324 2746 9536 2774
rect 9508 800 9536 2746
rect 9784 800 9812 9646
rect 9876 9586 9904 9646
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 10230 9480 10286 9489
rect 10230 9415 10232 9424
rect 10284 9415 10286 9424
rect 10232 9386 10284 9392
rect 9956 9376 10008 9382
rect 9862 9344 9918 9353
rect 9956 9318 10008 9324
rect 9862 9279 9918 9288
rect 9876 8430 9904 9279
rect 9968 9178 9996 9318
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 9935 8732 10243 8752
rect 9935 8730 9941 8732
rect 9997 8730 10021 8732
rect 10077 8730 10101 8732
rect 10157 8730 10181 8732
rect 10237 8730 10243 8732
rect 9997 8678 9999 8730
rect 10179 8678 10181 8730
rect 9935 8676 9941 8678
rect 9997 8676 10021 8678
rect 10077 8676 10101 8678
rect 10157 8676 10181 8678
rect 10237 8676 10243 8678
rect 9935 8656 10243 8676
rect 10138 8528 10194 8537
rect 10138 8463 10194 8472
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 10046 8392 10102 8401
rect 9876 7410 9904 8366
rect 10046 8327 10102 8336
rect 10060 7886 10088 8327
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10152 7818 10180 8463
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 9935 7644 10243 7664
rect 9935 7642 9941 7644
rect 9997 7642 10021 7644
rect 10077 7642 10101 7644
rect 10157 7642 10181 7644
rect 10237 7642 10243 7644
rect 9997 7590 9999 7642
rect 10179 7590 10181 7642
rect 9935 7588 9941 7590
rect 9997 7588 10021 7590
rect 10077 7588 10101 7590
rect 10157 7588 10181 7590
rect 10237 7588 10243 7590
rect 9935 7568 10243 7588
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 9876 6440 9904 7346
rect 10244 6934 10272 7346
rect 10232 6928 10284 6934
rect 10232 6870 10284 6876
rect 9935 6556 10243 6576
rect 9935 6554 9941 6556
rect 9997 6554 10021 6556
rect 10077 6554 10101 6556
rect 10157 6554 10181 6556
rect 10237 6554 10243 6556
rect 9997 6502 9999 6554
rect 10179 6502 10181 6554
rect 9935 6500 9941 6502
rect 9997 6500 10021 6502
rect 10077 6500 10101 6502
rect 10157 6500 10181 6502
rect 10237 6500 10243 6502
rect 9935 6480 10243 6500
rect 9876 6412 9996 6440
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9876 5370 9904 6258
rect 9968 5681 9996 6412
rect 10230 6216 10286 6225
rect 10230 6151 10286 6160
rect 10244 5846 10272 6151
rect 10232 5840 10284 5846
rect 10232 5782 10284 5788
rect 9954 5672 10010 5681
rect 9954 5607 10010 5616
rect 9935 5468 10243 5488
rect 9935 5466 9941 5468
rect 9997 5466 10021 5468
rect 10077 5466 10101 5468
rect 10157 5466 10181 5468
rect 10237 5466 10243 5468
rect 9997 5414 9999 5466
rect 10179 5414 10181 5466
rect 9935 5412 9941 5414
rect 9997 5412 10021 5414
rect 10077 5412 10101 5414
rect 10157 5412 10181 5414
rect 10237 5412 10243 5414
rect 9935 5392 10243 5412
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 10230 5264 10286 5273
rect 10230 5199 10286 5208
rect 10244 4622 10272 5199
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 9876 2854 9904 4558
rect 9935 4380 10243 4400
rect 9935 4378 9941 4380
rect 9997 4378 10021 4380
rect 10077 4378 10101 4380
rect 10157 4378 10181 4380
rect 10237 4378 10243 4380
rect 9997 4326 9999 4378
rect 10179 4326 10181 4378
rect 9935 4324 9941 4326
rect 9997 4324 10021 4326
rect 10077 4324 10101 4326
rect 10157 4324 10181 4326
rect 10237 4324 10243 4326
rect 9935 4304 10243 4324
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 9968 3670 9996 4014
rect 10336 4010 10364 9687
rect 10440 9674 10468 9982
rect 10428 9646 10468 9674
rect 10428 7324 10456 9646
rect 10520 9450 10548 11086
rect 10508 9444 10560 9450
rect 10508 9386 10560 9392
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10520 8634 10548 8910
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10520 7426 10548 7822
rect 10612 7546 10640 12135
rect 10704 11354 10732 13466
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10980 13138 11008 14418
rect 11072 13462 11100 22066
rect 11242 21992 11298 22001
rect 11242 21927 11298 21936
rect 11256 20788 11284 21927
rect 11348 21690 11376 22578
rect 11336 21684 11388 21690
rect 11336 21626 11388 21632
rect 11336 21344 11388 21350
rect 11336 21286 11388 21292
rect 11348 20942 11376 21286
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 11256 20760 11376 20788
rect 11244 20528 11296 20534
rect 11244 20470 11296 20476
rect 11152 20324 11204 20330
rect 11152 20266 11204 20272
rect 11164 18086 11192 20266
rect 11256 18737 11284 20470
rect 11242 18728 11298 18737
rect 11242 18663 11298 18672
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 11242 18048 11298 18057
rect 11242 17983 11298 17992
rect 11256 15570 11284 17983
rect 11348 17513 11376 20760
rect 11334 17504 11390 17513
rect 11334 17439 11390 17448
rect 11336 17264 11388 17270
rect 11336 17206 11388 17212
rect 11348 16289 11376 17206
rect 11334 16280 11390 16289
rect 11334 16215 11390 16224
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11152 15496 11204 15502
rect 11440 15450 11468 26182
rect 11532 26042 11560 26930
rect 11520 26036 11572 26042
rect 11520 25978 11572 25984
rect 11796 25288 11848 25294
rect 11796 25230 11848 25236
rect 11520 24608 11572 24614
rect 11520 24550 11572 24556
rect 11532 23526 11560 24550
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 11612 24132 11664 24138
rect 11612 24074 11664 24080
rect 11624 23866 11652 24074
rect 11612 23860 11664 23866
rect 11612 23802 11664 23808
rect 11716 23662 11744 24142
rect 11704 23656 11756 23662
rect 11704 23598 11756 23604
rect 11808 23644 11836 25230
rect 11888 23656 11940 23662
rect 11808 23616 11888 23644
rect 11520 23520 11572 23526
rect 11520 23462 11572 23468
rect 11532 23118 11560 23462
rect 11520 23112 11572 23118
rect 11520 23054 11572 23060
rect 11704 23112 11756 23118
rect 11704 23054 11756 23060
rect 11612 22092 11664 22098
rect 11612 22034 11664 22040
rect 11520 21480 11572 21486
rect 11520 21422 11572 21428
rect 11532 21350 11560 21422
rect 11520 21344 11572 21350
rect 11520 21286 11572 21292
rect 11520 20800 11572 20806
rect 11520 20742 11572 20748
rect 11532 20058 11560 20742
rect 11520 20052 11572 20058
rect 11520 19994 11572 20000
rect 11624 19378 11652 22034
rect 11612 19372 11664 19378
rect 11612 19314 11664 19320
rect 11520 19168 11572 19174
rect 11520 19110 11572 19116
rect 11532 17882 11560 19110
rect 11610 18864 11666 18873
rect 11610 18799 11612 18808
rect 11664 18799 11666 18808
rect 11612 18770 11664 18776
rect 11612 18692 11664 18698
rect 11612 18634 11664 18640
rect 11520 17876 11572 17882
rect 11520 17818 11572 17824
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11152 15438 11204 15444
rect 11164 14550 11192 15438
rect 11256 15422 11468 15450
rect 11152 14544 11204 14550
rect 11152 14486 11204 14492
rect 11164 13870 11192 14486
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 10796 12918 10824 13126
rect 10980 13110 11100 13138
rect 10784 12912 10836 12918
rect 10784 12854 10836 12860
rect 10968 12912 11020 12918
rect 10968 12854 11020 12860
rect 10874 12336 10930 12345
rect 10874 12271 10930 12280
rect 10782 12200 10838 12209
rect 10782 12135 10838 12144
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10704 10674 10732 11018
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10690 10568 10746 10577
rect 10690 10503 10746 10512
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10520 7398 10640 7426
rect 10428 7296 10548 7324
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10428 6322 10456 6802
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 10428 5778 10456 6258
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10520 5234 10548 7296
rect 10612 6662 10640 7398
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10612 5114 10640 6598
rect 10428 5086 10640 5114
rect 10324 4004 10376 4010
rect 10324 3946 10376 3952
rect 10428 3942 10456 5086
rect 10600 4752 10652 4758
rect 10600 4694 10652 4700
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 9956 3664 10008 3670
rect 10520 3618 10548 4218
rect 9956 3606 10008 3612
rect 10336 3590 10548 3618
rect 9935 3292 10243 3312
rect 9935 3290 9941 3292
rect 9997 3290 10021 3292
rect 10077 3290 10101 3292
rect 10157 3290 10181 3292
rect 10237 3290 10243 3292
rect 9997 3238 9999 3290
rect 10179 3238 10181 3290
rect 9935 3236 9941 3238
rect 9997 3236 10021 3238
rect 10077 3236 10101 3238
rect 10157 3236 10181 3238
rect 10237 3236 10243 3238
rect 9935 3216 10243 3236
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 9876 2446 9904 2790
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 9935 2204 10243 2224
rect 9935 2202 9941 2204
rect 9997 2202 10021 2204
rect 10077 2202 10101 2204
rect 10157 2202 10181 2204
rect 10237 2202 10243 2204
rect 9997 2150 9999 2202
rect 10179 2150 10181 2202
rect 9935 2148 9941 2150
rect 9997 2148 10021 2150
rect 10077 2148 10101 2150
rect 10157 2148 10181 2150
rect 10237 2148 10243 2150
rect 9935 2128 10243 2148
rect 10336 2088 10364 3590
rect 10612 3534 10640 4694
rect 10704 4214 10732 10503
rect 10796 5352 10824 12135
rect 10888 5930 10916 12271
rect 10980 11218 11008 12854
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 10968 11008 11020 11014
rect 10968 10950 11020 10956
rect 10980 10849 11008 10950
rect 10966 10840 11022 10849
rect 10966 10775 11022 10784
rect 11072 10554 11100 13110
rect 11164 12986 11192 13670
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11164 10674 11192 12922
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 11072 10526 11192 10554
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10980 9926 11008 9998
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 10980 6118 11008 9590
rect 11072 9586 11100 10406
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11164 9382 11192 10526
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11072 8673 11100 8910
rect 11058 8664 11114 8673
rect 11058 8599 11114 8608
rect 11164 8498 11192 9318
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11072 7886 11100 8434
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 11072 7002 11100 7686
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 11150 6896 11206 6905
rect 11150 6831 11206 6840
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10888 5902 11008 5930
rect 10796 5324 10916 5352
rect 10782 5264 10838 5273
rect 10782 5199 10838 5208
rect 10796 4554 10824 5199
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10888 4282 10916 5324
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 10692 4004 10744 4010
rect 10692 3946 10744 3952
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 10416 2916 10468 2922
rect 10416 2858 10468 2864
rect 10060 2060 10364 2088
rect 10060 800 10088 2060
rect 10428 1034 10456 2858
rect 10520 2582 10548 3062
rect 10612 3058 10640 3470
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10508 2576 10560 2582
rect 10508 2518 10560 2524
rect 10612 2446 10640 2994
rect 10704 2990 10732 3946
rect 10692 2984 10744 2990
rect 10692 2926 10744 2932
rect 10796 2774 10824 4082
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10888 3466 10916 4014
rect 10980 3942 11008 5902
rect 11072 5370 11100 6326
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11058 5128 11114 5137
rect 11058 5063 11114 5072
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10876 3460 10928 3466
rect 10876 3402 10928 3408
rect 10888 3194 10916 3402
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10980 3040 11008 3674
rect 10704 2746 10824 2774
rect 10888 3012 11008 3040
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10704 1442 10732 2746
rect 10336 1006 10456 1034
rect 10612 1414 10732 1442
rect 10336 800 10364 1006
rect 10612 800 10640 1414
rect 10888 800 10916 3012
rect 11072 2904 11100 5063
rect 10980 2876 11100 2904
rect 10980 2650 11008 2876
rect 11058 2816 11114 2825
rect 11058 2751 11114 2760
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 10966 2544 11022 2553
rect 10966 2479 11022 2488
rect 10980 2378 11008 2479
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 11072 2310 11100 2751
rect 11164 2666 11192 6831
rect 11256 4010 11284 15422
rect 11336 15020 11388 15026
rect 11336 14962 11388 14968
rect 11348 14929 11376 14962
rect 11428 14952 11480 14958
rect 11334 14920 11390 14929
rect 11428 14894 11480 14900
rect 11334 14855 11390 14864
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11348 14346 11376 14758
rect 11336 14340 11388 14346
rect 11336 14282 11388 14288
rect 11348 13394 11376 14282
rect 11440 13938 11468 14894
rect 11532 14414 11560 17478
rect 11624 16794 11652 18634
rect 11716 18222 11744 23054
rect 11808 21894 11836 23616
rect 11888 23598 11940 23604
rect 11888 22704 11940 22710
rect 11888 22646 11940 22652
rect 11900 22098 11928 22646
rect 11888 22092 11940 22098
rect 11888 22034 11940 22040
rect 11796 21888 11848 21894
rect 11796 21830 11848 21836
rect 11808 20942 11836 21830
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 11888 20868 11940 20874
rect 11888 20810 11940 20816
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11808 18290 11836 20402
rect 11900 20398 11928 20810
rect 11888 20392 11940 20398
rect 11888 20334 11940 20340
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11900 19174 11928 19314
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11808 17542 11836 18022
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11796 17264 11848 17270
rect 11796 17206 11848 17212
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11612 16108 11664 16114
rect 11716 16096 11744 17138
rect 11664 16068 11744 16096
rect 11612 16050 11664 16056
rect 11520 14408 11572 14414
rect 11520 14350 11572 14356
rect 11518 14240 11574 14249
rect 11518 14175 11574 14184
rect 11532 14074 11560 14175
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11518 13968 11574 13977
rect 11428 13932 11480 13938
rect 11518 13903 11520 13912
rect 11428 13874 11480 13880
rect 11572 13903 11574 13912
rect 11520 13874 11572 13880
rect 11624 13870 11652 16050
rect 11808 15688 11836 17206
rect 11716 15660 11836 15688
rect 11716 14958 11744 15660
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11716 14618 11744 14758
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11808 14226 11836 15506
rect 11900 15314 11928 18906
rect 11992 17105 12020 28358
rect 12176 27713 12204 28358
rect 12820 28218 12848 28698
rect 13544 28688 13596 28694
rect 13544 28630 13596 28636
rect 13176 28552 13228 28558
rect 13176 28494 13228 28500
rect 13084 28416 13136 28422
rect 13084 28358 13136 28364
rect 12808 28212 12860 28218
rect 12808 28154 12860 28160
rect 12532 28076 12584 28082
rect 12532 28018 12584 28024
rect 12162 27704 12218 27713
rect 12162 27639 12218 27648
rect 12440 27328 12492 27334
rect 12440 27270 12492 27276
rect 12072 26784 12124 26790
rect 12072 26726 12124 26732
rect 12084 24818 12112 26726
rect 12256 26376 12308 26382
rect 12256 26318 12308 26324
rect 12268 25702 12296 26318
rect 12452 26042 12480 27270
rect 12544 27130 12572 28018
rect 13096 27674 13124 28358
rect 13188 27878 13216 28494
rect 13556 27878 13584 28630
rect 14004 28620 14056 28626
rect 14004 28562 14056 28568
rect 13728 28552 13780 28558
rect 13728 28494 13780 28500
rect 13176 27872 13228 27878
rect 13176 27814 13228 27820
rect 13544 27872 13596 27878
rect 13544 27814 13596 27820
rect 13084 27668 13136 27674
rect 13084 27610 13136 27616
rect 13188 27554 13216 27814
rect 13096 27526 13216 27554
rect 12716 27328 12768 27334
rect 12716 27270 12768 27276
rect 12532 27124 12584 27130
rect 12532 27066 12584 27072
rect 12728 26994 12756 27270
rect 12900 27056 12952 27062
rect 12900 26998 12952 27004
rect 12716 26988 12768 26994
rect 12716 26930 12768 26936
rect 12912 26450 12940 26998
rect 12532 26444 12584 26450
rect 12532 26386 12584 26392
rect 12900 26444 12952 26450
rect 12900 26386 12952 26392
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 12440 25900 12492 25906
rect 12440 25842 12492 25848
rect 12256 25696 12308 25702
rect 12256 25638 12308 25644
rect 12072 24812 12124 24818
rect 12072 24754 12124 24760
rect 12268 24682 12296 25638
rect 12452 25498 12480 25842
rect 12440 25492 12492 25498
rect 12440 25434 12492 25440
rect 12440 25356 12492 25362
rect 12440 25298 12492 25304
rect 12452 24954 12480 25298
rect 12440 24948 12492 24954
rect 12440 24890 12492 24896
rect 12348 24812 12400 24818
rect 12348 24754 12400 24760
rect 12072 24676 12124 24682
rect 12072 24618 12124 24624
rect 12256 24676 12308 24682
rect 12256 24618 12308 24624
rect 12084 23100 12112 24618
rect 12360 24614 12388 24754
rect 12348 24608 12400 24614
rect 12348 24550 12400 24556
rect 12544 24410 12572 26386
rect 12808 26036 12860 26042
rect 12808 25978 12860 25984
rect 12624 25968 12676 25974
rect 12624 25910 12676 25916
rect 12636 24886 12664 25910
rect 12820 25362 12848 25978
rect 12992 25900 13044 25906
rect 12992 25842 13044 25848
rect 13004 25498 13032 25842
rect 13096 25498 13124 27526
rect 13556 27470 13584 27814
rect 13544 27464 13596 27470
rect 13544 27406 13596 27412
rect 13634 27432 13690 27441
rect 13634 27367 13690 27376
rect 13176 26920 13228 26926
rect 13176 26862 13228 26868
rect 12992 25492 13044 25498
rect 12992 25434 13044 25440
rect 13084 25492 13136 25498
rect 13084 25434 13136 25440
rect 12808 25356 12860 25362
rect 12808 25298 12860 25304
rect 12624 24880 12676 24886
rect 12624 24822 12676 24828
rect 12820 24750 12848 25298
rect 12900 25288 12952 25294
rect 12900 25230 12952 25236
rect 12624 24744 12676 24750
rect 12624 24686 12676 24692
rect 12808 24744 12860 24750
rect 12808 24686 12860 24692
rect 12532 24404 12584 24410
rect 12452 24364 12532 24392
rect 12256 23112 12308 23118
rect 12084 23072 12256 23100
rect 12452 23100 12480 24364
rect 12532 24346 12584 24352
rect 12636 24138 12664 24686
rect 12912 24614 12940 25230
rect 13096 24954 13124 25434
rect 13084 24948 13136 24954
rect 13084 24890 13136 24896
rect 13188 24682 13216 26862
rect 13268 26852 13320 26858
rect 13268 26794 13320 26800
rect 13280 26489 13308 26794
rect 13266 26480 13322 26489
rect 13266 26415 13322 26424
rect 13360 26308 13412 26314
rect 13360 26250 13412 26256
rect 13268 25900 13320 25906
rect 13268 25842 13320 25848
rect 13280 25294 13308 25842
rect 13268 25288 13320 25294
rect 13268 25230 13320 25236
rect 13176 24676 13228 24682
rect 13176 24618 13228 24624
rect 12900 24608 12952 24614
rect 12900 24550 12952 24556
rect 13176 24200 13228 24206
rect 13176 24142 13228 24148
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 12532 23724 12584 23730
rect 12532 23666 12584 23672
rect 12544 23322 12572 23666
rect 12532 23316 12584 23322
rect 12532 23258 12584 23264
rect 12532 23112 12584 23118
rect 12452 23072 12532 23100
rect 12256 23054 12308 23060
rect 12532 23054 12584 23060
rect 12072 22636 12124 22642
rect 12072 22578 12124 22584
rect 12084 22030 12112 22578
rect 12164 22568 12216 22574
rect 12164 22510 12216 22516
rect 12176 22166 12204 22510
rect 12164 22160 12216 22166
rect 12164 22102 12216 22108
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 12176 21690 12204 22102
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 12268 21570 12296 23054
rect 12348 22976 12400 22982
rect 12348 22918 12400 22924
rect 12360 21622 12388 22918
rect 12544 22642 12572 23054
rect 12624 23044 12676 23050
rect 12624 22986 12676 22992
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12440 22568 12492 22574
rect 12440 22510 12492 22516
rect 12452 21894 12480 22510
rect 12636 22386 12664 22986
rect 12900 22772 12952 22778
rect 12900 22714 12952 22720
rect 12636 22358 12756 22386
rect 12532 21956 12584 21962
rect 12532 21898 12584 21904
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 12176 21542 12296 21570
rect 12348 21616 12400 21622
rect 12348 21558 12400 21564
rect 12176 21434 12204 21542
rect 12084 21406 12204 21434
rect 12256 21480 12308 21486
rect 12256 21422 12308 21428
rect 12084 20262 12112 21406
rect 12164 20800 12216 20806
rect 12164 20742 12216 20748
rect 12072 20256 12124 20262
rect 12072 20198 12124 20204
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 12084 19378 12112 19790
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 12176 18766 12204 20742
rect 12268 19718 12296 21422
rect 12348 20460 12400 20466
rect 12400 20420 12480 20448
rect 12348 20402 12400 20408
rect 12346 20360 12402 20369
rect 12346 20295 12402 20304
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12268 18902 12296 19654
rect 12256 18896 12308 18902
rect 12256 18838 12308 18844
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12084 18358 12112 18702
rect 12072 18352 12124 18358
rect 12072 18294 12124 18300
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 11978 17096 12034 17105
rect 11978 17031 12034 17040
rect 11900 15286 12020 15314
rect 11886 14648 11942 14657
rect 11886 14583 11942 14592
rect 11900 14346 11928 14583
rect 11888 14340 11940 14346
rect 11888 14282 11940 14288
rect 11808 14198 11928 14226
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11520 13456 11572 13462
rect 11520 13398 11572 13404
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 11348 10713 11376 13330
rect 11532 12850 11560 13398
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11428 11348 11480 11354
rect 11428 11290 11480 11296
rect 11440 11150 11468 11290
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11426 10976 11482 10985
rect 11426 10911 11482 10920
rect 11334 10704 11390 10713
rect 11334 10639 11390 10648
rect 11348 10062 11376 10639
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 11348 5710 11376 7754
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11440 5352 11468 10911
rect 11532 9489 11560 12786
rect 11624 12170 11652 13806
rect 11716 12306 11744 13806
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11716 11558 11744 12242
rect 11900 12102 11928 14198
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11992 11898 12020 15286
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11716 10606 11744 11494
rect 11900 11150 11928 11494
rect 11888 11144 11940 11150
rect 11808 11104 11888 11132
rect 11808 10810 11836 11104
rect 11888 11086 11940 11092
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11716 10169 11744 10542
rect 11808 10266 11836 10746
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 11702 10160 11758 10169
rect 11702 10095 11758 10104
rect 11518 9480 11574 9489
rect 11518 9415 11574 9424
rect 11716 8974 11744 10095
rect 11900 9926 11928 10406
rect 11992 10266 12020 10610
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 11888 9716 11940 9722
rect 11888 9658 11940 9664
rect 11796 9648 11848 9654
rect 11796 9590 11848 9596
rect 11808 9353 11836 9590
rect 11794 9344 11850 9353
rect 11794 9279 11850 9288
rect 11900 8974 11928 9658
rect 11704 8968 11756 8974
rect 11888 8968 11940 8974
rect 11704 8910 11756 8916
rect 11794 8936 11850 8945
rect 11888 8910 11940 8916
rect 11794 8871 11850 8880
rect 11612 8560 11664 8566
rect 11664 8520 11744 8548
rect 11612 8502 11664 8508
rect 11610 8392 11666 8401
rect 11610 8327 11666 8336
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11532 6390 11560 7278
rect 11520 6384 11572 6390
rect 11520 6326 11572 6332
rect 11532 6254 11560 6326
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11348 5324 11468 5352
rect 11244 4004 11296 4010
rect 11244 3946 11296 3952
rect 11348 3618 11376 5324
rect 11428 5228 11480 5234
rect 11428 5170 11480 5176
rect 11440 3738 11468 5170
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11532 4826 11560 5102
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11532 4146 11560 4762
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11256 3590 11376 3618
rect 11256 2922 11284 3590
rect 11440 3534 11468 3674
rect 11624 3602 11652 8327
rect 11716 8294 11744 8520
rect 11808 8498 11836 8871
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 11716 7954 11744 8230
rect 12084 8022 12112 18158
rect 12176 17338 12204 18702
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12162 17232 12218 17241
rect 12162 17167 12164 17176
rect 12216 17167 12218 17176
rect 12164 17138 12216 17144
rect 12164 17060 12216 17066
rect 12164 17002 12216 17008
rect 12176 16522 12204 17002
rect 12164 16516 12216 16522
rect 12164 16458 12216 16464
rect 12176 16114 12204 16458
rect 12268 16250 12296 18838
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 12164 16108 12216 16114
rect 12164 16050 12216 16056
rect 12360 15994 12388 20295
rect 12452 19310 12480 20420
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 12544 19242 12572 21898
rect 12624 21888 12676 21894
rect 12624 21830 12676 21836
rect 12636 20330 12664 21830
rect 12624 20324 12676 20330
rect 12624 20266 12676 20272
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12532 19236 12584 19242
rect 12532 19178 12584 19184
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12452 17354 12480 19110
rect 12544 19009 12572 19178
rect 12530 19000 12586 19009
rect 12530 18935 12586 18944
rect 12544 18766 12572 18935
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12636 18630 12664 19314
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12624 18148 12676 18154
rect 12624 18090 12676 18096
rect 12532 18080 12584 18086
rect 12532 18022 12584 18028
rect 12544 17610 12572 18022
rect 12532 17604 12584 17610
rect 12532 17546 12584 17552
rect 12636 17513 12664 18090
rect 12622 17504 12678 17513
rect 12622 17439 12678 17448
rect 12452 17326 12664 17354
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12176 15966 12388 15994
rect 12176 14890 12204 15966
rect 12254 15872 12310 15881
rect 12254 15807 12310 15816
rect 12164 14884 12216 14890
rect 12164 14826 12216 14832
rect 12162 14784 12218 14793
rect 12162 14719 12218 14728
rect 12176 14482 12204 14719
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12268 12850 12296 15807
rect 12348 15632 12400 15638
rect 12348 15574 12400 15580
rect 12360 15094 12388 15574
rect 12348 15088 12400 15094
rect 12348 15030 12400 15036
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12360 13734 12388 14554
rect 12348 13728 12400 13734
rect 12348 13670 12400 13676
rect 12360 13326 12388 13670
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 12176 11558 12204 12718
rect 12164 11552 12216 11558
rect 12164 11494 12216 11500
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12176 10130 12204 11290
rect 12268 11014 12296 12786
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 12360 10810 12388 12582
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12360 10033 12388 10610
rect 12346 10024 12402 10033
rect 12256 9988 12308 9994
rect 12346 9959 12402 9968
rect 12256 9930 12308 9936
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12176 8838 12204 9454
rect 12268 9450 12296 9930
rect 12256 9444 12308 9450
rect 12256 9386 12308 9392
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12360 9081 12388 9114
rect 12346 9072 12402 9081
rect 12346 9007 12402 9016
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12348 8424 12400 8430
rect 12346 8392 12348 8401
rect 12400 8392 12402 8401
rect 12346 8327 12402 8336
rect 11888 8016 11940 8022
rect 11888 7958 11940 7964
rect 12072 8016 12124 8022
rect 12124 7976 12296 8004
rect 12072 7958 12124 7964
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11702 6760 11758 6769
rect 11702 6695 11704 6704
rect 11756 6695 11758 6704
rect 11704 6666 11756 6672
rect 11808 6662 11836 7346
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11716 4842 11744 6054
rect 11808 5030 11836 6598
rect 11900 6066 11928 7958
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11992 6186 12020 7822
rect 11980 6180 12032 6186
rect 11980 6122 12032 6128
rect 12164 6112 12216 6118
rect 11900 6038 12112 6066
rect 12164 6054 12216 6060
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11900 5302 11928 5510
rect 11888 5296 11940 5302
rect 11888 5238 11940 5244
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11716 4814 11836 4842
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11716 4282 11744 4558
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 11704 4004 11756 4010
rect 11704 3946 11756 3952
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 11244 2916 11296 2922
rect 11244 2858 11296 2864
rect 11164 2638 11284 2666
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11164 800 11192 2518
rect 11256 1442 11284 2638
rect 11348 2582 11376 3470
rect 11336 2576 11388 2582
rect 11336 2518 11388 2524
rect 11256 1414 11468 1442
rect 11440 800 11468 1414
rect 11716 800 11744 3946
rect 11808 2650 11836 4814
rect 11888 4752 11940 4758
rect 11888 4694 11940 4700
rect 11900 4128 11928 4694
rect 11992 4690 12020 4966
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11980 4140 12032 4146
rect 11900 4100 11980 4128
rect 11900 3534 11928 4100
rect 11980 4082 12032 4088
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11980 3460 12032 3466
rect 11980 3402 12032 3408
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 11796 2644 11848 2650
rect 11796 2586 11848 2592
rect 11900 2446 11928 3334
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11900 1970 11928 2246
rect 11888 1964 11940 1970
rect 11888 1906 11940 1912
rect 11992 800 12020 3402
rect 12084 3058 12112 6038
rect 12072 3052 12124 3058
rect 12072 2994 12124 3000
rect 12176 2825 12204 6054
rect 12268 5234 12296 7976
rect 12348 7812 12400 7818
rect 12348 7754 12400 7760
rect 12360 7342 12388 7754
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12348 6792 12400 6798
rect 12452 6780 12480 16390
rect 12544 16153 12572 16934
rect 12530 16144 12586 16153
rect 12530 16079 12586 16088
rect 12636 15745 12664 17326
rect 12622 15736 12678 15745
rect 12622 15671 12678 15680
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12636 15026 12664 15506
rect 12728 15416 12756 22358
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 12820 20505 12848 21966
rect 12912 20602 12940 22714
rect 12992 22568 13044 22574
rect 12992 22510 13044 22516
rect 13004 22234 13032 22510
rect 12992 22228 13044 22234
rect 12992 22170 13044 22176
rect 13084 21888 13136 21894
rect 13084 21830 13136 21836
rect 13096 21049 13124 21830
rect 13082 21040 13138 21049
rect 13082 20975 13138 20984
rect 13084 20936 13136 20942
rect 13084 20878 13136 20884
rect 12900 20596 12952 20602
rect 12900 20538 12952 20544
rect 13096 20534 13124 20878
rect 13084 20528 13136 20534
rect 12806 20496 12862 20505
rect 13084 20470 13136 20476
rect 12806 20431 12862 20440
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 12820 19922 12848 20334
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12990 19680 13046 19689
rect 12808 19372 12860 19378
rect 12808 19314 12860 19320
rect 12820 18465 12848 19314
rect 12806 18456 12862 18465
rect 12806 18391 12862 18400
rect 12820 17320 12848 18391
rect 12912 18290 12940 19654
rect 12990 19615 13046 19624
rect 13004 19446 13032 19615
rect 12992 19440 13044 19446
rect 12992 19382 13044 19388
rect 13096 19174 13124 20470
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 12992 18692 13044 18698
rect 12992 18634 13044 18640
rect 13004 18601 13032 18634
rect 12990 18592 13046 18601
rect 12990 18527 13046 18536
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 12820 17292 12940 17320
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 12820 16794 12848 17138
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12820 15570 12848 16730
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12728 15388 12848 15416
rect 12714 15328 12770 15337
rect 12714 15263 12770 15272
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12636 14346 12664 14962
rect 12728 14521 12756 15263
rect 12714 14512 12770 14521
rect 12714 14447 12770 14456
rect 12624 14340 12676 14346
rect 12624 14282 12676 14288
rect 12636 14074 12664 14282
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12544 11558 12572 12038
rect 12728 11914 12756 14010
rect 12820 12730 12848 15388
rect 12912 14074 12940 17292
rect 13004 14464 13032 18527
rect 13096 18329 13124 18770
rect 13082 18320 13138 18329
rect 13082 18255 13138 18264
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 13096 17202 13124 18158
rect 13188 17882 13216 24142
rect 13268 24064 13320 24070
rect 13268 24006 13320 24012
rect 13280 19854 13308 24006
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13280 18873 13308 19450
rect 13372 19394 13400 26250
rect 13648 25888 13676 27367
rect 13740 27316 13768 28494
rect 13820 28416 13872 28422
rect 13820 28358 13872 28364
rect 13832 27470 13860 28358
rect 13912 28008 13964 28014
rect 13912 27950 13964 27956
rect 13924 27606 13952 27950
rect 13912 27600 13964 27606
rect 13912 27542 13964 27548
rect 14016 27538 14044 28562
rect 15016 28552 15068 28558
rect 15016 28494 15068 28500
rect 14832 28416 14884 28422
rect 14832 28358 14884 28364
rect 14844 27985 14872 28358
rect 14830 27976 14886 27985
rect 14830 27911 14886 27920
rect 14428 27772 14736 27792
rect 14428 27770 14434 27772
rect 14490 27770 14514 27772
rect 14570 27770 14594 27772
rect 14650 27770 14674 27772
rect 14730 27770 14736 27772
rect 14490 27718 14492 27770
rect 14672 27718 14674 27770
rect 14428 27716 14434 27718
rect 14490 27716 14514 27718
rect 14570 27716 14594 27718
rect 14650 27716 14674 27718
rect 14730 27716 14736 27718
rect 14428 27696 14736 27716
rect 14004 27532 14056 27538
rect 14004 27474 14056 27480
rect 13820 27464 13872 27470
rect 13912 27464 13964 27470
rect 13820 27406 13872 27412
rect 13910 27432 13912 27441
rect 13964 27432 13966 27441
rect 13910 27367 13966 27376
rect 13740 27288 13952 27316
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 13832 26042 13860 26930
rect 13820 26036 13872 26042
rect 13820 25978 13872 25984
rect 13924 25906 13952 27288
rect 14016 26994 14044 27474
rect 14096 27396 14148 27402
rect 14096 27338 14148 27344
rect 14004 26988 14056 26994
rect 14004 26930 14056 26936
rect 14016 26518 14044 26930
rect 14004 26512 14056 26518
rect 14004 26454 14056 26460
rect 14108 26382 14136 27338
rect 14924 27328 14976 27334
rect 14924 27270 14976 27276
rect 14740 26988 14792 26994
rect 14740 26930 14792 26936
rect 14752 26874 14780 26930
rect 14752 26846 14872 26874
rect 14280 26784 14332 26790
rect 14280 26726 14332 26732
rect 14292 26586 14320 26726
rect 14428 26684 14736 26704
rect 14428 26682 14434 26684
rect 14490 26682 14514 26684
rect 14570 26682 14594 26684
rect 14650 26682 14674 26684
rect 14730 26682 14736 26684
rect 14490 26630 14492 26682
rect 14672 26630 14674 26682
rect 14428 26628 14434 26630
rect 14490 26628 14514 26630
rect 14570 26628 14594 26630
rect 14650 26628 14674 26630
rect 14730 26628 14736 26630
rect 14428 26608 14736 26628
rect 14844 26586 14872 26846
rect 14280 26580 14332 26586
rect 14280 26522 14332 26528
rect 14832 26580 14884 26586
rect 14832 26522 14884 26528
rect 14554 26480 14610 26489
rect 14554 26415 14610 26424
rect 14568 26382 14596 26415
rect 14096 26376 14148 26382
rect 14096 26318 14148 26324
rect 14556 26376 14608 26382
rect 14556 26318 14608 26324
rect 14004 26240 14056 26246
rect 14004 26182 14056 26188
rect 13912 25900 13964 25906
rect 13648 25860 13860 25888
rect 13728 25764 13780 25770
rect 13728 25706 13780 25712
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 13556 23730 13584 24754
rect 13636 24608 13688 24614
rect 13636 24550 13688 24556
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 13556 23118 13584 23666
rect 13544 23112 13596 23118
rect 13544 23054 13596 23060
rect 13544 22976 13596 22982
rect 13544 22918 13596 22924
rect 13556 22710 13584 22918
rect 13544 22704 13596 22710
rect 13544 22646 13596 22652
rect 13648 22556 13676 24550
rect 13740 23866 13768 25706
rect 13728 23860 13780 23866
rect 13728 23802 13780 23808
rect 13728 23520 13780 23526
rect 13728 23462 13780 23468
rect 13740 23322 13768 23462
rect 13728 23316 13780 23322
rect 13728 23258 13780 23264
rect 13556 22528 13676 22556
rect 13452 21684 13504 21690
rect 13556 21672 13584 22528
rect 13634 22400 13690 22409
rect 13634 22335 13690 22344
rect 13504 21644 13584 21672
rect 13452 21626 13504 21632
rect 13464 20058 13492 21626
rect 13544 20800 13596 20806
rect 13544 20742 13596 20748
rect 13556 20330 13584 20742
rect 13544 20324 13596 20330
rect 13544 20266 13596 20272
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 13450 19544 13506 19553
rect 13450 19479 13452 19488
rect 13504 19479 13506 19488
rect 13452 19450 13504 19456
rect 13372 19366 13492 19394
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13266 18864 13322 18873
rect 13266 18799 13322 18808
rect 13268 18420 13320 18426
rect 13268 18362 13320 18368
rect 13280 18086 13308 18362
rect 13268 18080 13320 18086
rect 13268 18022 13320 18028
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 13268 17876 13320 17882
rect 13268 17818 13320 17824
rect 13188 17338 13216 17818
rect 13176 17332 13228 17338
rect 13176 17274 13228 17280
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 13082 16416 13138 16425
rect 13082 16351 13138 16360
rect 13096 16114 13124 16351
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 13188 16046 13216 17274
rect 13280 17134 13308 17818
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 13082 15600 13138 15609
rect 13082 15535 13138 15544
rect 13096 15026 13124 15535
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 13280 14958 13308 17070
rect 13372 16590 13400 19110
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13358 16144 13414 16153
rect 13358 16079 13414 16088
rect 13372 15706 13400 16079
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 13372 15094 13400 15642
rect 13360 15088 13412 15094
rect 13360 15030 13412 15036
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13096 14618 13124 14758
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 13004 14436 13400 14464
rect 13176 14340 13228 14346
rect 13176 14282 13228 14288
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 13188 13977 13216 14282
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13174 13968 13230 13977
rect 13174 13903 13230 13912
rect 12820 12702 12940 12730
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 12820 12102 12848 12582
rect 12912 12102 12940 12702
rect 13082 12472 13138 12481
rect 12992 12436 13044 12442
rect 13082 12407 13138 12416
rect 12992 12378 13044 12384
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12728 11886 12940 11914
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12544 10985 12572 11494
rect 12728 11150 12756 11698
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12530 10976 12586 10985
rect 12530 10911 12586 10920
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12544 9926 12572 10610
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12544 9178 12572 9386
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12530 9072 12586 9081
rect 12530 9007 12532 9016
rect 12584 9007 12586 9016
rect 12532 8978 12584 8984
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12544 8498 12572 8774
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12544 7546 12572 8298
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12636 7478 12664 11018
rect 12728 10198 12756 11086
rect 12716 10192 12768 10198
rect 12716 10134 12768 10140
rect 12820 9042 12848 11494
rect 12912 9466 12940 11886
rect 13004 11762 13032 12378
rect 13096 11762 13124 12407
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 13096 11257 13124 11562
rect 13082 11248 13138 11257
rect 13082 11183 13138 11192
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 13096 10441 13124 10474
rect 13082 10432 13138 10441
rect 13082 10367 13138 10376
rect 13096 9994 13124 10367
rect 13084 9988 13136 9994
rect 13084 9930 13136 9936
rect 13188 9602 13216 13903
rect 13280 13433 13308 14214
rect 13266 13424 13322 13433
rect 13266 13359 13322 13368
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 13280 12442 13308 12786
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13096 9574 13216 9602
rect 12912 9438 13032 9466
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12912 8974 12940 9318
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12716 8560 12768 8566
rect 12716 8502 12768 8508
rect 12728 8362 12756 8502
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12624 7472 12676 7478
rect 12624 7414 12676 7420
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12400 6752 12480 6780
rect 12348 6734 12400 6740
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12452 5302 12480 6598
rect 12544 6390 12572 7142
rect 12728 7002 12756 7754
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 13004 6934 13032 9438
rect 12992 6928 13044 6934
rect 12636 6876 12992 6882
rect 12636 6870 13044 6876
rect 12636 6854 13032 6870
rect 12636 6798 12664 6854
rect 13004 6805 13032 6854
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 12532 6384 12584 6390
rect 12532 6326 12584 6332
rect 12440 5296 12492 5302
rect 12440 5238 12492 5244
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12544 4554 12572 6326
rect 12728 6254 12756 6666
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12728 5846 12756 6190
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12728 5098 12756 5646
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12820 5370 12848 5510
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 12912 5234 12940 6734
rect 12990 6352 13046 6361
rect 12990 6287 13046 6296
rect 13004 5914 13032 6287
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 13004 5302 13032 5510
rect 12992 5296 13044 5302
rect 12992 5238 13044 5244
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 12716 5092 12768 5098
rect 12716 5034 12768 5040
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12532 4548 12584 4554
rect 12532 4490 12584 4496
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12440 4004 12492 4010
rect 12440 3946 12492 3952
rect 12452 3534 12480 3946
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12256 3120 12308 3126
rect 12256 3062 12308 3068
rect 12162 2816 12218 2825
rect 12162 2751 12218 2760
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 12176 2310 12204 2586
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 12268 800 12296 3062
rect 12452 2446 12480 3470
rect 12544 3194 12572 4490
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12624 3120 12676 3126
rect 12622 3088 12624 3097
rect 12676 3088 12678 3097
rect 12622 3023 12678 3032
rect 12532 2916 12584 2922
rect 12532 2858 12584 2864
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 12544 800 12572 2858
rect 12728 800 12756 4490
rect 12820 3670 12848 4558
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 12808 3664 12860 3670
rect 12808 3606 12860 3612
rect 13004 800 13032 3878
rect 13096 3058 13124 9574
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13188 9110 13216 9454
rect 13176 9104 13228 9110
rect 13176 9046 13228 9052
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13188 8634 13216 8910
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13188 8401 13216 8434
rect 13174 8392 13230 8401
rect 13174 8327 13230 8336
rect 13174 8256 13230 8265
rect 13174 8191 13230 8200
rect 13188 4554 13216 8191
rect 13280 8090 13308 12242
rect 13372 8838 13400 14436
rect 13464 12306 13492 19366
rect 13556 17202 13584 20266
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13544 16720 13596 16726
rect 13544 16662 13596 16668
rect 13556 16114 13584 16662
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13556 15910 13584 16050
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13542 14920 13598 14929
rect 13542 14855 13598 14864
rect 13556 14006 13584 14855
rect 13544 14000 13596 14006
rect 13544 13942 13596 13948
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13556 12782 13584 13262
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13464 11150 13492 11630
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13450 10976 13506 10985
rect 13450 10911 13506 10920
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13464 8498 13492 10911
rect 13556 10674 13584 11154
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13542 10024 13598 10033
rect 13542 9959 13598 9968
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13372 7954 13400 8230
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13360 6928 13412 6934
rect 13360 6870 13412 6876
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13280 6390 13308 6598
rect 13372 6390 13400 6870
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 13360 6384 13412 6390
rect 13360 6326 13412 6332
rect 13464 5930 13492 8026
rect 13556 8022 13584 9959
rect 13648 9602 13676 22335
rect 13832 22094 13860 25860
rect 13912 25842 13964 25848
rect 13924 24614 13952 25842
rect 14016 25838 14044 26182
rect 14108 26042 14136 26318
rect 14096 26036 14148 26042
rect 14096 25978 14148 25984
rect 14280 25968 14332 25974
rect 14280 25910 14332 25916
rect 14004 25832 14056 25838
rect 14004 25774 14056 25780
rect 14292 25430 14320 25910
rect 14832 25696 14884 25702
rect 14832 25638 14884 25644
rect 14428 25596 14736 25616
rect 14428 25594 14434 25596
rect 14490 25594 14514 25596
rect 14570 25594 14594 25596
rect 14650 25594 14674 25596
rect 14730 25594 14736 25596
rect 14490 25542 14492 25594
rect 14672 25542 14674 25594
rect 14428 25540 14434 25542
rect 14490 25540 14514 25542
rect 14570 25540 14594 25542
rect 14650 25540 14674 25542
rect 14730 25540 14736 25542
rect 14428 25520 14736 25540
rect 14844 25430 14872 25638
rect 14280 25424 14332 25430
rect 14280 25366 14332 25372
rect 14832 25424 14884 25430
rect 14832 25366 14884 25372
rect 14188 25220 14240 25226
rect 14188 25162 14240 25168
rect 14200 24818 14228 25162
rect 14188 24812 14240 24818
rect 14188 24754 14240 24760
rect 13912 24608 13964 24614
rect 13912 24550 13964 24556
rect 14428 24508 14736 24528
rect 14428 24506 14434 24508
rect 14490 24506 14514 24508
rect 14570 24506 14594 24508
rect 14650 24506 14674 24508
rect 14730 24506 14736 24508
rect 14490 24454 14492 24506
rect 14672 24454 14674 24506
rect 14428 24452 14434 24454
rect 14490 24452 14514 24454
rect 14570 24452 14594 24454
rect 14650 24452 14674 24454
rect 14730 24452 14736 24454
rect 14428 24432 14736 24452
rect 14832 24404 14884 24410
rect 14832 24346 14884 24352
rect 14188 24200 14240 24206
rect 14188 24142 14240 24148
rect 14740 24200 14792 24206
rect 14740 24142 14792 24148
rect 14004 23520 14056 23526
rect 14004 23462 14056 23468
rect 14016 23186 14044 23462
rect 14004 23180 14056 23186
rect 14004 23122 14056 23128
rect 14016 22438 14044 23122
rect 14096 23044 14148 23050
rect 14096 22986 14148 22992
rect 14108 22642 14136 22986
rect 14200 22964 14228 24142
rect 14752 23730 14780 24142
rect 14740 23724 14792 23730
rect 14740 23666 14792 23672
rect 14280 23588 14332 23594
rect 14280 23530 14332 23536
rect 14292 23118 14320 23530
rect 14428 23420 14736 23440
rect 14428 23418 14434 23420
rect 14490 23418 14514 23420
rect 14570 23418 14594 23420
rect 14650 23418 14674 23420
rect 14730 23418 14736 23420
rect 14490 23366 14492 23418
rect 14672 23366 14674 23418
rect 14428 23364 14434 23366
rect 14490 23364 14514 23366
rect 14570 23364 14594 23366
rect 14650 23364 14674 23366
rect 14730 23364 14736 23366
rect 14428 23344 14736 23364
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 14280 22976 14332 22982
rect 14200 22936 14280 22964
rect 14280 22918 14332 22924
rect 14464 22976 14516 22982
rect 14464 22918 14516 22924
rect 14096 22636 14148 22642
rect 14096 22578 14148 22584
rect 14188 22636 14240 22642
rect 14188 22578 14240 22584
rect 14004 22432 14056 22438
rect 14004 22374 14056 22380
rect 14016 22234 14044 22374
rect 14004 22228 14056 22234
rect 14004 22170 14056 22176
rect 14108 22166 14136 22578
rect 14200 22234 14228 22578
rect 14188 22228 14240 22234
rect 14188 22170 14240 22176
rect 14096 22160 14148 22166
rect 14096 22102 14148 22108
rect 13832 22066 14044 22094
rect 13912 22024 13964 22030
rect 13912 21966 13964 21972
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13832 20874 13860 21490
rect 13820 20868 13872 20874
rect 13820 20810 13872 20816
rect 13832 20466 13860 20810
rect 13820 20460 13872 20466
rect 13820 20402 13872 20408
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13728 19780 13780 19786
rect 13728 19722 13780 19728
rect 13740 19242 13768 19722
rect 13832 19378 13860 20198
rect 13924 19553 13952 21966
rect 14016 21146 14044 22066
rect 14096 22024 14148 22030
rect 14148 21984 14228 22012
rect 14096 21966 14148 21972
rect 14096 21888 14148 21894
rect 14096 21830 14148 21836
rect 14004 21140 14056 21146
rect 14004 21082 14056 21088
rect 14016 21049 14044 21082
rect 14002 21040 14058 21049
rect 14002 20975 14058 20984
rect 14004 20528 14056 20534
rect 14004 20470 14056 20476
rect 14016 20058 14044 20470
rect 14004 20052 14056 20058
rect 14004 19994 14056 20000
rect 14108 19825 14136 21830
rect 14200 21060 14228 21984
rect 14292 21350 14320 22918
rect 14476 22642 14504 22918
rect 14464 22636 14516 22642
rect 14464 22578 14516 22584
rect 14428 22332 14736 22352
rect 14428 22330 14434 22332
rect 14490 22330 14514 22332
rect 14570 22330 14594 22332
rect 14650 22330 14674 22332
rect 14730 22330 14736 22332
rect 14490 22278 14492 22330
rect 14672 22278 14674 22330
rect 14428 22276 14434 22278
rect 14490 22276 14514 22278
rect 14570 22276 14594 22278
rect 14650 22276 14674 22278
rect 14730 22276 14736 22278
rect 14428 22256 14736 22276
rect 14372 22160 14424 22166
rect 14372 22102 14424 22108
rect 14384 22030 14412 22102
rect 14372 22024 14424 22030
rect 14372 21966 14424 21972
rect 14740 22024 14792 22030
rect 14740 21966 14792 21972
rect 14752 21400 14780 21966
rect 14844 21962 14872 24346
rect 14832 21956 14884 21962
rect 14832 21898 14884 21904
rect 14844 21554 14872 21898
rect 14832 21548 14884 21554
rect 14832 21490 14884 21496
rect 14752 21372 14872 21400
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 14428 21244 14736 21264
rect 14428 21242 14434 21244
rect 14490 21242 14514 21244
rect 14570 21242 14594 21244
rect 14650 21242 14674 21244
rect 14730 21242 14736 21244
rect 14490 21190 14492 21242
rect 14672 21190 14674 21242
rect 14428 21188 14434 21190
rect 14490 21188 14514 21190
rect 14570 21188 14594 21190
rect 14650 21188 14674 21190
rect 14730 21188 14736 21190
rect 14428 21168 14736 21188
rect 14200 21032 14320 21060
rect 14188 20460 14240 20466
rect 14188 20402 14240 20408
rect 14200 20097 14228 20402
rect 14186 20088 14242 20097
rect 14186 20023 14242 20032
rect 14292 19990 14320 21032
rect 14428 20156 14736 20176
rect 14428 20154 14434 20156
rect 14490 20154 14514 20156
rect 14570 20154 14594 20156
rect 14650 20154 14674 20156
rect 14730 20154 14736 20156
rect 14490 20102 14492 20154
rect 14672 20102 14674 20154
rect 14428 20100 14434 20102
rect 14490 20100 14514 20102
rect 14570 20100 14594 20102
rect 14650 20100 14674 20102
rect 14730 20100 14736 20102
rect 14428 20080 14736 20100
rect 14844 20040 14872 21372
rect 14752 20012 14872 20040
rect 14280 19984 14332 19990
rect 14280 19926 14332 19932
rect 14370 19952 14426 19961
rect 14292 19854 14320 19926
rect 14370 19887 14372 19896
rect 14424 19887 14426 19896
rect 14372 19858 14424 19864
rect 14280 19848 14332 19854
rect 14094 19816 14150 19825
rect 14280 19790 14332 19796
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14094 19751 14150 19760
rect 14186 19680 14242 19689
rect 14186 19615 14242 19624
rect 13910 19544 13966 19553
rect 13910 19479 13966 19488
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 13910 19272 13966 19281
rect 13728 19236 13780 19242
rect 13910 19207 13966 19216
rect 13728 19178 13780 19184
rect 13740 17882 13768 19178
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 13832 18222 13860 18702
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13728 17604 13780 17610
rect 13728 17546 13780 17552
rect 13740 17338 13768 17546
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13740 16522 13768 17138
rect 13728 16516 13780 16522
rect 13728 16458 13780 16464
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13740 15502 13768 16186
rect 13818 16144 13874 16153
rect 13818 16079 13820 16088
rect 13872 16079 13874 16088
rect 13820 16050 13872 16056
rect 13924 15994 13952 19207
rect 14016 18970 14044 19450
rect 14200 19378 14228 19615
rect 14476 19514 14504 19790
rect 14648 19712 14700 19718
rect 14646 19680 14648 19689
rect 14700 19680 14702 19689
rect 14646 19615 14702 19624
rect 14464 19508 14516 19514
rect 14464 19450 14516 19456
rect 14188 19372 14240 19378
rect 14240 19332 14320 19360
rect 14188 19314 14240 19320
rect 14096 19168 14148 19174
rect 14094 19136 14096 19145
rect 14148 19136 14150 19145
rect 14094 19071 14150 19080
rect 14186 19000 14242 19009
rect 14004 18964 14056 18970
rect 14004 18906 14056 18912
rect 14096 18964 14148 18970
rect 14186 18935 14242 18944
rect 14096 18906 14148 18912
rect 14004 18828 14056 18834
rect 14004 18770 14056 18776
rect 14016 18358 14044 18770
rect 14108 18766 14136 18906
rect 14200 18902 14228 18935
rect 14188 18896 14240 18902
rect 14188 18838 14240 18844
rect 14292 18834 14320 19332
rect 14476 19242 14504 19450
rect 14464 19236 14516 19242
rect 14464 19178 14516 19184
rect 14752 19156 14780 20012
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14844 19281 14872 19314
rect 14830 19272 14886 19281
rect 14830 19207 14886 19216
rect 14752 19128 14872 19156
rect 14428 19068 14736 19088
rect 14428 19066 14434 19068
rect 14490 19066 14514 19068
rect 14570 19066 14594 19068
rect 14650 19066 14674 19068
rect 14730 19066 14736 19068
rect 14490 19014 14492 19066
rect 14672 19014 14674 19066
rect 14428 19012 14434 19014
rect 14490 19012 14514 19014
rect 14570 19012 14594 19014
rect 14650 19012 14674 19014
rect 14730 19012 14736 19014
rect 14428 18992 14736 19012
rect 14844 18952 14872 19128
rect 14752 18924 14872 18952
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14096 18760 14148 18766
rect 14096 18702 14148 18708
rect 14004 18352 14056 18358
rect 14004 18294 14056 18300
rect 14108 18290 14136 18702
rect 14752 18306 14780 18924
rect 14830 18728 14886 18737
rect 14830 18663 14886 18672
rect 14844 18426 14872 18663
rect 14832 18420 14884 18426
rect 14832 18362 14884 18368
rect 14096 18284 14148 18290
rect 14752 18278 14872 18306
rect 14096 18226 14148 18232
rect 14094 18048 14150 18057
rect 14094 17983 14150 17992
rect 14004 16720 14056 16726
rect 14004 16662 14056 16668
rect 13832 15966 13952 15994
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13740 15162 13768 15438
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13740 14385 13768 14962
rect 13726 14376 13782 14385
rect 13726 14311 13782 14320
rect 13740 12481 13768 14311
rect 13726 12472 13782 12481
rect 13726 12407 13782 12416
rect 13832 12102 13860 15966
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13924 14482 13952 15846
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 14016 12986 14044 16662
rect 14108 13530 14136 17983
rect 14428 17980 14736 18000
rect 14428 17978 14434 17980
rect 14490 17978 14514 17980
rect 14570 17978 14594 17980
rect 14650 17978 14674 17980
rect 14730 17978 14736 17980
rect 14490 17926 14492 17978
rect 14672 17926 14674 17978
rect 14428 17924 14434 17926
rect 14490 17924 14514 17926
rect 14570 17924 14594 17926
rect 14650 17924 14674 17926
rect 14730 17924 14736 17926
rect 14428 17904 14736 17924
rect 14844 17882 14872 18278
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14844 17270 14872 17818
rect 14832 17264 14884 17270
rect 14370 17232 14426 17241
rect 14832 17206 14884 17212
rect 14370 17167 14372 17176
rect 14424 17167 14426 17176
rect 14372 17138 14424 17144
rect 14428 16892 14736 16912
rect 14428 16890 14434 16892
rect 14490 16890 14514 16892
rect 14570 16890 14594 16892
rect 14650 16890 14674 16892
rect 14730 16890 14736 16892
rect 14490 16838 14492 16890
rect 14672 16838 14674 16890
rect 14428 16836 14434 16838
rect 14490 16836 14514 16838
rect 14570 16836 14594 16838
rect 14650 16836 14674 16838
rect 14730 16836 14736 16838
rect 14428 16816 14736 16836
rect 14832 16584 14884 16590
rect 14832 16526 14884 16532
rect 14372 16516 14424 16522
rect 14372 16458 14424 16464
rect 14384 16250 14412 16458
rect 14844 16425 14872 16526
rect 14830 16416 14886 16425
rect 14830 16351 14886 16360
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 14384 16017 14412 16050
rect 14370 16008 14426 16017
rect 14370 15943 14426 15952
rect 14428 15804 14736 15824
rect 14428 15802 14434 15804
rect 14490 15802 14514 15804
rect 14570 15802 14594 15804
rect 14650 15802 14674 15804
rect 14730 15802 14736 15804
rect 14490 15750 14492 15802
rect 14672 15750 14674 15802
rect 14428 15748 14434 15750
rect 14490 15748 14514 15750
rect 14570 15748 14594 15750
rect 14650 15748 14674 15750
rect 14730 15748 14736 15750
rect 14428 15728 14736 15748
rect 14646 15600 14702 15609
rect 14646 15535 14702 15544
rect 14188 15496 14240 15502
rect 14372 15496 14424 15502
rect 14188 15438 14240 15444
rect 14292 15456 14372 15484
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14002 12880 14058 12889
rect 14002 12815 14058 12824
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13740 11626 13768 12038
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13820 11552 13872 11558
rect 13740 11500 13820 11506
rect 13740 11494 13872 11500
rect 13740 11478 13860 11494
rect 13740 11354 13768 11478
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13648 9574 13768 9602
rect 13636 8900 13688 8906
rect 13636 8842 13688 8848
rect 13648 8634 13676 8842
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13544 8016 13596 8022
rect 13544 7958 13596 7964
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13556 7410 13584 7822
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13556 6118 13584 6938
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13372 5902 13492 5930
rect 13176 4548 13228 4554
rect 13176 4490 13228 4496
rect 13268 4480 13320 4486
rect 13268 4422 13320 4428
rect 13176 4276 13228 4282
rect 13176 4218 13228 4224
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 13188 2854 13216 4218
rect 13280 4078 13308 4422
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 13372 4010 13400 5902
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 13556 5710 13584 5782
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13648 5148 13676 8434
rect 13740 6866 13768 9574
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13740 5914 13768 6054
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13832 5760 13860 11290
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13924 10810 13952 11086
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13924 9926 13952 10746
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13910 8664 13966 8673
rect 13910 8599 13966 8608
rect 13924 8498 13952 8599
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13924 7206 13952 8230
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 13912 6384 13964 6390
rect 13912 6326 13964 6332
rect 13924 6118 13952 6326
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 13740 5732 13860 5760
rect 13740 5250 13768 5732
rect 13912 5636 13964 5642
rect 13912 5578 13964 5584
rect 13740 5222 13860 5250
rect 13924 5234 13952 5578
rect 13648 5120 13768 5148
rect 13360 4004 13412 4010
rect 13360 3946 13412 3952
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13280 3194 13308 3470
rect 13544 3392 13596 3398
rect 13464 3352 13544 3380
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 13280 2446 13308 2586
rect 13372 2514 13400 2926
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13464 2292 13492 3352
rect 13544 3334 13596 3340
rect 13648 2774 13676 3878
rect 13280 2264 13492 2292
rect 13556 2746 13676 2774
rect 13280 800 13308 2264
rect 13556 800 13584 2746
rect 13740 2650 13768 5120
rect 13832 5114 13860 5222
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 13832 5086 13952 5114
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13832 4146 13860 4422
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 13924 2514 13952 5086
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 14016 2394 14044 12815
rect 14108 11914 14136 13126
rect 14200 12073 14228 15438
rect 14292 13512 14320 15456
rect 14372 15438 14424 15444
rect 14554 15464 14610 15473
rect 14660 15434 14688 15535
rect 14740 15496 14792 15502
rect 14844 15484 14872 16351
rect 14792 15456 14872 15484
rect 14740 15438 14792 15444
rect 14554 15399 14556 15408
rect 14608 15399 14610 15408
rect 14648 15428 14700 15434
rect 14556 15370 14608 15376
rect 14648 15370 14700 15376
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 14428 14716 14736 14736
rect 14428 14714 14434 14716
rect 14490 14714 14514 14716
rect 14570 14714 14594 14716
rect 14650 14714 14674 14716
rect 14730 14714 14736 14716
rect 14490 14662 14492 14714
rect 14672 14662 14674 14714
rect 14428 14660 14434 14662
rect 14490 14660 14514 14662
rect 14570 14660 14594 14662
rect 14650 14660 14674 14662
rect 14730 14660 14736 14662
rect 14428 14640 14736 14660
rect 14844 14600 14872 14962
rect 14752 14572 14872 14600
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14476 14074 14504 14350
rect 14646 14104 14702 14113
rect 14464 14068 14516 14074
rect 14646 14039 14702 14048
rect 14464 14010 14516 14016
rect 14660 14006 14688 14039
rect 14648 14000 14700 14006
rect 14648 13942 14700 13948
rect 14752 13802 14780 14572
rect 14832 14476 14884 14482
rect 14832 14418 14884 14424
rect 14740 13796 14792 13802
rect 14740 13738 14792 13744
rect 14428 13628 14736 13648
rect 14428 13626 14434 13628
rect 14490 13626 14514 13628
rect 14570 13626 14594 13628
rect 14650 13626 14674 13628
rect 14730 13626 14736 13628
rect 14490 13574 14492 13626
rect 14672 13574 14674 13626
rect 14428 13572 14434 13574
rect 14490 13572 14514 13574
rect 14570 13572 14594 13574
rect 14650 13572 14674 13574
rect 14730 13572 14736 13574
rect 14428 13552 14736 13572
rect 14292 13484 14412 13512
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14292 12918 14320 13262
rect 14280 12912 14332 12918
rect 14280 12854 14332 12860
rect 14384 12714 14412 13484
rect 14844 12850 14872 14418
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14372 12708 14424 12714
rect 14936 12696 14964 27270
rect 15028 21457 15056 28494
rect 15568 28416 15620 28422
rect 15568 28358 15620 28364
rect 15292 27872 15344 27878
rect 15292 27814 15344 27820
rect 15200 27328 15252 27334
rect 15200 27270 15252 27276
rect 15212 26353 15240 27270
rect 15198 26344 15254 26353
rect 15198 26279 15254 26288
rect 15304 26228 15332 27814
rect 15384 26784 15436 26790
rect 15384 26726 15436 26732
rect 15396 26246 15424 26726
rect 15212 26200 15332 26228
rect 15384 26240 15436 26246
rect 15108 25696 15160 25702
rect 15108 25638 15160 25644
rect 15120 25498 15148 25638
rect 15108 25492 15160 25498
rect 15108 25434 15160 25440
rect 15212 25158 15240 26200
rect 15384 26182 15436 26188
rect 15292 25424 15344 25430
rect 15292 25366 15344 25372
rect 15200 25152 15252 25158
rect 15200 25094 15252 25100
rect 15212 24818 15240 25094
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15200 24200 15252 24206
rect 15200 24142 15252 24148
rect 15108 24064 15160 24070
rect 15108 24006 15160 24012
rect 15120 23118 15148 24006
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 15212 22710 15240 24142
rect 15200 22704 15252 22710
rect 15200 22646 15252 22652
rect 15304 22098 15332 25366
rect 15384 24676 15436 24682
rect 15384 24618 15436 24624
rect 15396 23798 15424 24618
rect 15384 23792 15436 23798
rect 15384 23734 15436 23740
rect 15108 22092 15160 22098
rect 15108 22034 15160 22040
rect 15292 22092 15344 22098
rect 15292 22034 15344 22040
rect 15014 21448 15070 21457
rect 15014 21383 15070 21392
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 15028 19854 15056 21286
rect 15120 20262 15148 22034
rect 15200 20868 15252 20874
rect 15200 20810 15252 20816
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 15212 20058 15240 20810
rect 15292 20460 15344 20466
rect 15292 20402 15344 20408
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15016 19848 15068 19854
rect 15016 19790 15068 19796
rect 15028 18766 15056 19790
rect 15304 19718 15332 20402
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15120 18952 15148 19654
rect 15120 18924 15164 18952
rect 15136 18884 15164 18924
rect 15120 18856 15164 18884
rect 15120 18816 15148 18856
rect 15120 18788 15332 18816
rect 15016 18760 15068 18766
rect 15016 18702 15068 18708
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 15212 18290 15240 18566
rect 15108 18284 15160 18290
rect 15108 18226 15160 18232
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 15016 18216 15068 18222
rect 15120 18193 15148 18226
rect 15016 18158 15068 18164
rect 15106 18184 15162 18193
rect 15028 17610 15056 18158
rect 15106 18119 15162 18128
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 15108 17808 15160 17814
rect 15108 17750 15160 17756
rect 15016 17604 15068 17610
rect 15016 17546 15068 17552
rect 15028 17270 15056 17546
rect 15016 17264 15068 17270
rect 15016 17206 15068 17212
rect 15016 16516 15068 16522
rect 15016 16458 15068 16464
rect 15028 16046 15056 16458
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 15028 15502 15056 15982
rect 15120 15745 15148 17750
rect 15106 15736 15162 15745
rect 15106 15671 15162 15680
rect 15108 15632 15160 15638
rect 15108 15574 15160 15580
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 15016 14816 15068 14822
rect 15016 14758 15068 14764
rect 15028 14550 15056 14758
rect 15016 14544 15068 14550
rect 15016 14486 15068 14492
rect 15016 14340 15068 14346
rect 15016 14282 15068 14288
rect 15028 14249 15056 14282
rect 15014 14240 15070 14249
rect 15014 14175 15070 14184
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 15028 13977 15056 14010
rect 15014 13968 15070 13977
rect 15014 13903 15070 13912
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 14372 12650 14424 12656
rect 14844 12668 14964 12696
rect 14428 12540 14736 12560
rect 14428 12538 14434 12540
rect 14490 12538 14514 12540
rect 14570 12538 14594 12540
rect 14650 12538 14674 12540
rect 14730 12538 14736 12540
rect 14490 12486 14492 12538
rect 14672 12486 14674 12538
rect 14428 12484 14434 12486
rect 14490 12484 14514 12486
rect 14570 12484 14594 12486
rect 14650 12484 14674 12486
rect 14730 12484 14736 12486
rect 14428 12464 14736 12484
rect 14186 12064 14242 12073
rect 14186 11999 14242 12008
rect 14646 11928 14702 11937
rect 14108 11898 14504 11914
rect 14108 11892 14516 11898
rect 14108 11886 14464 11892
rect 14108 11354 14136 11886
rect 14646 11863 14648 11872
rect 14464 11834 14516 11840
rect 14700 11863 14702 11872
rect 14648 11834 14700 11840
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 14292 11150 14320 11494
rect 14428 11452 14736 11472
rect 14428 11450 14434 11452
rect 14490 11450 14514 11452
rect 14570 11450 14594 11452
rect 14650 11450 14674 11452
rect 14730 11450 14736 11452
rect 14490 11398 14492 11450
rect 14672 11398 14674 11450
rect 14428 11396 14434 11398
rect 14490 11396 14514 11398
rect 14570 11396 14594 11398
rect 14650 11396 14674 11398
rect 14730 11396 14736 11398
rect 14428 11376 14736 11396
rect 14280 11144 14332 11150
rect 14332 11092 14412 11098
rect 14280 11086 14412 11092
rect 14292 11070 14412 11086
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14108 10266 14136 10610
rect 14200 10266 14228 10950
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14094 10160 14150 10169
rect 14094 10095 14150 10104
rect 14108 8265 14136 10095
rect 14292 10062 14320 10950
rect 14384 10742 14412 11070
rect 14372 10736 14424 10742
rect 14372 10678 14424 10684
rect 14428 10364 14736 10384
rect 14428 10362 14434 10364
rect 14490 10362 14514 10364
rect 14570 10362 14594 10364
rect 14650 10362 14674 10364
rect 14730 10362 14736 10364
rect 14490 10310 14492 10362
rect 14672 10310 14674 10362
rect 14428 10308 14434 10310
rect 14490 10308 14514 10310
rect 14570 10308 14594 10310
rect 14650 10308 14674 10310
rect 14730 10308 14736 10310
rect 14428 10288 14736 10308
rect 14844 10169 14872 12668
rect 15028 12628 15056 13466
rect 14936 12600 15056 12628
rect 14830 10160 14886 10169
rect 14648 10124 14700 10130
rect 14830 10095 14886 10104
rect 14648 10066 14700 10072
rect 14280 10056 14332 10062
rect 14186 10024 14242 10033
rect 14280 9998 14332 10004
rect 14186 9959 14242 9968
rect 14200 9926 14228 9959
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 14554 9888 14610 9897
rect 14554 9823 14610 9832
rect 14568 9466 14596 9823
rect 14660 9586 14688 10066
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14292 9438 14596 9466
rect 14094 8256 14150 8265
rect 14094 8191 14150 8200
rect 14186 8120 14242 8129
rect 14186 8055 14242 8064
rect 14200 8022 14228 8055
rect 14188 8016 14240 8022
rect 14188 7958 14240 7964
rect 14292 7562 14320 9438
rect 14832 9376 14884 9382
rect 14832 9318 14884 9324
rect 14428 9276 14736 9296
rect 14428 9274 14434 9276
rect 14490 9274 14514 9276
rect 14570 9274 14594 9276
rect 14650 9274 14674 9276
rect 14730 9274 14736 9276
rect 14490 9222 14492 9274
rect 14672 9222 14674 9274
rect 14428 9220 14434 9222
rect 14490 9220 14514 9222
rect 14570 9220 14594 9222
rect 14650 9220 14674 9222
rect 14730 9220 14736 9222
rect 14428 9200 14736 9220
rect 14844 8838 14872 9318
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 14428 8188 14736 8208
rect 14428 8186 14434 8188
rect 14490 8186 14514 8188
rect 14570 8186 14594 8188
rect 14650 8186 14674 8188
rect 14730 8186 14736 8188
rect 14490 8134 14492 8186
rect 14672 8134 14674 8186
rect 14428 8132 14434 8134
rect 14490 8132 14514 8134
rect 14570 8132 14594 8134
rect 14650 8132 14674 8134
rect 14730 8132 14736 8134
rect 14428 8112 14736 8132
rect 14844 8022 14872 8434
rect 14832 8016 14884 8022
rect 14370 7984 14426 7993
rect 14832 7958 14884 7964
rect 14370 7919 14426 7928
rect 14384 7886 14412 7919
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 14108 7534 14320 7562
rect 14108 4622 14136 7534
rect 14188 7472 14240 7478
rect 14188 7414 14240 7420
rect 14200 5846 14228 7414
rect 14428 7100 14736 7120
rect 14428 7098 14434 7100
rect 14490 7098 14514 7100
rect 14570 7098 14594 7100
rect 14650 7098 14674 7100
rect 14730 7098 14736 7100
rect 14490 7046 14492 7098
rect 14672 7046 14674 7098
rect 14428 7044 14434 7046
rect 14490 7044 14514 7046
rect 14570 7044 14594 7046
rect 14650 7044 14674 7046
rect 14730 7044 14736 7046
rect 14428 7024 14736 7044
rect 14936 7002 14964 12600
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 15028 10130 15056 10542
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 15120 9058 15148 15574
rect 15212 14346 15240 18022
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 15304 14074 15332 18788
rect 15396 16590 15424 23734
rect 15476 23112 15528 23118
rect 15476 23054 15528 23060
rect 15488 22710 15516 23054
rect 15476 22704 15528 22710
rect 15476 22646 15528 22652
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15488 19357 15516 20198
rect 15474 19348 15530 19357
rect 15474 19283 15530 19292
rect 15580 18952 15608 28358
rect 15660 27328 15712 27334
rect 15660 27270 15712 27276
rect 15672 27130 15700 27270
rect 15660 27124 15712 27130
rect 15660 27066 15712 27072
rect 15660 24608 15712 24614
rect 15660 24550 15712 24556
rect 15672 23866 15700 24550
rect 15660 23860 15712 23866
rect 15660 23802 15712 23808
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15672 22642 15700 23054
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 15672 21593 15700 22578
rect 15658 21584 15714 21593
rect 15658 21519 15714 21528
rect 15660 20528 15712 20534
rect 15660 20470 15712 20476
rect 15672 19990 15700 20470
rect 15660 19984 15712 19990
rect 15660 19926 15712 19932
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15672 19224 15700 19790
rect 15764 19352 15792 28698
rect 16488 28552 16540 28558
rect 16488 28494 16540 28500
rect 16120 28212 16172 28218
rect 16120 28154 16172 28160
rect 16028 27464 16080 27470
rect 16028 27406 16080 27412
rect 15844 26784 15896 26790
rect 15844 26726 15896 26732
rect 15936 26784 15988 26790
rect 15936 26726 15988 26732
rect 15856 25906 15884 26726
rect 15948 26330 15976 26726
rect 16040 26586 16068 27406
rect 16028 26580 16080 26586
rect 16028 26522 16080 26528
rect 15948 26302 16068 26330
rect 15936 26240 15988 26246
rect 15936 26182 15988 26188
rect 15844 25900 15896 25906
rect 15844 25842 15896 25848
rect 15948 25702 15976 26182
rect 15936 25696 15988 25702
rect 15936 25638 15988 25644
rect 15844 25288 15896 25294
rect 15844 25230 15896 25236
rect 15856 24274 15884 25230
rect 15844 24268 15896 24274
rect 15844 24210 15896 24216
rect 15936 24132 15988 24138
rect 15936 24074 15988 24080
rect 15844 22092 15896 22098
rect 15844 22034 15896 22040
rect 15856 20398 15884 22034
rect 15844 20392 15896 20398
rect 15844 20334 15896 20340
rect 15948 19961 15976 24074
rect 16040 22506 16068 26302
rect 16028 22500 16080 22506
rect 16028 22442 16080 22448
rect 16132 22094 16160 28154
rect 16500 26518 16528 28494
rect 16580 27328 16632 27334
rect 16580 27270 16632 27276
rect 16488 26512 16540 26518
rect 16488 26454 16540 26460
rect 16488 25696 16540 25702
rect 16488 25638 16540 25644
rect 16304 25424 16356 25430
rect 16304 25366 16356 25372
rect 16132 22066 16252 22094
rect 16120 21888 16172 21894
rect 16120 21830 16172 21836
rect 16132 21554 16160 21830
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 16028 20324 16080 20330
rect 16028 20266 16080 20272
rect 15934 19952 15990 19961
rect 15934 19887 15990 19896
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15752 19346 15804 19352
rect 15856 19334 15884 19654
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 15856 19306 15900 19334
rect 15752 19288 15804 19294
rect 15672 19196 15792 19224
rect 15580 18924 15700 18952
rect 15672 18612 15700 18924
rect 15580 18584 15700 18612
rect 15474 16824 15530 16833
rect 15474 16759 15530 16768
rect 15384 16584 15436 16590
rect 15384 16526 15436 16532
rect 15384 15632 15436 15638
rect 15384 15574 15436 15580
rect 15396 15337 15424 15574
rect 15382 15328 15438 15337
rect 15382 15263 15438 15272
rect 15488 14929 15516 16759
rect 15474 14920 15530 14929
rect 15384 14884 15436 14890
rect 15474 14855 15530 14864
rect 15384 14826 15436 14832
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15200 12708 15252 12714
rect 15200 12650 15252 12656
rect 15212 11694 15240 12650
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 15304 11558 15332 13670
rect 15396 13326 15424 14826
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15488 14074 15516 14214
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15474 13968 15530 13977
rect 15474 13903 15530 13912
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15488 13172 15516 13903
rect 15396 13144 15516 13172
rect 15292 11552 15344 11558
rect 15198 11520 15254 11529
rect 15292 11494 15344 11500
rect 15198 11455 15254 11464
rect 15028 9030 15148 9058
rect 14924 6996 14976 7002
rect 14924 6938 14976 6944
rect 15028 6848 15056 9030
rect 15108 8900 15160 8906
rect 15108 8842 15160 8848
rect 15120 8090 15148 8842
rect 15212 8566 15240 11455
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15304 10062 15332 10406
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15200 8560 15252 8566
rect 15200 8502 15252 8508
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15304 7886 15332 8298
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15028 6820 15148 6848
rect 14924 6792 14976 6798
rect 14976 6752 15056 6780
rect 14924 6734 14976 6740
rect 14280 6724 14332 6730
rect 14280 6666 14332 6672
rect 14188 5840 14240 5846
rect 14188 5782 14240 5788
rect 14292 5234 14320 6666
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 14740 6248 14792 6254
rect 14738 6216 14740 6225
rect 14792 6216 14794 6225
rect 14738 6151 14794 6160
rect 14428 6012 14736 6032
rect 14428 6010 14434 6012
rect 14490 6010 14514 6012
rect 14570 6010 14594 6012
rect 14650 6010 14674 6012
rect 14730 6010 14736 6012
rect 14490 5958 14492 6010
rect 14672 5958 14674 6010
rect 14428 5956 14434 5958
rect 14490 5956 14514 5958
rect 14570 5956 14594 5958
rect 14650 5956 14674 5958
rect 14730 5956 14736 5958
rect 14428 5936 14736 5956
rect 14370 5808 14426 5817
rect 14844 5778 14872 6258
rect 14370 5743 14426 5752
rect 14832 5772 14884 5778
rect 14280 5228 14332 5234
rect 14200 5188 14280 5216
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14096 4004 14148 4010
rect 14096 3946 14148 3952
rect 13832 2366 14044 2394
rect 13832 800 13860 2366
rect 14108 800 14136 3946
rect 14200 3534 14228 5188
rect 14280 5170 14332 5176
rect 14384 5114 14412 5743
rect 14832 5714 14884 5720
rect 14292 5086 14412 5114
rect 14188 3528 14240 3534
rect 14292 3516 14320 5086
rect 14428 4924 14736 4944
rect 14428 4922 14434 4924
rect 14490 4922 14514 4924
rect 14570 4922 14594 4924
rect 14650 4922 14674 4924
rect 14730 4922 14736 4924
rect 14490 4870 14492 4922
rect 14672 4870 14674 4922
rect 14428 4868 14434 4870
rect 14490 4868 14514 4870
rect 14570 4868 14594 4870
rect 14650 4868 14674 4870
rect 14730 4868 14736 4870
rect 14428 4848 14736 4868
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14428 3836 14736 3856
rect 14428 3834 14434 3836
rect 14490 3834 14514 3836
rect 14570 3834 14594 3836
rect 14650 3834 14674 3836
rect 14730 3834 14736 3836
rect 14490 3782 14492 3834
rect 14672 3782 14674 3834
rect 14428 3780 14434 3782
rect 14490 3780 14514 3782
rect 14570 3780 14594 3782
rect 14650 3780 14674 3782
rect 14730 3780 14736 3782
rect 14428 3760 14736 3780
rect 14372 3528 14424 3534
rect 14292 3488 14372 3516
rect 14188 3470 14240 3476
rect 14372 3470 14424 3476
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14292 1986 14320 3130
rect 14428 2748 14736 2768
rect 14428 2746 14434 2748
rect 14490 2746 14514 2748
rect 14570 2746 14594 2748
rect 14650 2746 14674 2748
rect 14730 2746 14736 2748
rect 14490 2694 14492 2746
rect 14672 2694 14674 2746
rect 14428 2692 14434 2694
rect 14490 2692 14514 2694
rect 14570 2692 14594 2694
rect 14650 2692 14674 2694
rect 14730 2692 14736 2694
rect 14428 2672 14736 2692
rect 14844 2258 14872 4422
rect 14936 4146 14964 6598
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 15028 4026 15056 6752
rect 15120 5817 15148 6820
rect 15212 6440 15240 7346
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15304 6730 15332 7142
rect 15292 6724 15344 6730
rect 15292 6666 15344 6672
rect 15292 6452 15344 6458
rect 15212 6412 15292 6440
rect 15292 6394 15344 6400
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15304 5930 15332 6190
rect 15212 5902 15332 5930
rect 15106 5808 15162 5817
rect 15106 5743 15162 5752
rect 15108 5636 15160 5642
rect 15212 5624 15240 5902
rect 15160 5596 15240 5624
rect 15292 5636 15344 5642
rect 15108 5578 15160 5584
rect 15396 5624 15424 13144
rect 15474 13016 15530 13025
rect 15474 12951 15530 12960
rect 15488 8838 15516 12951
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15488 7750 15516 8774
rect 15580 8480 15608 18584
rect 15764 18426 15792 19196
rect 15872 19145 15900 19306
rect 15858 19136 15914 19145
rect 15858 19071 15914 19080
rect 15948 18766 15976 19450
rect 15936 18760 15988 18766
rect 15936 18702 15988 18708
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 15750 18048 15806 18057
rect 15750 17983 15806 17992
rect 15660 17876 15712 17882
rect 15660 17818 15712 17824
rect 15672 16697 15700 17818
rect 15658 16688 15714 16697
rect 15658 16623 15714 16632
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 15672 15502 15700 16526
rect 15764 16522 15792 17983
rect 15948 17882 15976 18226
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 15936 17196 15988 17202
rect 15936 17138 15988 17144
rect 15948 16794 15976 17138
rect 15936 16788 15988 16794
rect 15936 16730 15988 16736
rect 15948 16658 15976 16730
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 15934 16552 15990 16561
rect 15752 16516 15804 16522
rect 15934 16487 15936 16496
rect 15752 16458 15804 16464
rect 15988 16487 15990 16496
rect 15936 16458 15988 16464
rect 15750 16416 15806 16425
rect 16040 16402 16068 20266
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 15750 16351 15806 16360
rect 15856 16374 16068 16402
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15658 15192 15714 15201
rect 15658 15127 15714 15136
rect 15672 14006 15700 15127
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15672 12782 15700 13262
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15672 10538 15700 10610
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15672 9994 15700 10474
rect 15660 9988 15712 9994
rect 15660 9930 15712 9936
rect 15580 8452 15700 8480
rect 15568 8356 15620 8362
rect 15568 8298 15620 8304
rect 15580 7818 15608 8298
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15672 7426 15700 8452
rect 15764 7562 15792 16351
rect 15856 15706 15884 16374
rect 16132 16046 16160 19314
rect 16224 19258 16252 22066
rect 16316 22030 16344 25366
rect 16396 25288 16448 25294
rect 16396 25230 16448 25236
rect 16408 23322 16436 25230
rect 16396 23316 16448 23322
rect 16396 23258 16448 23264
rect 16500 23118 16528 25638
rect 16592 23508 16620 27270
rect 16684 24857 16712 28698
rect 18328 28688 18380 28694
rect 18328 28630 18380 28636
rect 20168 28688 20220 28694
rect 20168 28630 20220 28636
rect 22100 28688 22152 28694
rect 22100 28630 22152 28636
rect 17592 28552 17644 28558
rect 17592 28494 17644 28500
rect 18144 28552 18196 28558
rect 18144 28494 18196 28500
rect 16856 28416 16908 28422
rect 16856 28358 16908 28364
rect 17316 28416 17368 28422
rect 17316 28358 17368 28364
rect 16764 28076 16816 28082
rect 16868 28064 16896 28358
rect 16948 28076 17000 28082
rect 16868 28036 16948 28064
rect 16764 28018 16816 28024
rect 16948 28018 17000 28024
rect 16776 26994 16804 28018
rect 17132 27396 17184 27402
rect 17132 27338 17184 27344
rect 17040 27328 17092 27334
rect 17040 27270 17092 27276
rect 16764 26988 16816 26994
rect 16764 26930 16816 26936
rect 16670 24848 16726 24857
rect 16670 24783 16726 24792
rect 16672 24200 16724 24206
rect 16672 24142 16724 24148
rect 16684 23662 16712 24142
rect 16672 23656 16724 23662
rect 16672 23598 16724 23604
rect 16592 23480 16712 23508
rect 16488 23112 16540 23118
rect 16488 23054 16540 23060
rect 16500 22574 16528 23054
rect 16488 22568 16540 22574
rect 16488 22510 16540 22516
rect 16488 22432 16540 22438
rect 16488 22374 16540 22380
rect 16500 22098 16528 22374
rect 16488 22092 16540 22098
rect 16488 22034 16540 22040
rect 16304 22024 16356 22030
rect 16304 21966 16356 21972
rect 16304 20936 16356 20942
rect 16304 20878 16356 20884
rect 16316 19854 16344 20878
rect 16396 20392 16448 20398
rect 16396 20334 16448 20340
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 16316 19446 16344 19790
rect 16304 19440 16356 19446
rect 16304 19382 16356 19388
rect 16224 19230 16344 19258
rect 16212 18896 16264 18902
rect 16212 18838 16264 18844
rect 16224 18465 16252 18838
rect 16210 18456 16266 18465
rect 16210 18391 16266 18400
rect 16212 16720 16264 16726
rect 16212 16662 16264 16668
rect 16224 16182 16252 16662
rect 16212 16176 16264 16182
rect 16212 16118 16264 16124
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 15936 15972 15988 15978
rect 15936 15914 15988 15920
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15844 15564 15896 15570
rect 15844 15506 15896 15512
rect 15856 15162 15884 15506
rect 15948 15366 15976 15914
rect 16028 15700 16080 15706
rect 16028 15642 16080 15648
rect 15936 15360 15988 15366
rect 15936 15302 15988 15308
rect 15844 15156 15896 15162
rect 15844 15098 15896 15104
rect 15856 14346 15884 15098
rect 16040 14822 16068 15642
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 16040 14618 16068 14758
rect 16028 14612 16080 14618
rect 16028 14554 16080 14560
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 15844 14340 15896 14346
rect 15844 14282 15896 14288
rect 15842 13832 15898 13841
rect 15842 13767 15898 13776
rect 15856 13734 15884 13767
rect 15844 13728 15896 13734
rect 15844 13670 15896 13676
rect 15948 13394 15976 14350
rect 15936 13388 15988 13394
rect 15936 13330 15988 13336
rect 15844 13252 15896 13258
rect 15844 13194 15896 13200
rect 15936 13252 15988 13258
rect 15936 13194 15988 13200
rect 15856 12889 15884 13194
rect 15842 12880 15898 12889
rect 15842 12815 15898 12824
rect 15948 12442 15976 13194
rect 16040 12918 16068 14350
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 16028 12640 16080 12646
rect 16028 12582 16080 12588
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 15934 12336 15990 12345
rect 15934 12271 15990 12280
rect 15948 12170 15976 12271
rect 15936 12164 15988 12170
rect 15936 12106 15988 12112
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15856 11626 15884 12038
rect 15936 11824 15988 11830
rect 15936 11766 15988 11772
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 15948 11529 15976 11766
rect 15934 11520 15990 11529
rect 15934 11455 15990 11464
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 15856 10810 15884 11290
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15856 10674 15884 10746
rect 16040 10713 16068 12582
rect 16132 11286 16160 15982
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 16224 15201 16252 15642
rect 16210 15192 16266 15201
rect 16210 15127 16266 15136
rect 16212 14884 16264 14890
rect 16212 14826 16264 14832
rect 16224 12646 16252 14826
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16120 11280 16172 11286
rect 16120 11222 16172 11228
rect 16026 10704 16082 10713
rect 15844 10668 15896 10674
rect 16026 10639 16082 10648
rect 15844 10610 15896 10616
rect 16132 10130 16160 11222
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 16224 10010 16252 12038
rect 16132 9982 16252 10010
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 15856 9178 15884 9522
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15842 9072 15898 9081
rect 15842 9007 15898 9016
rect 15856 8566 15884 9007
rect 15948 8634 15976 9114
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 15844 8560 15896 8566
rect 15844 8502 15896 8508
rect 15844 8424 15896 8430
rect 15842 8392 15844 8401
rect 15896 8392 15898 8401
rect 15842 8327 15898 8336
rect 15764 7534 16068 7562
rect 15672 7398 15884 7426
rect 15660 7336 15712 7342
rect 15660 7278 15712 7284
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15344 5596 15424 5624
rect 15292 5578 15344 5584
rect 15396 5030 15424 5596
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15488 4622 15516 7142
rect 15568 6724 15620 6730
rect 15568 6666 15620 6672
rect 15580 6361 15608 6666
rect 15566 6352 15622 6361
rect 15566 6287 15622 6296
rect 15672 5846 15700 7278
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 15660 5840 15712 5846
rect 15660 5782 15712 5788
rect 15764 5710 15792 6938
rect 15752 5704 15804 5710
rect 15658 5672 15714 5681
rect 15752 5646 15804 5652
rect 15658 5607 15714 5616
rect 15672 5574 15700 5607
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 15672 5370 15700 5510
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 15476 4616 15528 4622
rect 15476 4558 15528 4564
rect 15292 4548 15344 4554
rect 15292 4490 15344 4496
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 14936 3998 15056 4026
rect 14936 2650 14964 3998
rect 15108 3664 15160 3670
rect 15108 3606 15160 3612
rect 15016 3460 15068 3466
rect 15016 3402 15068 3408
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 14660 2230 14872 2258
rect 14292 1958 14412 1986
rect 14384 800 14412 1958
rect 14660 800 14688 2230
rect 15028 1714 15056 3402
rect 15120 3194 15148 3606
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 14936 1686 15056 1714
rect 14936 800 14964 1686
rect 15212 800 15240 4422
rect 15304 3194 15332 4490
rect 15752 4004 15804 4010
rect 15752 3946 15804 3952
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15476 3120 15528 3126
rect 15476 3062 15528 3068
rect 15384 2916 15436 2922
rect 15384 2858 15436 2864
rect 15396 2650 15424 2858
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 15488 800 15516 3062
rect 15764 800 15792 3946
rect 15856 3398 15884 7398
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15948 6225 15976 6598
rect 15934 6216 15990 6225
rect 15934 6151 15990 6160
rect 15844 3392 15896 3398
rect 15844 3334 15896 3340
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 15948 2650 15976 2926
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 16040 800 16068 7534
rect 16132 7528 16160 9982
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16224 7886 16252 8366
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 16316 7818 16344 19230
rect 16408 17882 16436 20334
rect 16500 19786 16528 22034
rect 16580 20256 16632 20262
rect 16580 20198 16632 20204
rect 16592 19854 16620 20198
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 16488 19780 16540 19786
rect 16488 19722 16540 19728
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16488 19304 16540 19310
rect 16486 19272 16488 19281
rect 16540 19272 16542 19281
rect 16486 19207 16542 19216
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 16500 18970 16528 19110
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16500 18426 16528 18702
rect 16488 18420 16540 18426
rect 16488 18362 16540 18368
rect 16488 18216 16540 18222
rect 16488 18158 16540 18164
rect 16396 17876 16448 17882
rect 16396 17818 16448 17824
rect 16500 17785 16528 18158
rect 16486 17776 16542 17785
rect 16486 17711 16542 17720
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16500 17513 16528 17546
rect 16486 17504 16542 17513
rect 16486 17439 16542 17448
rect 16396 17128 16448 17134
rect 16396 17070 16448 17076
rect 16408 16833 16436 17070
rect 16488 17060 16540 17066
rect 16488 17002 16540 17008
rect 16394 16824 16450 16833
rect 16394 16759 16450 16768
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16408 13870 16436 14758
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 16408 11082 16436 12854
rect 16500 11150 16528 17002
rect 16592 15026 16620 19654
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16684 14890 16712 23480
rect 16776 20942 16804 26930
rect 16856 25220 16908 25226
rect 16856 25162 16908 25168
rect 16868 24614 16896 25162
rect 16948 25152 17000 25158
rect 16948 25094 17000 25100
rect 16856 24608 16908 24614
rect 16856 24550 16908 24556
rect 16868 24342 16896 24550
rect 16856 24336 16908 24342
rect 16856 24278 16908 24284
rect 16868 23118 16896 24278
rect 16960 24206 16988 25094
rect 16948 24200 17000 24206
rect 16948 24142 17000 24148
rect 16960 23526 16988 24142
rect 16948 23520 17000 23526
rect 16948 23462 17000 23468
rect 16856 23112 16908 23118
rect 16856 23054 16908 23060
rect 16868 21962 16896 23054
rect 16856 21956 16908 21962
rect 16856 21898 16908 21904
rect 16868 21146 16896 21898
rect 16856 21140 16908 21146
rect 16856 21082 16908 21088
rect 16764 20936 16816 20942
rect 16764 20878 16816 20884
rect 17052 20754 17080 27270
rect 16868 20726 17080 20754
rect 16764 20460 16816 20466
rect 16764 20402 16816 20408
rect 16776 19718 16804 20402
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16764 19372 16816 19378
rect 16764 19314 16816 19320
rect 16776 17338 16804 19314
rect 16764 17332 16816 17338
rect 16764 17274 16816 17280
rect 16762 17232 16818 17241
rect 16762 17167 16818 17176
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16578 14648 16634 14657
rect 16578 14583 16580 14592
rect 16632 14583 16634 14592
rect 16580 14554 16632 14560
rect 16670 14512 16726 14521
rect 16670 14447 16726 14456
rect 16684 14346 16712 14447
rect 16672 14340 16724 14346
rect 16672 14282 16724 14288
rect 16580 14000 16632 14006
rect 16580 13942 16632 13948
rect 16592 13530 16620 13942
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16684 12986 16712 13806
rect 16672 12980 16724 12986
rect 16672 12922 16724 12928
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16396 11076 16448 11082
rect 16396 11018 16448 11024
rect 16408 10810 16436 11018
rect 16488 11008 16540 11014
rect 16488 10950 16540 10956
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 16408 10266 16436 10610
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16500 10062 16528 10950
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16304 7812 16356 7818
rect 16304 7754 16356 7760
rect 16132 7500 16252 7528
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16132 3738 16160 7346
rect 16224 6390 16252 7500
rect 16304 7268 16356 7274
rect 16304 7210 16356 7216
rect 16212 6384 16264 6390
rect 16212 6326 16264 6332
rect 16212 5568 16264 5574
rect 16212 5510 16264 5516
rect 16224 4622 16252 5510
rect 16316 5166 16344 7210
rect 16408 7206 16436 9862
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16408 6322 16436 7142
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16408 5846 16436 6054
rect 16396 5840 16448 5846
rect 16396 5782 16448 5788
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16224 3942 16252 4014
rect 16408 3942 16436 4626
rect 16212 3936 16264 3942
rect 16212 3878 16264 3884
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16224 2774 16252 3878
rect 16500 3534 16528 9998
rect 16592 7478 16620 12786
rect 16684 12170 16712 12922
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 16684 11286 16712 12106
rect 16672 11280 16724 11286
rect 16672 11222 16724 11228
rect 16684 10674 16712 11222
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 16670 10160 16726 10169
rect 16670 10095 16726 10104
rect 16684 9654 16712 10095
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16580 7472 16632 7478
rect 16580 7414 16632 7420
rect 16684 6633 16712 9454
rect 16776 7562 16804 17167
rect 16868 17105 16896 20726
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 16854 17096 16910 17105
rect 16854 17031 16910 17040
rect 16856 16992 16908 16998
rect 16960 16969 16988 20538
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 17052 20058 17080 20402
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 17040 19848 17092 19854
rect 17040 19790 17092 19796
rect 17052 18737 17080 19790
rect 17038 18728 17094 18737
rect 17038 18663 17094 18672
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 16856 16934 16908 16940
rect 16946 16960 17002 16969
rect 16868 16114 16896 16934
rect 17052 16946 17080 18566
rect 17144 17241 17172 27338
rect 17224 24744 17276 24750
rect 17224 24686 17276 24692
rect 17236 24410 17264 24686
rect 17224 24404 17276 24410
rect 17224 24346 17276 24352
rect 17224 24268 17276 24274
rect 17224 24210 17276 24216
rect 17236 23730 17264 24210
rect 17224 23724 17276 23730
rect 17224 23666 17276 23672
rect 17224 21344 17276 21350
rect 17224 21286 17276 21292
rect 17236 20942 17264 21286
rect 17224 20936 17276 20942
rect 17224 20878 17276 20884
rect 17236 20398 17264 20878
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 17224 19304 17276 19310
rect 17224 19246 17276 19252
rect 17236 18737 17264 19246
rect 17222 18728 17278 18737
rect 17222 18663 17278 18672
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17236 18193 17264 18566
rect 17222 18184 17278 18193
rect 17222 18119 17278 18128
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17130 17232 17186 17241
rect 17130 17167 17186 17176
rect 17236 17134 17264 17818
rect 17328 17202 17356 28358
rect 17500 26376 17552 26382
rect 17500 26318 17552 26324
rect 17512 26042 17540 26318
rect 17500 26036 17552 26042
rect 17500 25978 17552 25984
rect 17408 25764 17460 25770
rect 17408 25706 17460 25712
rect 17420 20602 17448 25706
rect 17500 24812 17552 24818
rect 17500 24754 17552 24760
rect 17512 24138 17540 24754
rect 17500 24132 17552 24138
rect 17500 24074 17552 24080
rect 17604 22094 17632 28494
rect 18052 27872 18104 27878
rect 18052 27814 18104 27820
rect 17684 26988 17736 26994
rect 17684 26930 17736 26936
rect 17696 26382 17724 26930
rect 17960 26920 18012 26926
rect 17960 26862 18012 26868
rect 17972 26382 18000 26862
rect 17684 26376 17736 26382
rect 17684 26318 17736 26324
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 17696 26246 17724 26318
rect 17776 26308 17828 26314
rect 17776 26250 17828 26256
rect 17684 26240 17736 26246
rect 17684 26182 17736 26188
rect 17696 25906 17724 26182
rect 17684 25900 17736 25906
rect 17684 25842 17736 25848
rect 17696 24818 17724 25842
rect 17684 24812 17736 24818
rect 17684 24754 17736 24760
rect 17788 24410 17816 26250
rect 17972 25906 18000 26318
rect 18064 26314 18092 27814
rect 18156 27674 18184 28494
rect 18144 27668 18196 27674
rect 18144 27610 18196 27616
rect 18236 27600 18288 27606
rect 18236 27542 18288 27548
rect 18144 26784 18196 26790
rect 18144 26726 18196 26732
rect 18052 26308 18104 26314
rect 18052 26250 18104 26256
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 17868 25424 17920 25430
rect 17868 25366 17920 25372
rect 17776 24404 17828 24410
rect 17776 24346 17828 24352
rect 17684 24336 17736 24342
rect 17880 24290 17908 25366
rect 17972 25362 18000 25842
rect 18156 25838 18184 26726
rect 18144 25832 18196 25838
rect 18144 25774 18196 25780
rect 17960 25356 18012 25362
rect 17960 25298 18012 25304
rect 18248 24970 18276 27542
rect 17684 24278 17736 24284
rect 17696 22778 17724 24278
rect 17788 24262 17908 24290
rect 17972 24942 18276 24970
rect 17684 22772 17736 22778
rect 17684 22714 17736 22720
rect 17788 22094 17816 24262
rect 17868 23860 17920 23866
rect 17868 23802 17920 23808
rect 17880 22658 17908 23802
rect 17972 22778 18000 24942
rect 18236 24812 18288 24818
rect 18236 24754 18288 24760
rect 18248 24206 18276 24754
rect 18236 24200 18288 24206
rect 18236 24142 18288 24148
rect 18236 24064 18288 24070
rect 18236 24006 18288 24012
rect 18248 23526 18276 24006
rect 18052 23520 18104 23526
rect 18052 23462 18104 23468
rect 18236 23520 18288 23526
rect 18236 23462 18288 23468
rect 18064 23322 18092 23462
rect 18340 23338 18368 28630
rect 19248 28620 19300 28626
rect 19248 28562 19300 28568
rect 18696 28552 18748 28558
rect 18696 28494 18748 28500
rect 18604 28416 18656 28422
rect 18604 28358 18656 28364
rect 18616 28082 18644 28358
rect 18604 28076 18656 28082
rect 18604 28018 18656 28024
rect 18708 27538 18736 28494
rect 18920 28316 19228 28336
rect 18920 28314 18926 28316
rect 18982 28314 19006 28316
rect 19062 28314 19086 28316
rect 19142 28314 19166 28316
rect 19222 28314 19228 28316
rect 18982 28262 18984 28314
rect 19164 28262 19166 28314
rect 18920 28260 18926 28262
rect 18982 28260 19006 28262
rect 19062 28260 19086 28262
rect 19142 28260 19166 28262
rect 19222 28260 19228 28262
rect 18920 28240 19228 28260
rect 18696 27532 18748 27538
rect 18696 27474 18748 27480
rect 18512 27464 18564 27470
rect 18512 27406 18564 27412
rect 18524 27130 18552 27406
rect 18708 27146 18736 27474
rect 18920 27228 19228 27248
rect 18920 27226 18926 27228
rect 18982 27226 19006 27228
rect 19062 27226 19086 27228
rect 19142 27226 19166 27228
rect 19222 27226 19228 27228
rect 18982 27174 18984 27226
rect 19164 27174 19166 27226
rect 18920 27172 18926 27174
rect 18982 27172 19006 27174
rect 19062 27172 19086 27174
rect 19142 27172 19166 27174
rect 19222 27172 19228 27174
rect 18920 27152 19228 27172
rect 18512 27124 18564 27130
rect 18708 27118 18828 27146
rect 18512 27066 18564 27072
rect 18696 26988 18748 26994
rect 18696 26930 18748 26936
rect 18420 26308 18472 26314
rect 18420 26250 18472 26256
rect 18432 24070 18460 26250
rect 18708 26058 18736 26930
rect 18800 26450 18828 27118
rect 18788 26444 18840 26450
rect 18788 26386 18840 26392
rect 19260 26353 19288 28562
rect 19800 28552 19852 28558
rect 19800 28494 19852 28500
rect 19616 28416 19668 28422
rect 19616 28358 19668 28364
rect 19628 28082 19656 28358
rect 19708 28144 19760 28150
rect 19708 28086 19760 28092
rect 19616 28076 19668 28082
rect 19616 28018 19668 28024
rect 19432 27872 19484 27878
rect 19352 27832 19432 27860
rect 19352 27062 19380 27832
rect 19432 27814 19484 27820
rect 19340 27056 19392 27062
rect 19340 26998 19392 27004
rect 19246 26344 19302 26353
rect 19246 26279 19302 26288
rect 19248 26240 19300 26246
rect 19352 26217 19380 26998
rect 19616 26920 19668 26926
rect 19616 26862 19668 26868
rect 19628 26382 19656 26862
rect 19432 26376 19484 26382
rect 19616 26376 19668 26382
rect 19484 26336 19564 26364
rect 19432 26318 19484 26324
rect 19536 26217 19564 26336
rect 19616 26318 19668 26324
rect 19248 26182 19300 26188
rect 19338 26208 19394 26217
rect 18920 26140 19228 26160
rect 18920 26138 18926 26140
rect 18982 26138 19006 26140
rect 19062 26138 19086 26140
rect 19142 26138 19166 26140
rect 19222 26138 19228 26140
rect 18982 26086 18984 26138
rect 19164 26086 19166 26138
rect 18920 26084 18926 26086
rect 18982 26084 19006 26086
rect 19062 26084 19086 26086
rect 19142 26084 19166 26086
rect 19222 26084 19228 26086
rect 18920 26064 19228 26084
rect 18708 26030 18828 26058
rect 18696 25968 18748 25974
rect 18696 25910 18748 25916
rect 18604 25832 18656 25838
rect 18604 25774 18656 25780
rect 18512 25764 18564 25770
rect 18512 25706 18564 25712
rect 18420 24064 18472 24070
rect 18420 24006 18472 24012
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 18156 23310 18368 23338
rect 17960 22772 18012 22778
rect 17960 22714 18012 22720
rect 17880 22642 18000 22658
rect 17880 22636 18012 22642
rect 17880 22630 17960 22636
rect 17960 22578 18012 22584
rect 17512 22066 17632 22094
rect 17696 22066 17816 22094
rect 17868 22092 17920 22098
rect 17408 20596 17460 20602
rect 17408 20538 17460 20544
rect 17408 19372 17460 19378
rect 17408 19314 17460 19320
rect 17420 18766 17448 19314
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 17420 18057 17448 18362
rect 17406 18048 17462 18057
rect 17406 17983 17462 17992
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 17224 17128 17276 17134
rect 17224 17070 17276 17076
rect 17316 16992 17368 16998
rect 17052 16918 17172 16946
rect 17316 16934 17368 16940
rect 16946 16895 17002 16904
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16868 15026 16896 15846
rect 16960 15706 16988 16526
rect 17144 16046 17172 16918
rect 17328 16794 17356 16934
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17224 16720 17276 16726
rect 17224 16662 17276 16668
rect 17236 16153 17264 16662
rect 17420 16454 17448 17983
rect 17408 16448 17460 16454
rect 17408 16390 17460 16396
rect 17222 16144 17278 16153
rect 17222 16079 17278 16088
rect 17132 16040 17184 16046
rect 17184 16000 17264 16028
rect 17132 15982 17184 15988
rect 16948 15700 17000 15706
rect 16948 15642 17000 15648
rect 16948 15360 17000 15366
rect 16948 15302 17000 15308
rect 17130 15328 17186 15337
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16856 14884 16908 14890
rect 16856 14826 16908 14832
rect 16868 13172 16896 14826
rect 16960 13326 16988 15302
rect 17130 15263 17186 15272
rect 17144 13512 17172 15263
rect 17236 14414 17264 16000
rect 17408 15020 17460 15026
rect 17408 14962 17460 14968
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17144 13484 17264 13512
rect 17130 13424 17186 13433
rect 17130 13359 17186 13368
rect 17144 13326 17172 13359
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 16868 13144 16988 13172
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16868 8514 16896 12582
rect 16960 12322 16988 13144
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 16960 12294 17080 12322
rect 16946 12200 17002 12209
rect 16946 12135 17002 12144
rect 16960 9518 16988 12135
rect 17052 9722 17080 12294
rect 17040 9716 17092 9722
rect 17040 9658 17092 9664
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16960 8974 16988 9318
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 17052 8634 17080 9522
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 16868 8486 17080 8514
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 16868 8294 16896 8325
rect 16856 8288 16908 8294
rect 16960 8242 16988 8366
rect 16908 8236 16988 8242
rect 16856 8230 16988 8236
rect 16868 8214 16988 8230
rect 16868 7721 16896 8214
rect 16948 7744 17000 7750
rect 16854 7712 16910 7721
rect 16948 7686 17000 7692
rect 16854 7647 16910 7656
rect 16776 7534 16896 7562
rect 16762 7440 16818 7449
rect 16762 7375 16764 7384
rect 16816 7375 16818 7384
rect 16764 7346 16816 7352
rect 16764 7268 16816 7274
rect 16764 7210 16816 7216
rect 16670 6624 16726 6633
rect 16670 6559 16726 6568
rect 16684 6458 16712 6559
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 16776 6338 16804 7210
rect 16684 6310 16804 6338
rect 16684 4554 16712 6310
rect 16762 6216 16818 6225
rect 16762 6151 16818 6160
rect 16776 5710 16804 6151
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 16672 4548 16724 4554
rect 16672 4490 16724 4496
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 16500 3058 16528 3334
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16592 2774 16620 4422
rect 16776 4146 16804 5510
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16672 3120 16724 3126
rect 16672 3062 16724 3068
rect 16132 2746 16252 2774
rect 16316 2746 16620 2774
rect 16132 2446 16160 2746
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 16316 800 16344 2746
rect 16684 2666 16712 3062
rect 16868 2774 16896 7534
rect 16960 7410 16988 7686
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16946 7304 17002 7313
rect 16946 7239 17002 7248
rect 16960 3194 16988 7239
rect 17052 5710 17080 8486
rect 17040 5704 17092 5710
rect 17040 5646 17092 5652
rect 17038 5536 17094 5545
rect 17038 5471 17094 5480
rect 17052 3670 17080 5471
rect 17144 4826 17172 12786
rect 17236 11354 17264 13484
rect 17316 12708 17368 12714
rect 17316 12650 17368 12656
rect 17328 11898 17356 12650
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17314 11656 17370 11665
rect 17314 11591 17370 11600
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 17328 11234 17356 11591
rect 17236 11206 17356 11234
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 17040 3664 17092 3670
rect 17040 3606 17092 3612
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 16868 2746 17080 2774
rect 16592 2638 16712 2666
rect 16592 800 16620 2638
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 16776 2106 16804 2246
rect 16764 2100 16816 2106
rect 16764 2042 16816 2048
rect 16868 2038 16896 2246
rect 16856 2032 16908 2038
rect 16856 1974 16908 1980
rect 16764 1964 16816 1970
rect 16764 1906 16816 1912
rect 16776 800 16804 1906
rect 17052 800 17080 2746
rect 17144 1970 17172 3606
rect 17236 3058 17264 11206
rect 17314 11112 17370 11121
rect 17314 11047 17370 11056
rect 17328 10810 17356 11047
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17328 9178 17356 9998
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17316 8832 17368 8838
rect 17316 8774 17368 8780
rect 17328 7954 17356 8774
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17328 6798 17356 7890
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17328 5778 17356 6734
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 17328 5302 17356 5714
rect 17316 5296 17368 5302
rect 17316 5238 17368 5244
rect 17328 4690 17356 5238
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17420 3534 17448 14962
rect 17512 12186 17540 22066
rect 17592 20800 17644 20806
rect 17592 20742 17644 20748
rect 17604 18193 17632 20742
rect 17696 19718 17724 22066
rect 17868 22034 17920 22040
rect 17880 21486 17908 22034
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 17972 21554 18000 21966
rect 18052 21888 18104 21894
rect 18052 21830 18104 21836
rect 18064 21554 18092 21830
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 17868 21480 17920 21486
rect 17868 21422 17920 21428
rect 18064 20942 18092 21490
rect 18052 20936 18104 20942
rect 18052 20878 18104 20884
rect 17868 20800 17920 20806
rect 17868 20742 17920 20748
rect 17880 20534 17908 20742
rect 17868 20528 17920 20534
rect 17774 20496 17830 20505
rect 17868 20470 17920 20476
rect 17960 20528 18012 20534
rect 17960 20470 18012 20476
rect 17774 20431 17830 20440
rect 17684 19712 17736 19718
rect 17684 19654 17736 19660
rect 17684 19508 17736 19514
rect 17684 19450 17736 19456
rect 17590 18184 17646 18193
rect 17590 18119 17646 18128
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17604 17338 17632 17546
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17696 17218 17724 19450
rect 17788 19360 17816 20431
rect 17868 19372 17920 19378
rect 17788 19332 17868 19360
rect 17868 19314 17920 19320
rect 17880 19242 17908 19314
rect 17868 19236 17920 19242
rect 17868 19178 17920 19184
rect 17880 18766 17908 19178
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17868 18760 17920 18766
rect 17868 18702 17920 18708
rect 17788 18290 17816 18702
rect 17776 18284 17828 18290
rect 17776 18226 17828 18232
rect 17880 18222 17908 18702
rect 17868 18216 17920 18222
rect 17868 18158 17920 18164
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17880 17921 17908 18022
rect 17866 17912 17922 17921
rect 17866 17847 17922 17856
rect 17972 17762 18000 20470
rect 18052 20460 18104 20466
rect 18052 20402 18104 20408
rect 18064 20058 18092 20402
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 18052 19916 18104 19922
rect 18052 19858 18104 19864
rect 17880 17734 18000 17762
rect 17776 17536 17828 17542
rect 17776 17478 17828 17484
rect 17604 17190 17724 17218
rect 17604 15065 17632 17190
rect 17684 17128 17736 17134
rect 17684 17070 17736 17076
rect 17590 15056 17646 15065
rect 17590 14991 17646 15000
rect 17592 14544 17644 14550
rect 17592 14486 17644 14492
rect 17604 13705 17632 14486
rect 17590 13696 17646 13705
rect 17590 13631 17646 13640
rect 17592 13524 17644 13530
rect 17592 13466 17644 13472
rect 17604 12345 17632 13466
rect 17590 12336 17646 12345
rect 17590 12271 17646 12280
rect 17512 12158 17632 12186
rect 17604 12073 17632 12158
rect 17696 12102 17724 17070
rect 17788 17066 17816 17478
rect 17776 17060 17828 17066
rect 17776 17002 17828 17008
rect 17788 16590 17816 17002
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17880 16454 17908 17734
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 17868 16448 17920 16454
rect 17868 16390 17920 16396
rect 17788 16266 17816 16390
rect 17788 16238 17908 16266
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17788 15706 17816 16050
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17880 15586 17908 16238
rect 17972 16114 18000 17614
rect 18064 16998 18092 19858
rect 18156 18034 18184 23310
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 18248 22030 18276 22578
rect 18340 22166 18368 23054
rect 18328 22160 18380 22166
rect 18328 22102 18380 22108
rect 18236 22024 18288 22030
rect 18236 21966 18288 21972
rect 18234 21856 18290 21865
rect 18234 21791 18290 21800
rect 18248 18465 18276 21791
rect 18328 21072 18380 21078
rect 18328 21014 18380 21020
rect 18340 19961 18368 21014
rect 18326 19952 18382 19961
rect 18326 19887 18382 19896
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 18340 19514 18368 19790
rect 18328 19508 18380 19514
rect 18328 19450 18380 19456
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 18340 19174 18368 19246
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18340 18902 18368 19110
rect 18328 18896 18380 18902
rect 18328 18838 18380 18844
rect 18234 18456 18290 18465
rect 18234 18391 18290 18400
rect 18340 18290 18368 18838
rect 18432 18766 18460 24006
rect 18524 23798 18552 25706
rect 18616 24886 18644 25774
rect 18708 24954 18736 25910
rect 18696 24948 18748 24954
rect 18696 24890 18748 24896
rect 18604 24880 18656 24886
rect 18604 24822 18656 24828
rect 18512 23792 18564 23798
rect 18512 23734 18564 23740
rect 18512 23656 18564 23662
rect 18512 23598 18564 23604
rect 18524 23118 18552 23598
rect 18512 23112 18564 23118
rect 18512 23054 18564 23060
rect 18616 23066 18644 24822
rect 18800 24410 18828 26030
rect 19260 25906 19288 26182
rect 19338 26143 19394 26152
rect 19522 26208 19578 26217
rect 19522 26143 19578 26152
rect 19340 26036 19392 26042
rect 19720 26024 19748 28086
rect 19812 26586 19840 28494
rect 19892 27464 19944 27470
rect 19892 27406 19944 27412
rect 19904 26994 19932 27406
rect 20076 27328 20128 27334
rect 20076 27270 20128 27276
rect 19892 26988 19944 26994
rect 19892 26930 19944 26936
rect 19800 26580 19852 26586
rect 19800 26522 19852 26528
rect 19800 26376 19852 26382
rect 19800 26318 19852 26324
rect 19392 25996 19748 26024
rect 19340 25978 19392 25984
rect 19338 25936 19394 25945
rect 19248 25900 19300 25906
rect 19338 25871 19394 25880
rect 19522 25936 19578 25945
rect 19522 25871 19578 25880
rect 19248 25842 19300 25848
rect 18920 25052 19228 25072
rect 18920 25050 18926 25052
rect 18982 25050 19006 25052
rect 19062 25050 19086 25052
rect 19142 25050 19166 25052
rect 19222 25050 19228 25052
rect 18982 24998 18984 25050
rect 19164 24998 19166 25050
rect 18920 24996 18926 24998
rect 18982 24996 19006 24998
rect 19062 24996 19086 24998
rect 19142 24996 19166 24998
rect 19222 24996 19228 24998
rect 18920 24976 19228 24996
rect 19248 24744 19300 24750
rect 19248 24686 19300 24692
rect 18788 24404 18840 24410
rect 18788 24346 18840 24352
rect 18920 23964 19228 23984
rect 18920 23962 18926 23964
rect 18982 23962 19006 23964
rect 19062 23962 19086 23964
rect 19142 23962 19166 23964
rect 19222 23962 19228 23964
rect 18982 23910 18984 23962
rect 19164 23910 19166 23962
rect 18920 23908 18926 23910
rect 18982 23908 19006 23910
rect 19062 23908 19086 23910
rect 19142 23908 19166 23910
rect 19222 23908 19228 23910
rect 18920 23888 19228 23908
rect 19260 23866 19288 24686
rect 19352 24070 19380 25871
rect 19536 24954 19564 25871
rect 19616 25832 19668 25838
rect 19616 25774 19668 25780
rect 19628 25498 19656 25774
rect 19616 25492 19668 25498
rect 19616 25434 19668 25440
rect 19524 24948 19576 24954
rect 19524 24890 19576 24896
rect 19430 24848 19486 24857
rect 19430 24783 19486 24792
rect 19444 24614 19472 24783
rect 19432 24608 19484 24614
rect 19432 24550 19484 24556
rect 19432 24404 19484 24410
rect 19432 24346 19484 24352
rect 19340 24064 19392 24070
rect 19340 24006 19392 24012
rect 19248 23860 19300 23866
rect 19248 23802 19300 23808
rect 19156 23792 19208 23798
rect 19156 23734 19208 23740
rect 18696 23656 18748 23662
rect 18696 23598 18748 23604
rect 18708 23186 18736 23598
rect 18696 23180 18748 23186
rect 18696 23122 18748 23128
rect 18616 23038 18736 23066
rect 19168 23050 19196 23734
rect 19248 23656 19300 23662
rect 19248 23598 19300 23604
rect 18512 22772 18564 22778
rect 18512 22714 18564 22720
rect 18604 22772 18656 22778
rect 18604 22714 18656 22720
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18524 18578 18552 22714
rect 18616 20534 18644 22714
rect 18604 20528 18656 20534
rect 18604 20470 18656 20476
rect 18708 20380 18736 23038
rect 19156 23044 19208 23050
rect 19156 22986 19208 22992
rect 18920 22876 19228 22896
rect 18920 22874 18926 22876
rect 18982 22874 19006 22876
rect 19062 22874 19086 22876
rect 19142 22874 19166 22876
rect 19222 22874 19228 22876
rect 18982 22822 18984 22874
rect 19164 22822 19166 22874
rect 18920 22820 18926 22822
rect 18982 22820 19006 22822
rect 19062 22820 19086 22822
rect 19142 22820 19166 22822
rect 19222 22820 19228 22822
rect 18920 22800 19228 22820
rect 18972 22432 19024 22438
rect 18972 22374 19024 22380
rect 18984 22234 19012 22374
rect 18972 22228 19024 22234
rect 18972 22170 19024 22176
rect 18920 21788 19228 21808
rect 18920 21786 18926 21788
rect 18982 21786 19006 21788
rect 19062 21786 19086 21788
rect 19142 21786 19166 21788
rect 19222 21786 19228 21788
rect 18982 21734 18984 21786
rect 19164 21734 19166 21786
rect 18920 21732 18926 21734
rect 18982 21732 19006 21734
rect 19062 21732 19086 21734
rect 19142 21732 19166 21734
rect 19222 21732 19228 21734
rect 18920 21712 19228 21732
rect 18788 21616 18840 21622
rect 18788 21558 18840 21564
rect 18432 18550 18552 18578
rect 18616 20352 18736 20380
rect 18328 18284 18380 18290
rect 18328 18226 18380 18232
rect 18156 18006 18368 18034
rect 18142 17912 18198 17921
rect 18142 17847 18198 17856
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 18052 16720 18104 16726
rect 18052 16662 18104 16668
rect 18064 16114 18092 16662
rect 18156 16590 18184 17847
rect 18234 17096 18290 17105
rect 18234 17031 18290 17040
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 17788 15558 17908 15586
rect 17788 14278 17816 15558
rect 17972 15502 18000 16050
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17972 15026 18000 15438
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17880 14550 17908 14894
rect 17868 14544 17920 14550
rect 17868 14486 17920 14492
rect 18052 14544 18104 14550
rect 18052 14486 18104 14492
rect 17880 14414 17908 14486
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17776 14272 17828 14278
rect 17776 14214 17828 14220
rect 17868 13796 17920 13802
rect 17868 13738 17920 13744
rect 17776 13728 17828 13734
rect 17776 13670 17828 13676
rect 17788 13326 17816 13670
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17880 13190 17908 13738
rect 17960 13728 18012 13734
rect 17960 13670 18012 13676
rect 17972 13258 18000 13670
rect 18064 13297 18092 14486
rect 18050 13288 18106 13297
rect 17960 13252 18012 13258
rect 18050 13223 18106 13232
rect 17960 13194 18012 13200
rect 17868 13184 17920 13190
rect 17774 13152 17830 13161
rect 17868 13126 17920 13132
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 17774 13087 17830 13096
rect 17788 12170 17816 13087
rect 17958 13016 18014 13025
rect 17868 12980 17920 12986
rect 17958 12951 18014 12960
rect 17868 12922 17920 12928
rect 17880 12889 17908 12922
rect 17866 12880 17922 12889
rect 17866 12815 17922 12824
rect 17776 12164 17828 12170
rect 17776 12106 17828 12112
rect 17684 12096 17736 12102
rect 17590 12064 17646 12073
rect 17684 12038 17736 12044
rect 17590 11999 17646 12008
rect 17590 11928 17646 11937
rect 17500 11892 17552 11898
rect 17590 11863 17646 11872
rect 17500 11834 17552 11840
rect 17512 6798 17540 11834
rect 17604 10062 17632 11863
rect 17682 11792 17738 11801
rect 17788 11762 17816 12106
rect 17682 11727 17738 11736
rect 17776 11756 17828 11762
rect 17696 10062 17724 11727
rect 17776 11698 17828 11704
rect 17866 10840 17922 10849
rect 17866 10775 17922 10784
rect 17880 10606 17908 10775
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17592 10056 17644 10062
rect 17592 9998 17644 10004
rect 17684 10056 17736 10062
rect 17868 10056 17920 10062
rect 17684 9998 17736 10004
rect 17774 10024 17830 10033
rect 17868 9998 17920 10004
rect 17774 9959 17830 9968
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17604 7886 17632 9862
rect 17788 9722 17816 9959
rect 17684 9716 17736 9722
rect 17684 9658 17736 9664
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17696 8378 17724 9658
rect 17788 9450 17816 9658
rect 17776 9444 17828 9450
rect 17776 9386 17828 9392
rect 17776 8832 17828 8838
rect 17776 8774 17828 8780
rect 17788 8566 17816 8774
rect 17776 8560 17828 8566
rect 17776 8502 17828 8508
rect 17696 8350 17816 8378
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17604 6458 17632 7346
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 17604 6202 17632 6258
rect 17512 6174 17632 6202
rect 17512 3738 17540 6174
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17604 5574 17632 6054
rect 17592 5568 17644 5574
rect 17592 5510 17644 5516
rect 17592 4820 17644 4826
rect 17592 4762 17644 4768
rect 17604 4214 17632 4762
rect 17592 4208 17644 4214
rect 17592 4150 17644 4156
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 17696 2774 17724 7686
rect 17604 2746 17724 2774
rect 17788 2774 17816 8350
rect 17880 7546 17908 9998
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17868 7268 17920 7274
rect 17868 7210 17920 7216
rect 17880 6769 17908 7210
rect 17866 6760 17922 6769
rect 17866 6695 17922 6704
rect 17868 6656 17920 6662
rect 17866 6624 17868 6633
rect 17920 6624 17922 6633
rect 17866 6559 17922 6568
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 17880 6361 17908 6394
rect 17972 6390 18000 12951
rect 18064 12442 18092 13126
rect 18156 12918 18184 16390
rect 18144 12912 18196 12918
rect 18144 12854 18196 12860
rect 18248 12764 18276 17031
rect 18340 13025 18368 18006
rect 18432 17082 18460 18550
rect 18510 18456 18566 18465
rect 18616 18426 18644 20352
rect 18696 20052 18748 20058
rect 18696 19994 18748 20000
rect 18708 19378 18736 19994
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18800 19281 18828 21558
rect 18972 21344 19024 21350
rect 18972 21286 19024 21292
rect 18984 21146 19012 21286
rect 18972 21140 19024 21146
rect 18972 21082 19024 21088
rect 18920 20700 19228 20720
rect 18920 20698 18926 20700
rect 18982 20698 19006 20700
rect 19062 20698 19086 20700
rect 19142 20698 19166 20700
rect 19222 20698 19228 20700
rect 18982 20646 18984 20698
rect 19164 20646 19166 20698
rect 18920 20644 18926 20646
rect 18982 20644 19006 20646
rect 19062 20644 19086 20646
rect 19142 20644 19166 20646
rect 19222 20644 19228 20646
rect 18920 20624 19228 20644
rect 19156 20256 19208 20262
rect 19156 20198 19208 20204
rect 19168 19854 19196 20198
rect 19156 19848 19208 19854
rect 19154 19816 19156 19825
rect 19208 19816 19210 19825
rect 19154 19751 19210 19760
rect 18920 19612 19228 19632
rect 18920 19610 18926 19612
rect 18982 19610 19006 19612
rect 19062 19610 19086 19612
rect 19142 19610 19166 19612
rect 19222 19610 19228 19612
rect 18982 19558 18984 19610
rect 19164 19558 19166 19610
rect 18920 19556 18926 19558
rect 18982 19556 19006 19558
rect 19062 19556 19086 19558
rect 19142 19556 19166 19558
rect 19222 19556 19228 19558
rect 18920 19536 19228 19556
rect 18970 19408 19026 19417
rect 18880 19372 18932 19378
rect 18970 19343 19026 19352
rect 18880 19314 18932 19320
rect 18786 19272 18842 19281
rect 18708 19230 18786 19258
rect 18510 18391 18566 18400
rect 18604 18420 18656 18426
rect 18524 17202 18552 18391
rect 18604 18362 18656 18368
rect 18602 18184 18658 18193
rect 18602 18119 18658 18128
rect 18512 17196 18564 17202
rect 18512 17138 18564 17144
rect 18432 17054 18552 17082
rect 18418 16960 18474 16969
rect 18524 16946 18552 17054
rect 18616 17048 18644 18119
rect 18708 17202 18736 19230
rect 18786 19207 18842 19216
rect 18892 19145 18920 19314
rect 18878 19136 18934 19145
rect 18878 19071 18934 19080
rect 18984 19009 19012 19343
rect 19260 19334 19288 23598
rect 19352 20058 19380 24006
rect 19444 22778 19472 24346
rect 19522 24304 19578 24313
rect 19522 24239 19578 24248
rect 19616 24268 19668 24274
rect 19536 24206 19564 24239
rect 19616 24210 19668 24216
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19522 23760 19578 23769
rect 19522 23695 19524 23704
rect 19576 23695 19578 23704
rect 19524 23666 19576 23672
rect 19524 23588 19576 23594
rect 19524 23530 19576 23536
rect 19536 23118 19564 23530
rect 19524 23112 19576 23118
rect 19524 23054 19576 23060
rect 19628 22982 19656 24210
rect 19720 23882 19748 25996
rect 19812 25906 19840 26318
rect 20088 26314 20116 27270
rect 20076 26308 20128 26314
rect 20076 26250 20128 26256
rect 19800 25900 19852 25906
rect 19800 25842 19852 25848
rect 19984 25900 20036 25906
rect 19984 25842 20036 25848
rect 19800 25696 19852 25702
rect 19800 25638 19852 25644
rect 19812 24274 19840 25638
rect 19892 25288 19944 25294
rect 19892 25230 19944 25236
rect 19800 24268 19852 24274
rect 19800 24210 19852 24216
rect 19720 23854 19840 23882
rect 19708 23724 19760 23730
rect 19708 23666 19760 23672
rect 19720 23050 19748 23666
rect 19708 23044 19760 23050
rect 19708 22986 19760 22992
rect 19616 22976 19668 22982
rect 19522 22944 19578 22953
rect 19616 22918 19668 22924
rect 19522 22879 19578 22888
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 19444 21350 19472 22578
rect 19536 22506 19564 22879
rect 19720 22794 19748 22986
rect 19628 22766 19748 22794
rect 19812 22778 19840 23854
rect 19904 23730 19932 25230
rect 19892 23724 19944 23730
rect 19892 23666 19944 23672
rect 19892 23180 19944 23186
rect 19892 23122 19944 23128
rect 19800 22772 19852 22778
rect 19524 22500 19576 22506
rect 19524 22442 19576 22448
rect 19522 22264 19578 22273
rect 19628 22234 19656 22766
rect 19800 22714 19852 22720
rect 19708 22704 19760 22710
rect 19708 22646 19760 22652
rect 19522 22199 19578 22208
rect 19616 22228 19668 22234
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19432 20868 19484 20874
rect 19432 20810 19484 20816
rect 19444 20262 19472 20810
rect 19536 20466 19564 22199
rect 19616 22170 19668 22176
rect 19628 21962 19656 22170
rect 19616 21956 19668 21962
rect 19616 21898 19668 21904
rect 19628 21486 19656 21898
rect 19720 21593 19748 22646
rect 19800 22568 19852 22574
rect 19800 22510 19852 22516
rect 19812 21729 19840 22510
rect 19904 22094 19932 23122
rect 19996 22273 20024 25842
rect 20088 24818 20116 26250
rect 20180 25242 20208 28630
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 21640 28552 21692 28558
rect 21640 28494 21692 28500
rect 20352 27872 20404 27878
rect 20352 27814 20404 27820
rect 20364 27402 20392 27814
rect 20352 27396 20404 27402
rect 20352 27338 20404 27344
rect 20352 27056 20404 27062
rect 20352 26998 20404 27004
rect 20364 25362 20392 26998
rect 20536 26444 20588 26450
rect 20536 26386 20588 26392
rect 20444 26376 20496 26382
rect 20444 26318 20496 26324
rect 20456 26042 20484 26318
rect 20444 26036 20496 26042
rect 20444 25978 20496 25984
rect 20548 25702 20576 26386
rect 20640 26228 20668 28494
rect 20720 28416 20772 28422
rect 20720 28358 20772 28364
rect 20732 26353 20760 28358
rect 20996 27872 21048 27878
rect 20996 27814 21048 27820
rect 20812 26784 20864 26790
rect 20812 26726 20864 26732
rect 20718 26344 20774 26353
rect 20718 26279 20774 26288
rect 20640 26200 20760 26228
rect 20626 26072 20682 26081
rect 20626 26007 20682 26016
rect 20640 25906 20668 26007
rect 20628 25900 20680 25906
rect 20628 25842 20680 25848
rect 20536 25696 20588 25702
rect 20536 25638 20588 25644
rect 20352 25356 20404 25362
rect 20352 25298 20404 25304
rect 20180 25214 20300 25242
rect 20168 25152 20220 25158
rect 20168 25094 20220 25100
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 19982 22264 20038 22273
rect 19982 22199 20038 22208
rect 19904 22066 20024 22094
rect 19892 22024 19944 22030
rect 19892 21966 19944 21972
rect 19798 21720 19854 21729
rect 19904 21690 19932 21966
rect 19798 21655 19854 21664
rect 19892 21684 19944 21690
rect 19892 21626 19944 21632
rect 19706 21584 19762 21593
rect 19706 21519 19762 21528
rect 19890 21584 19946 21593
rect 19890 21519 19946 21528
rect 19904 21486 19932 21519
rect 19616 21480 19668 21486
rect 19616 21422 19668 21428
rect 19892 21480 19944 21486
rect 19892 21422 19944 21428
rect 19892 21072 19944 21078
rect 19892 21014 19944 21020
rect 19616 20936 19668 20942
rect 19616 20878 19668 20884
rect 19524 20460 19576 20466
rect 19524 20402 19576 20408
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19168 19306 19288 19334
rect 19064 19236 19116 19242
rect 19168 19224 19196 19306
rect 19168 19196 19288 19224
rect 19064 19178 19116 19184
rect 18970 19000 19026 19009
rect 18970 18935 19026 18944
rect 18880 18896 18932 18902
rect 19076 18873 19104 19178
rect 18880 18838 18932 18844
rect 19062 18864 19118 18873
rect 18788 18760 18840 18766
rect 18892 18737 18920 18838
rect 19062 18799 19118 18808
rect 18788 18702 18840 18708
rect 18878 18728 18934 18737
rect 18800 17678 18828 18702
rect 18878 18663 18934 18672
rect 18920 18524 19228 18544
rect 18920 18522 18926 18524
rect 18982 18522 19006 18524
rect 19062 18522 19086 18524
rect 19142 18522 19166 18524
rect 19222 18522 19228 18524
rect 18982 18470 18984 18522
rect 19164 18470 19166 18522
rect 18920 18468 18926 18470
rect 18982 18468 19006 18470
rect 19062 18468 19086 18470
rect 19142 18468 19166 18470
rect 19222 18468 19228 18470
rect 18920 18448 19228 18468
rect 18880 18352 18932 18358
rect 18878 18320 18880 18329
rect 18932 18320 18934 18329
rect 18878 18255 18934 18264
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 18880 18216 18932 18222
rect 18880 18158 18932 18164
rect 18892 17746 18920 18158
rect 18984 18057 19012 18226
rect 18970 18048 19026 18057
rect 18970 17983 19026 17992
rect 19064 17808 19116 17814
rect 19062 17776 19064 17785
rect 19116 17776 19118 17785
rect 18880 17740 18932 17746
rect 19062 17711 19118 17720
rect 18880 17682 18932 17688
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18800 17270 18828 17614
rect 18920 17436 19228 17456
rect 18920 17434 18926 17436
rect 18982 17434 19006 17436
rect 19062 17434 19086 17436
rect 19142 17434 19166 17436
rect 19222 17434 19228 17436
rect 18982 17382 18984 17434
rect 19164 17382 19166 17434
rect 18920 17380 18926 17382
rect 18982 17380 19006 17382
rect 19062 17380 19086 17382
rect 19142 17380 19166 17382
rect 19222 17380 19228 17382
rect 18920 17360 19228 17380
rect 18788 17264 18840 17270
rect 18788 17206 18840 17212
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18972 17060 19024 17066
rect 18616 17020 18736 17048
rect 18524 16918 18644 16946
rect 18418 16895 18474 16904
rect 18432 14278 18460 16895
rect 18510 16824 18566 16833
rect 18510 16759 18566 16768
rect 18524 16726 18552 16759
rect 18512 16720 18564 16726
rect 18512 16662 18564 16668
rect 18512 16584 18564 16590
rect 18510 16552 18512 16561
rect 18564 16552 18566 16561
rect 18510 16487 18566 16496
rect 18510 14376 18566 14385
rect 18510 14311 18566 14320
rect 18524 14278 18552 14311
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18512 14068 18564 14074
rect 18512 14010 18564 14016
rect 18418 13968 18474 13977
rect 18524 13938 18552 14010
rect 18418 13903 18420 13912
rect 18472 13903 18474 13912
rect 18512 13932 18564 13938
rect 18420 13874 18472 13880
rect 18512 13874 18564 13880
rect 18420 13184 18472 13190
rect 18512 13184 18564 13190
rect 18420 13126 18472 13132
rect 18510 13152 18512 13161
rect 18564 13152 18566 13161
rect 18326 13016 18382 13025
rect 18432 12986 18460 13126
rect 18510 13087 18566 13096
rect 18510 13016 18566 13025
rect 18326 12951 18382 12960
rect 18420 12980 18472 12986
rect 18510 12951 18566 12960
rect 18420 12922 18472 12928
rect 18328 12912 18380 12918
rect 18328 12854 18380 12860
rect 18156 12736 18276 12764
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 18064 11121 18092 12242
rect 18050 11112 18106 11121
rect 18050 11047 18106 11056
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 18064 10538 18092 10950
rect 18052 10532 18104 10538
rect 18052 10474 18104 10480
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 17960 6384 18012 6390
rect 17866 6352 17922 6361
rect 17960 6326 18012 6332
rect 17866 6287 17922 6296
rect 17958 6080 18014 6089
rect 17958 6015 18014 6024
rect 17972 4570 18000 6015
rect 18064 5302 18092 9318
rect 18156 7750 18184 12736
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 18248 10266 18276 10950
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 18248 6769 18276 9522
rect 18234 6760 18290 6769
rect 18234 6695 18290 6704
rect 18142 6352 18198 6361
rect 18142 6287 18198 6296
rect 18052 5296 18104 5302
rect 18052 5238 18104 5244
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 17880 4542 18000 4570
rect 17880 3482 17908 4542
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17972 3670 18000 4422
rect 18064 4078 18092 5102
rect 18156 4146 18184 6287
rect 18236 6180 18288 6186
rect 18236 6122 18288 6128
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 17960 3664 18012 3670
rect 17960 3606 18012 3612
rect 18144 3596 18196 3602
rect 18144 3538 18196 3544
rect 17880 3454 18000 3482
rect 17972 3398 18000 3454
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 18156 3194 18184 3538
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 18156 2990 18184 3130
rect 18144 2984 18196 2990
rect 18144 2926 18196 2932
rect 17788 2746 18184 2774
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 17132 1964 17184 1970
rect 17132 1906 17184 1912
rect 17328 800 17356 2246
rect 17604 800 17632 2746
rect 17868 2304 17920 2310
rect 17868 2246 17920 2252
rect 17880 800 17908 2246
rect 18156 800 18184 2746
rect 18248 2378 18276 6122
rect 18340 2774 18368 12854
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18432 10266 18460 12786
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18432 8634 18460 10202
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18432 5234 18460 6258
rect 18420 5228 18472 5234
rect 18420 5170 18472 5176
rect 18420 5024 18472 5030
rect 18420 4966 18472 4972
rect 18432 3194 18460 4966
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 18524 3040 18552 12951
rect 18616 12322 18644 16918
rect 18708 15026 18736 17020
rect 18972 17002 19024 17008
rect 18984 16697 19012 17002
rect 18970 16688 19026 16697
rect 18970 16623 19026 16632
rect 18788 16516 18840 16522
rect 18788 16458 18840 16464
rect 18696 15020 18748 15026
rect 18696 14962 18748 14968
rect 18800 14618 18828 16458
rect 18920 16348 19228 16368
rect 18920 16346 18926 16348
rect 18982 16346 19006 16348
rect 19062 16346 19086 16348
rect 19142 16346 19166 16348
rect 19222 16346 19228 16348
rect 18982 16294 18984 16346
rect 19164 16294 19166 16346
rect 18920 16292 18926 16294
rect 18982 16292 19006 16294
rect 19062 16292 19086 16294
rect 19142 16292 19166 16294
rect 19222 16292 19228 16294
rect 18920 16272 19228 16292
rect 18920 15260 19228 15280
rect 18920 15258 18926 15260
rect 18982 15258 19006 15260
rect 19062 15258 19086 15260
rect 19142 15258 19166 15260
rect 19222 15258 19228 15260
rect 18982 15206 18984 15258
rect 19164 15206 19166 15258
rect 18920 15204 18926 15206
rect 18982 15204 19006 15206
rect 19062 15204 19086 15206
rect 19142 15204 19166 15206
rect 19222 15204 19228 15206
rect 18920 15184 19228 15204
rect 19156 14816 19208 14822
rect 19156 14758 19208 14764
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 18696 14408 18748 14414
rect 18696 14350 18748 14356
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18708 13025 18736 14350
rect 18800 14074 18828 14350
rect 19168 14346 19196 14758
rect 19156 14340 19208 14346
rect 19156 14282 19208 14288
rect 19260 14226 19288 19196
rect 19444 18952 19472 19790
rect 19352 18924 19472 18952
rect 19352 17218 19380 18924
rect 19536 18816 19564 20402
rect 19628 19514 19656 20878
rect 19708 20596 19760 20602
rect 19708 20538 19760 20544
rect 19720 20346 19748 20538
rect 19904 20466 19932 21014
rect 19892 20460 19944 20466
rect 19892 20402 19944 20408
rect 19720 20318 19932 20346
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 19616 19508 19668 19514
rect 19616 19450 19668 19456
rect 19616 19168 19668 19174
rect 19616 19110 19668 19116
rect 19444 18788 19564 18816
rect 19444 18290 19472 18788
rect 19515 18736 19567 18742
rect 19515 18678 19567 18684
rect 19527 18652 19564 18678
rect 19536 18426 19564 18652
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 19522 18320 19578 18329
rect 19432 18284 19484 18290
rect 19628 18290 19656 19110
rect 19720 18290 19748 19858
rect 19800 19712 19852 19718
rect 19800 19654 19852 19660
rect 19522 18255 19578 18264
rect 19616 18284 19668 18290
rect 19432 18226 19484 18232
rect 19536 17338 19564 18255
rect 19616 18226 19668 18232
rect 19708 18284 19760 18290
rect 19708 18226 19760 18232
rect 19720 17354 19748 18226
rect 19524 17332 19576 17338
rect 19524 17274 19576 17280
rect 19628 17326 19748 17354
rect 19352 17190 19564 17218
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19352 16658 19380 17070
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 19352 15978 19380 16594
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19340 15972 19392 15978
rect 19340 15914 19392 15920
rect 19340 15360 19392 15366
rect 19340 15302 19392 15308
rect 19352 15162 19380 15302
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 19352 14346 19380 14418
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19260 14198 19380 14226
rect 18920 14172 19228 14192
rect 18920 14170 18926 14172
rect 18982 14170 19006 14172
rect 19062 14170 19086 14172
rect 19142 14170 19166 14172
rect 19222 14170 19228 14172
rect 18982 14118 18984 14170
rect 19164 14118 19166 14170
rect 18920 14116 18926 14118
rect 18982 14116 19006 14118
rect 19062 14116 19086 14118
rect 19142 14116 19166 14118
rect 19222 14116 19228 14118
rect 18920 14096 19228 14116
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19154 13968 19210 13977
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 19064 13932 19116 13938
rect 19154 13903 19210 13912
rect 19064 13874 19116 13880
rect 18788 13524 18840 13530
rect 18788 13466 18840 13472
rect 18800 13326 18828 13466
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 18892 13172 18920 13874
rect 19076 13530 19104 13874
rect 19168 13870 19196 13903
rect 19156 13864 19208 13870
rect 19156 13806 19208 13812
rect 19154 13560 19210 13569
rect 19064 13524 19116 13530
rect 19154 13495 19210 13504
rect 19064 13466 19116 13472
rect 19168 13258 19196 13495
rect 19156 13252 19208 13258
rect 19156 13194 19208 13200
rect 18800 13144 18920 13172
rect 18694 13016 18750 13025
rect 18694 12951 18750 12960
rect 18616 12294 18736 12322
rect 18604 12164 18656 12170
rect 18604 12106 18656 12112
rect 18616 11898 18644 12106
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18604 9988 18656 9994
rect 18604 9930 18656 9936
rect 18616 7954 18644 9930
rect 18708 9110 18736 12294
rect 18800 11354 18828 13144
rect 18920 13084 19228 13104
rect 18920 13082 18926 13084
rect 18982 13082 19006 13084
rect 19062 13082 19086 13084
rect 19142 13082 19166 13084
rect 19222 13082 19228 13084
rect 18982 13030 18984 13082
rect 19164 13030 19166 13082
rect 18920 13028 18926 13030
rect 18982 13028 19006 13030
rect 19062 13028 19086 13030
rect 19142 13028 19166 13030
rect 19222 13028 19228 13030
rect 18920 13008 19228 13028
rect 19260 12968 19288 14010
rect 18984 12940 19288 12968
rect 18984 12209 19012 12940
rect 19352 12866 19380 14198
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 19168 12838 19380 12866
rect 19076 12306 19104 12786
rect 19064 12300 19116 12306
rect 19064 12242 19116 12248
rect 18970 12200 19026 12209
rect 19168 12170 19196 12838
rect 19444 12434 19472 16526
rect 19536 14482 19564 17190
rect 19628 16794 19656 17326
rect 19708 17264 19760 17270
rect 19708 17206 19760 17212
rect 19616 16788 19668 16794
rect 19616 16730 19668 16736
rect 19628 15638 19656 16730
rect 19616 15632 19668 15638
rect 19616 15574 19668 15580
rect 19616 14544 19668 14550
rect 19616 14486 19668 14492
rect 19524 14476 19576 14482
rect 19524 14418 19576 14424
rect 19524 14000 19576 14006
rect 19522 13968 19524 13977
rect 19576 13968 19578 13977
rect 19628 13938 19656 14486
rect 19522 13903 19578 13912
rect 19616 13932 19668 13938
rect 19616 13874 19668 13880
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 19536 13376 19564 13670
rect 19527 13348 19564 13376
rect 19527 13258 19555 13348
rect 19616 13298 19668 13304
rect 19524 13252 19576 13258
rect 19616 13240 19668 13246
rect 19524 13194 19576 13200
rect 19522 13152 19578 13161
rect 19522 13087 19578 13096
rect 19536 12986 19564 13087
rect 19628 12986 19656 13240
rect 19524 12980 19576 12986
rect 19524 12922 19576 12928
rect 19616 12980 19668 12986
rect 19616 12922 19668 12928
rect 19720 12434 19748 17206
rect 19352 12406 19472 12434
rect 19628 12406 19748 12434
rect 19352 12220 19380 12406
rect 19260 12192 19380 12220
rect 18970 12135 19026 12144
rect 19156 12164 19208 12170
rect 19156 12106 19208 12112
rect 18920 11996 19228 12016
rect 18920 11994 18926 11996
rect 18982 11994 19006 11996
rect 19062 11994 19086 11996
rect 19142 11994 19166 11996
rect 19222 11994 19228 11996
rect 18982 11942 18984 11994
rect 19164 11942 19166 11994
rect 18920 11940 18926 11942
rect 18982 11940 19006 11942
rect 19062 11940 19086 11942
rect 19142 11940 19166 11942
rect 19222 11940 19228 11942
rect 18920 11920 19228 11940
rect 18878 11792 18934 11801
rect 18878 11727 18880 11736
rect 18932 11727 18934 11736
rect 19156 11756 19208 11762
rect 18880 11698 18932 11704
rect 19156 11698 19208 11704
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18892 11234 18920 11698
rect 18800 11206 18920 11234
rect 18800 9364 18828 11206
rect 19168 11082 19196 11698
rect 19156 11076 19208 11082
rect 19156 11018 19208 11024
rect 18920 10908 19228 10928
rect 18920 10906 18926 10908
rect 18982 10906 19006 10908
rect 19062 10906 19086 10908
rect 19142 10906 19166 10908
rect 19222 10906 19228 10908
rect 18982 10854 18984 10906
rect 19164 10854 19166 10906
rect 18920 10852 18926 10854
rect 18982 10852 19006 10854
rect 19062 10852 19086 10854
rect 19142 10852 19166 10854
rect 19222 10852 19228 10854
rect 18920 10832 19228 10852
rect 19260 10792 19288 12192
rect 19432 11824 19484 11830
rect 19432 11766 19484 11772
rect 19444 11082 19472 11766
rect 19524 11620 19576 11626
rect 19524 11562 19576 11568
rect 19536 11082 19564 11562
rect 19432 11076 19484 11082
rect 19432 11018 19484 11024
rect 19524 11076 19576 11082
rect 19524 11018 19576 11024
rect 19168 10764 19288 10792
rect 19168 10606 19196 10764
rect 19246 10704 19302 10713
rect 19246 10639 19302 10648
rect 19524 10668 19576 10674
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 18920 9820 19228 9840
rect 18920 9818 18926 9820
rect 18982 9818 19006 9820
rect 19062 9818 19086 9820
rect 19142 9818 19166 9820
rect 19222 9818 19228 9820
rect 18982 9766 18984 9818
rect 19164 9766 19166 9818
rect 18920 9764 18926 9766
rect 18982 9764 19006 9766
rect 19062 9764 19086 9766
rect 19142 9764 19166 9766
rect 19222 9764 19228 9766
rect 18920 9744 19228 9764
rect 19260 9602 19288 10639
rect 19524 10610 19576 10616
rect 19430 10568 19486 10577
rect 19430 10503 19486 10512
rect 19338 10160 19394 10169
rect 19444 10146 19472 10503
rect 19536 10266 19564 10610
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 19444 10118 19564 10146
rect 19338 10095 19394 10104
rect 19352 10062 19380 10095
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 19430 10024 19486 10033
rect 19352 9654 19380 9998
rect 19430 9959 19432 9968
rect 19484 9959 19486 9968
rect 19432 9930 19484 9936
rect 19168 9574 19288 9602
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 18800 9336 18920 9364
rect 18696 9104 18748 9110
rect 18696 9046 18748 9052
rect 18694 8936 18750 8945
rect 18892 8888 18920 9336
rect 18694 8871 18750 8880
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18616 4010 18644 6054
rect 18604 4004 18656 4010
rect 18604 3946 18656 3952
rect 18616 3602 18644 3946
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 18708 3534 18736 8871
rect 18800 8860 18920 8888
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18800 3398 18828 8860
rect 19168 8820 19196 9574
rect 19246 9072 19302 9081
rect 19246 9007 19302 9016
rect 19260 8974 19288 9007
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19352 8906 19380 9590
rect 19444 8974 19472 9930
rect 19536 9722 19564 10118
rect 19524 9716 19576 9722
rect 19524 9658 19576 9664
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 19340 8900 19392 8906
rect 19340 8842 19392 8848
rect 19168 8792 19288 8820
rect 18920 8732 19228 8752
rect 18920 8730 18926 8732
rect 18982 8730 19006 8732
rect 19062 8730 19086 8732
rect 19142 8730 19166 8732
rect 19222 8730 19228 8732
rect 18982 8678 18984 8730
rect 19164 8678 19166 8730
rect 18920 8676 18926 8678
rect 18982 8676 19006 8678
rect 19062 8676 19086 8678
rect 19142 8676 19166 8678
rect 19222 8676 19228 8678
rect 18920 8656 19228 8676
rect 19260 8022 19288 8792
rect 19536 8786 19564 9522
rect 19444 8758 19564 8786
rect 19444 8430 19472 8758
rect 19524 8628 19576 8634
rect 19524 8570 19576 8576
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19430 8256 19486 8265
rect 19430 8191 19486 8200
rect 19248 8016 19300 8022
rect 19248 7958 19300 7964
rect 19248 7812 19300 7818
rect 19248 7754 19300 7760
rect 19340 7812 19392 7818
rect 19340 7754 19392 7760
rect 18920 7644 19228 7664
rect 18920 7642 18926 7644
rect 18982 7642 19006 7644
rect 19062 7642 19086 7644
rect 19142 7642 19166 7644
rect 19222 7642 19228 7644
rect 18982 7590 18984 7642
rect 19164 7590 19166 7642
rect 18920 7588 18926 7590
rect 18982 7588 19006 7590
rect 19062 7588 19086 7590
rect 19142 7588 19166 7590
rect 19222 7588 19228 7590
rect 18920 7568 19228 7588
rect 19260 7546 19288 7754
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 19076 7206 19104 7346
rect 19352 7342 19380 7754
rect 19444 7410 19472 8191
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19064 7200 19116 7206
rect 19064 7142 19116 7148
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19076 6798 19104 7142
rect 19352 6934 19380 7142
rect 19340 6928 19392 6934
rect 19340 6870 19392 6876
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 18920 6556 19228 6576
rect 18920 6554 18926 6556
rect 18982 6554 19006 6556
rect 19062 6554 19086 6556
rect 19142 6554 19166 6556
rect 19222 6554 19228 6556
rect 18982 6502 18984 6554
rect 19164 6502 19166 6554
rect 18920 6500 18926 6502
rect 18982 6500 19006 6502
rect 19062 6500 19086 6502
rect 19142 6500 19166 6502
rect 19222 6500 19228 6502
rect 18920 6480 19228 6500
rect 19352 6254 19380 6870
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19340 6248 19392 6254
rect 19340 6190 19392 6196
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19248 5568 19300 5574
rect 19248 5510 19300 5516
rect 18920 5468 19228 5488
rect 18920 5466 18926 5468
rect 18982 5466 19006 5468
rect 19062 5466 19086 5468
rect 19142 5466 19166 5468
rect 19222 5466 19228 5468
rect 18982 5414 18984 5466
rect 19164 5414 19166 5466
rect 18920 5412 18926 5414
rect 18982 5412 19006 5414
rect 19062 5412 19086 5414
rect 19142 5412 19166 5414
rect 19222 5412 19228 5414
rect 18920 5392 19228 5412
rect 19260 5250 19288 5510
rect 19076 5222 19288 5250
rect 19076 4554 19104 5222
rect 19064 4548 19116 4554
rect 19064 4490 19116 4496
rect 18920 4380 19228 4400
rect 18920 4378 18926 4380
rect 18982 4378 19006 4380
rect 19062 4378 19086 4380
rect 19142 4378 19166 4380
rect 19222 4378 19228 4380
rect 18982 4326 18984 4378
rect 19164 4326 19166 4378
rect 18920 4324 18926 4326
rect 18982 4324 19006 4326
rect 19062 4324 19086 4326
rect 19142 4324 19166 4326
rect 19222 4324 19228 4326
rect 18920 4304 19228 4324
rect 19352 4146 19380 5646
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 19444 4078 19472 6258
rect 19536 4214 19564 8570
rect 19628 7528 19656 12406
rect 19706 12336 19762 12345
rect 19706 12271 19708 12280
rect 19760 12271 19762 12280
rect 19708 12242 19760 12248
rect 19812 11898 19840 19654
rect 19904 18630 19932 20318
rect 19996 19854 20024 22066
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 19892 18624 19944 18630
rect 19892 18566 19944 18572
rect 19904 18222 19932 18566
rect 19996 18222 20024 19790
rect 20088 19378 20116 24754
rect 20180 24274 20208 25094
rect 20168 24268 20220 24274
rect 20168 24210 20220 24216
rect 20272 24154 20300 25214
rect 20352 24948 20404 24954
rect 20352 24890 20404 24896
rect 20180 24126 20300 24154
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 20074 19272 20130 19281
rect 20074 19207 20130 19216
rect 20088 19174 20116 19207
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 19892 18216 19944 18222
rect 19892 18158 19944 18164
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 19904 17354 19932 18158
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19996 17746 20024 18022
rect 20076 17808 20128 17814
rect 20076 17750 20128 17756
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 19904 17326 20024 17354
rect 19892 16108 19944 16114
rect 19892 16050 19944 16056
rect 19904 15706 19932 16050
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19890 15056 19946 15065
rect 19890 14991 19946 15000
rect 19904 14958 19932 14991
rect 19892 14952 19944 14958
rect 19892 14894 19944 14900
rect 19890 14648 19946 14657
rect 19890 14583 19892 14592
rect 19944 14583 19946 14592
rect 19892 14554 19944 14560
rect 19892 14000 19944 14006
rect 19892 13942 19944 13948
rect 19904 13841 19932 13942
rect 19890 13832 19946 13841
rect 19890 13767 19946 13776
rect 19996 13716 20024 17326
rect 20088 17134 20116 17750
rect 20180 17270 20208 24126
rect 20260 24064 20312 24070
rect 20260 24006 20312 24012
rect 20168 17264 20220 17270
rect 20168 17206 20220 17212
rect 20076 17128 20128 17134
rect 20076 17070 20128 17076
rect 20168 16448 20220 16454
rect 20168 16390 20220 16396
rect 20076 15496 20128 15502
rect 20076 15438 20128 15444
rect 19904 13688 20024 13716
rect 19904 13394 19932 13688
rect 20088 13410 20116 15438
rect 19892 13388 19944 13394
rect 19892 13330 19944 13336
rect 19996 13382 20116 13410
rect 19996 12730 20024 13382
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 20088 13190 20116 13262
rect 20076 13184 20128 13190
rect 20076 13126 20128 13132
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 19904 12702 20024 12730
rect 19904 12646 19932 12702
rect 19892 12640 19944 12646
rect 19892 12582 19944 12588
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 19800 11892 19852 11898
rect 19800 11834 19852 11840
rect 19800 11688 19852 11694
rect 19800 11630 19852 11636
rect 19708 11144 19760 11150
rect 19708 11086 19760 11092
rect 19720 10674 19748 11086
rect 19812 11082 19840 11630
rect 19890 11248 19946 11257
rect 19890 11183 19946 11192
rect 19800 11076 19852 11082
rect 19800 11018 19852 11024
rect 19708 10668 19760 10674
rect 19708 10610 19760 10616
rect 19904 9586 19932 11183
rect 19800 9580 19852 9586
rect 19800 9522 19852 9528
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19720 8498 19748 9318
rect 19812 9178 19840 9522
rect 19800 9172 19852 9178
rect 19800 9114 19852 9120
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19708 8492 19760 8498
rect 19708 8434 19760 8440
rect 19904 7886 19932 8910
rect 19996 8634 20024 12582
rect 20088 12374 20116 12922
rect 20076 12368 20128 12374
rect 20076 12310 20128 12316
rect 20076 12164 20128 12170
rect 20076 12106 20128 12112
rect 20088 11898 20116 12106
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 20088 10554 20116 11834
rect 20180 10742 20208 16390
rect 20272 11744 20300 24006
rect 20364 22710 20392 24890
rect 20626 24848 20682 24857
rect 20626 24783 20682 24792
rect 20536 24744 20588 24750
rect 20536 24686 20588 24692
rect 20444 24200 20496 24206
rect 20444 24142 20496 24148
rect 20352 22704 20404 22710
rect 20352 22646 20404 22652
rect 20352 22568 20404 22574
rect 20352 22510 20404 22516
rect 20364 20942 20392 22510
rect 20352 20936 20404 20942
rect 20352 20878 20404 20884
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 20364 19854 20392 20742
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 20350 19272 20406 19281
rect 20350 19207 20406 19216
rect 20364 13802 20392 19207
rect 20352 13796 20404 13802
rect 20352 13738 20404 13744
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 20364 12850 20392 13466
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20364 11898 20392 12582
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20272 11716 20392 11744
rect 20260 11620 20312 11626
rect 20260 11562 20312 11568
rect 20168 10736 20220 10742
rect 20168 10678 20220 10684
rect 20088 10526 20208 10554
rect 20076 8900 20128 8906
rect 20076 8842 20128 8848
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 20088 8362 20116 8842
rect 20076 8356 20128 8362
rect 20076 8298 20128 8304
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19628 7500 19840 7528
rect 19616 7404 19668 7410
rect 19616 7346 19668 7352
rect 19628 6866 19656 7346
rect 19616 6860 19668 6866
rect 19616 6802 19668 6808
rect 19708 6792 19760 6798
rect 19708 6734 19760 6740
rect 19720 6390 19748 6734
rect 19708 6384 19760 6390
rect 19708 6326 19760 6332
rect 19708 6180 19760 6186
rect 19708 6122 19760 6128
rect 19616 5772 19668 5778
rect 19616 5714 19668 5720
rect 19524 4208 19576 4214
rect 19524 4150 19576 4156
rect 19432 4072 19484 4078
rect 19338 4040 19394 4049
rect 19432 4014 19484 4020
rect 19524 4072 19576 4078
rect 19524 4014 19576 4020
rect 19338 3975 19394 3984
rect 19352 3466 19380 3975
rect 19430 3904 19486 3913
rect 19430 3839 19486 3848
rect 19444 3534 19472 3839
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18920 3292 19228 3312
rect 18920 3290 18926 3292
rect 18982 3290 19006 3292
rect 19062 3290 19086 3292
rect 19142 3290 19166 3292
rect 19222 3290 19228 3292
rect 18982 3238 18984 3290
rect 19164 3238 19166 3290
rect 18920 3236 18926 3238
rect 18982 3236 19006 3238
rect 19062 3236 19086 3238
rect 19142 3236 19166 3238
rect 19222 3236 19228 3238
rect 18786 3224 18842 3233
rect 18920 3216 19228 3236
rect 18786 3159 18842 3168
rect 18696 3052 18748 3058
rect 18524 3012 18696 3040
rect 18696 2994 18748 3000
rect 18340 2746 18736 2774
rect 18236 2372 18288 2378
rect 18236 2314 18288 2320
rect 18420 2304 18472 2310
rect 18420 2246 18472 2252
rect 18432 800 18460 2246
rect 18708 800 18736 2746
rect 18800 1086 18828 3159
rect 19536 2922 19564 4014
rect 19524 2916 19576 2922
rect 19524 2858 19576 2864
rect 19248 2576 19300 2582
rect 19248 2518 19300 2524
rect 18920 2204 19228 2224
rect 18920 2202 18926 2204
rect 18982 2202 19006 2204
rect 19062 2202 19086 2204
rect 19142 2202 19166 2204
rect 19222 2202 19228 2204
rect 18982 2150 18984 2202
rect 19164 2150 19166 2202
rect 18920 2148 18926 2150
rect 18982 2148 19006 2150
rect 19062 2148 19086 2150
rect 19142 2148 19166 2150
rect 19222 2148 19228 2150
rect 18920 2128 19228 2148
rect 19260 1170 19288 2518
rect 19628 2446 19656 5714
rect 19720 2922 19748 6122
rect 19708 2916 19760 2922
rect 19708 2858 19760 2864
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19524 1964 19576 1970
rect 19524 1906 19576 1912
rect 18984 1142 19288 1170
rect 18788 1080 18840 1086
rect 18788 1022 18840 1028
rect 18984 800 19012 1142
rect 19248 1080 19300 1086
rect 19248 1022 19300 1028
rect 19260 800 19288 1022
rect 19536 800 19564 1906
rect 19812 800 19840 7500
rect 19904 6798 19932 7822
rect 20180 7528 20208 10526
rect 20272 9674 20300 11562
rect 20364 11150 20392 11716
rect 20456 11354 20484 24142
rect 20548 23866 20576 24686
rect 20536 23860 20588 23866
rect 20536 23802 20588 23808
rect 20640 23474 20668 24783
rect 20732 24410 20760 26200
rect 20824 25838 20852 26726
rect 20904 25968 20956 25974
rect 20904 25910 20956 25916
rect 20812 25832 20864 25838
rect 20812 25774 20864 25780
rect 20824 25226 20852 25774
rect 20812 25220 20864 25226
rect 20812 25162 20864 25168
rect 20720 24404 20772 24410
rect 20720 24346 20772 24352
rect 20720 24064 20772 24070
rect 20720 24006 20772 24012
rect 20548 23446 20668 23474
rect 20548 22658 20576 23446
rect 20628 23316 20680 23322
rect 20628 23258 20680 23264
rect 20640 22778 20668 23258
rect 20732 23089 20760 24006
rect 20718 23080 20774 23089
rect 20718 23015 20774 23024
rect 20824 22964 20852 25162
rect 20916 23662 20944 25910
rect 20904 23656 20956 23662
rect 20904 23598 20956 23604
rect 20916 23254 20944 23598
rect 20904 23248 20956 23254
rect 20904 23190 20956 23196
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 20732 22936 20852 22964
rect 20628 22772 20680 22778
rect 20628 22714 20680 22720
rect 20548 22630 20668 22658
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 20548 22234 20576 22510
rect 20536 22228 20588 22234
rect 20536 22170 20588 22176
rect 20548 21486 20576 22170
rect 20640 21690 20668 22630
rect 20628 21684 20680 21690
rect 20628 21626 20680 21632
rect 20626 21584 20682 21593
rect 20626 21519 20682 21528
rect 20536 21480 20588 21486
rect 20536 21422 20588 21428
rect 20640 21350 20668 21519
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 20548 18426 20576 20878
rect 20640 20466 20668 21286
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 20640 19718 20668 20402
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20536 18420 20588 18426
rect 20536 18362 20588 18368
rect 20640 18306 20668 19450
rect 20548 18278 20668 18306
rect 20548 17202 20576 18278
rect 20732 17814 20760 22936
rect 20812 22772 20864 22778
rect 20812 22714 20864 22720
rect 20824 22574 20852 22714
rect 20812 22568 20864 22574
rect 20812 22510 20864 22516
rect 20824 21622 20852 22510
rect 20916 22506 20944 23054
rect 20904 22500 20956 22506
rect 20904 22442 20956 22448
rect 20916 22098 20944 22442
rect 20904 22092 20956 22098
rect 20904 22034 20956 22040
rect 20904 21956 20956 21962
rect 20904 21898 20956 21904
rect 20812 21616 20864 21622
rect 20812 21558 20864 21564
rect 20916 21350 20944 21898
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 20824 18358 20852 21082
rect 21008 21026 21036 27814
rect 21652 27674 21680 28494
rect 21824 28484 21876 28490
rect 21824 28426 21876 28432
rect 21836 27674 21864 28426
rect 21640 27668 21692 27674
rect 21640 27610 21692 27616
rect 21824 27668 21876 27674
rect 21824 27610 21876 27616
rect 21824 27532 21876 27538
rect 21824 27474 21876 27480
rect 21180 27464 21232 27470
rect 21180 27406 21232 27412
rect 21192 26382 21220 27406
rect 21548 27328 21600 27334
rect 21548 27270 21600 27276
rect 21272 26988 21324 26994
rect 21272 26930 21324 26936
rect 21180 26376 21232 26382
rect 21180 26318 21232 26324
rect 21088 25900 21140 25906
rect 21088 25842 21140 25848
rect 21180 25900 21232 25906
rect 21180 25842 21232 25848
rect 21100 25294 21128 25842
rect 21088 25288 21140 25294
rect 21088 25230 21140 25236
rect 21192 24954 21220 25842
rect 21180 24948 21232 24954
rect 21180 24890 21232 24896
rect 21284 24857 21312 26930
rect 21456 26852 21508 26858
rect 21456 26794 21508 26800
rect 21468 26586 21496 26794
rect 21456 26580 21508 26586
rect 21456 26522 21508 26528
rect 21364 25288 21416 25294
rect 21364 25230 21416 25236
rect 21270 24848 21326 24857
rect 21180 24812 21232 24818
rect 21270 24783 21326 24792
rect 21180 24754 21232 24760
rect 21088 24608 21140 24614
rect 21088 24550 21140 24556
rect 21100 23497 21128 24550
rect 21192 23769 21220 24754
rect 21272 24676 21324 24682
rect 21272 24618 21324 24624
rect 21284 24313 21312 24618
rect 21270 24304 21326 24313
rect 21270 24239 21326 24248
rect 21272 24132 21324 24138
rect 21272 24074 21324 24080
rect 21178 23760 21234 23769
rect 21178 23695 21234 23704
rect 21180 23588 21232 23594
rect 21180 23530 21232 23536
rect 21086 23488 21142 23497
rect 21086 23423 21142 23432
rect 21192 23254 21220 23530
rect 21180 23248 21232 23254
rect 21178 23216 21180 23225
rect 21232 23216 21234 23225
rect 21088 23180 21140 23186
rect 21178 23151 21234 23160
rect 21088 23122 21140 23128
rect 21100 23066 21128 23122
rect 21100 23038 21220 23066
rect 21086 22944 21142 22953
rect 21086 22879 21142 22888
rect 21100 21146 21128 22879
rect 21088 21140 21140 21146
rect 21088 21082 21140 21088
rect 20916 20998 21036 21026
rect 20916 20482 20944 20998
rect 21192 20942 21220 23038
rect 21284 22953 21312 24074
rect 21270 22944 21326 22953
rect 21270 22879 21326 22888
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 21180 20936 21232 20942
rect 21376 20890 21404 25230
rect 21456 24132 21508 24138
rect 21456 24074 21508 24080
rect 21468 24041 21496 24074
rect 21454 24032 21510 24041
rect 21454 23967 21510 23976
rect 21560 23361 21588 27270
rect 21640 26784 21692 26790
rect 21640 26726 21692 26732
rect 21652 24274 21680 26726
rect 21836 26450 21864 27474
rect 22112 27470 22140 28630
rect 22928 28552 22980 28558
rect 22928 28494 22980 28500
rect 27344 28552 27396 28558
rect 27344 28494 27396 28500
rect 22192 28416 22244 28422
rect 22192 28358 22244 28364
rect 22100 27464 22152 27470
rect 22100 27406 22152 27412
rect 22008 26988 22060 26994
rect 22008 26930 22060 26936
rect 21824 26444 21876 26450
rect 21824 26386 21876 26392
rect 22020 26042 22048 26930
rect 22008 26036 22060 26042
rect 22008 25978 22060 25984
rect 22100 25968 22152 25974
rect 21822 25936 21878 25945
rect 22100 25910 22152 25916
rect 21822 25871 21824 25880
rect 21876 25871 21878 25880
rect 21916 25900 21968 25906
rect 21824 25842 21876 25848
rect 21916 25842 21968 25848
rect 21836 25294 21864 25842
rect 21824 25288 21876 25294
rect 21824 25230 21876 25236
rect 21732 25152 21784 25158
rect 21732 25094 21784 25100
rect 21640 24268 21692 24274
rect 21640 24210 21692 24216
rect 21640 23724 21692 23730
rect 21640 23666 21692 23672
rect 21652 23633 21680 23666
rect 21638 23624 21694 23633
rect 21638 23559 21694 23568
rect 21546 23352 21602 23361
rect 21546 23287 21602 23296
rect 21548 23180 21600 23186
rect 21548 23122 21600 23128
rect 21456 23044 21508 23050
rect 21456 22986 21508 22992
rect 21180 20878 21232 20884
rect 20996 20868 21048 20874
rect 20996 20810 21048 20816
rect 21008 20602 21036 20810
rect 20996 20596 21048 20602
rect 20996 20538 21048 20544
rect 20916 20454 21036 20482
rect 20904 18692 20956 18698
rect 20904 18634 20956 18640
rect 20916 18426 20944 18634
rect 20904 18420 20956 18426
rect 20904 18362 20956 18368
rect 20812 18352 20864 18358
rect 20812 18294 20864 18300
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 20812 18148 20864 18154
rect 20812 18090 20864 18096
rect 20720 17808 20772 17814
rect 20720 17750 20772 17756
rect 20824 17678 20852 18090
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20628 17604 20680 17610
rect 20628 17546 20680 17552
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20548 14521 20576 17138
rect 20640 16182 20668 17546
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 20718 17232 20774 17241
rect 20718 17167 20774 17176
rect 20628 16176 20680 16182
rect 20628 16118 20680 16124
rect 20640 15638 20668 16118
rect 20628 15632 20680 15638
rect 20628 15574 20680 15580
rect 20732 15570 20760 17167
rect 20824 17066 20852 17274
rect 20812 17060 20864 17066
rect 20812 17002 20864 17008
rect 20812 16720 20864 16726
rect 20812 16662 20864 16668
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20824 15450 20852 16662
rect 20916 15706 20944 18226
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 21008 15586 21036 20454
rect 21100 20058 21128 20878
rect 21284 20862 21404 20890
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 21178 19136 21234 19145
rect 21178 19071 21234 19080
rect 21192 18154 21220 19071
rect 21180 18148 21232 18154
rect 21180 18090 21232 18096
rect 21088 18080 21140 18086
rect 21088 18022 21140 18028
rect 21100 17678 21128 18022
rect 21088 17672 21140 17678
rect 21088 17614 21140 17620
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 21100 17241 21128 17478
rect 21086 17232 21142 17241
rect 21192 17202 21220 18090
rect 21086 17167 21142 17176
rect 21180 17196 21232 17202
rect 21180 17138 21232 17144
rect 21088 17128 21140 17134
rect 21088 17070 21140 17076
rect 21100 16454 21128 17070
rect 21192 16969 21220 17138
rect 21178 16960 21234 16969
rect 21178 16895 21234 16904
rect 21192 16590 21220 16895
rect 21180 16584 21232 16590
rect 21180 16526 21232 16532
rect 21088 16448 21140 16454
rect 21088 16390 21140 16396
rect 21180 15904 21232 15910
rect 21180 15846 21232 15852
rect 20640 15422 20852 15450
rect 20916 15558 21036 15586
rect 21086 15600 21142 15609
rect 20640 15366 20668 15422
rect 20628 15360 20680 15366
rect 20628 15302 20680 15308
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20732 15201 20760 15302
rect 20718 15192 20774 15201
rect 20640 15150 20718 15178
rect 20534 14512 20590 14521
rect 20534 14447 20590 14456
rect 20640 13802 20668 15150
rect 20718 15127 20774 15136
rect 20720 15088 20772 15094
rect 20720 15030 20772 15036
rect 20732 14074 20760 15030
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20628 13796 20680 13802
rect 20628 13738 20680 13744
rect 20732 13734 20760 14010
rect 20720 13728 20772 13734
rect 20720 13670 20772 13676
rect 20534 13424 20590 13433
rect 20732 13394 20760 13670
rect 20534 13359 20590 13368
rect 20720 13388 20772 13394
rect 20548 12170 20576 13359
rect 20720 13330 20772 13336
rect 20628 13320 20680 13326
rect 20628 13262 20680 13268
rect 20640 13161 20668 13262
rect 20720 13184 20772 13190
rect 20626 13152 20682 13161
rect 20720 13126 20772 13132
rect 20626 13087 20682 13096
rect 20732 12850 20760 13126
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20536 12164 20588 12170
rect 20536 12106 20588 12112
rect 20628 12164 20680 12170
rect 20628 12106 20680 12112
rect 20640 11626 20668 12106
rect 20628 11620 20680 11626
rect 20628 11562 20680 11568
rect 20536 11552 20588 11558
rect 20536 11494 20588 11500
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 20352 11144 20404 11150
rect 20352 11086 20404 11092
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 20456 9761 20484 10202
rect 20442 9752 20498 9761
rect 20442 9687 20498 9696
rect 20272 9646 20392 9674
rect 20260 9104 20312 9110
rect 20260 9046 20312 9052
rect 20272 8634 20300 9046
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 19996 7500 20208 7528
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 19904 6322 19932 6734
rect 19892 6316 19944 6322
rect 19892 6258 19944 6264
rect 19892 6180 19944 6186
rect 19996 6168 20024 7500
rect 20364 7449 20392 9646
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20456 9178 20484 9318
rect 20444 9172 20496 9178
rect 20444 9114 20496 9120
rect 20442 8800 20498 8809
rect 20442 8735 20498 8744
rect 20350 7440 20406 7449
rect 20168 7404 20220 7410
rect 20456 7410 20484 8735
rect 20350 7375 20406 7384
rect 20444 7404 20496 7410
rect 20168 7346 20220 7352
rect 20444 7346 20496 7352
rect 20180 6390 20208 7346
rect 20548 7290 20576 11494
rect 20718 10840 20774 10849
rect 20718 10775 20720 10784
rect 20772 10775 20774 10784
rect 20720 10746 20772 10752
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20640 7546 20668 10406
rect 20732 9926 20760 10746
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20364 7262 20576 7290
rect 20168 6384 20220 6390
rect 20168 6326 20220 6332
rect 19944 6140 20024 6168
rect 19892 6122 19944 6128
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 19892 5568 19944 5574
rect 19892 5510 19944 5516
rect 19904 2514 19932 5510
rect 19982 5264 20038 5273
rect 19982 5199 20038 5208
rect 19996 3058 20024 5199
rect 20088 3194 20116 5646
rect 20364 5624 20392 7262
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 20180 5596 20392 5624
rect 20076 3188 20128 3194
rect 20076 3130 20128 3136
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 20074 2952 20130 2961
rect 20074 2887 20076 2896
rect 20128 2887 20130 2896
rect 20076 2858 20128 2864
rect 20076 2644 20128 2650
rect 20180 2632 20208 5596
rect 20258 5536 20314 5545
rect 20258 5471 20314 5480
rect 20272 4554 20300 5471
rect 20352 5296 20404 5302
rect 20352 5238 20404 5244
rect 20364 5137 20392 5238
rect 20350 5128 20406 5137
rect 20350 5063 20406 5072
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 20364 4826 20392 4966
rect 20352 4820 20404 4826
rect 20352 4762 20404 4768
rect 20260 4548 20312 4554
rect 20260 4490 20312 4496
rect 20456 4146 20484 7142
rect 20536 5568 20588 5574
rect 20640 5556 20668 7482
rect 20732 6390 20760 9522
rect 20824 9518 20852 14962
rect 20916 13852 20944 15558
rect 21086 15535 21142 15544
rect 21100 15434 21128 15535
rect 21192 15502 21220 15846
rect 21180 15496 21232 15502
rect 21180 15438 21232 15444
rect 21088 15428 21140 15434
rect 21088 15370 21140 15376
rect 21180 14952 21232 14958
rect 21180 14894 21232 14900
rect 21088 14816 21140 14822
rect 21088 14758 21140 14764
rect 20916 13824 21036 13852
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 20916 12850 20944 13466
rect 21008 13025 21036 13824
rect 20994 13016 21050 13025
rect 20994 12951 21050 12960
rect 20904 12844 20956 12850
rect 20956 12804 21036 12832
rect 20904 12786 20956 12792
rect 21008 11898 21036 12804
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 20904 11008 20956 11014
rect 20902 10976 20904 10985
rect 20996 11008 21048 11014
rect 20956 10976 20958 10985
rect 20996 10950 21048 10956
rect 20902 10911 20958 10920
rect 20904 10736 20956 10742
rect 20904 10678 20956 10684
rect 20916 10062 20944 10678
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 20916 8922 20944 9998
rect 21008 9994 21036 10950
rect 20996 9988 21048 9994
rect 20996 9930 21048 9936
rect 21100 8974 21128 14758
rect 21192 13938 21220 14894
rect 21180 13932 21232 13938
rect 21180 13874 21232 13880
rect 21192 13258 21220 13874
rect 21180 13252 21232 13258
rect 21180 13194 21232 13200
rect 21192 12850 21220 13194
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 21192 12306 21220 12786
rect 21284 12617 21312 20862
rect 21364 20800 21416 20806
rect 21364 20742 21416 20748
rect 21376 20602 21404 20742
rect 21364 20596 21416 20602
rect 21364 20538 21416 20544
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21376 20058 21404 20198
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21376 12986 21404 18566
rect 21468 14249 21496 22986
rect 21560 22642 21588 23122
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21652 22778 21680 23054
rect 21640 22772 21692 22778
rect 21640 22714 21692 22720
rect 21548 22636 21600 22642
rect 21548 22578 21600 22584
rect 21640 22432 21692 22438
rect 21640 22374 21692 22380
rect 21652 22030 21680 22374
rect 21640 22024 21692 22030
rect 21640 21966 21692 21972
rect 21652 21350 21680 21966
rect 21640 21344 21692 21350
rect 21640 21286 21692 21292
rect 21640 20800 21692 20806
rect 21640 20742 21692 20748
rect 21548 17740 21600 17746
rect 21548 17682 21600 17688
rect 21560 17649 21588 17682
rect 21546 17640 21602 17649
rect 21546 17575 21602 17584
rect 21546 17232 21602 17241
rect 21546 17167 21602 17176
rect 21560 14618 21588 17167
rect 21548 14612 21600 14618
rect 21548 14554 21600 14560
rect 21546 14512 21602 14521
rect 21546 14447 21548 14456
rect 21600 14447 21602 14456
rect 21548 14418 21600 14424
rect 21548 14272 21600 14278
rect 21454 14240 21510 14249
rect 21548 14214 21600 14220
rect 21454 14175 21510 14184
rect 21560 14006 21588 14214
rect 21548 14000 21600 14006
rect 21454 13968 21510 13977
rect 21548 13942 21600 13948
rect 21454 13903 21510 13912
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21364 12640 21416 12646
rect 21270 12608 21326 12617
rect 21364 12582 21416 12588
rect 21270 12543 21326 12552
rect 21270 12472 21326 12481
rect 21270 12407 21326 12416
rect 21180 12300 21232 12306
rect 21180 12242 21232 12248
rect 21178 11928 21234 11937
rect 21178 11863 21234 11872
rect 21192 11830 21220 11863
rect 21180 11824 21232 11830
rect 21180 11766 21232 11772
rect 21180 11688 21232 11694
rect 21180 11630 21232 11636
rect 21192 10656 21220 11630
rect 21284 11014 21312 12407
rect 21272 11008 21324 11014
rect 21272 10950 21324 10956
rect 21376 10674 21404 12582
rect 21468 10810 21496 13903
rect 21548 13796 21600 13802
rect 21548 13738 21600 13744
rect 21560 13705 21588 13738
rect 21546 13696 21602 13705
rect 21546 13631 21602 13640
rect 21548 12776 21600 12782
rect 21548 12718 21600 12724
rect 21560 12442 21588 12718
rect 21652 12646 21680 20742
rect 21744 13977 21772 25094
rect 21928 24410 21956 25842
rect 22008 25220 22060 25226
rect 22008 25162 22060 25168
rect 22020 24954 22048 25162
rect 22008 24948 22060 24954
rect 22008 24890 22060 24896
rect 21916 24404 21968 24410
rect 21916 24346 21968 24352
rect 21916 24200 21968 24206
rect 21916 24142 21968 24148
rect 21824 24132 21876 24138
rect 21824 24074 21876 24080
rect 21836 21894 21864 24074
rect 21928 24070 21956 24142
rect 21916 24064 21968 24070
rect 22112 24041 22140 25910
rect 21916 24006 21968 24012
rect 22098 24032 22154 24041
rect 22098 23967 22154 23976
rect 21916 23656 21968 23662
rect 21916 23598 21968 23604
rect 21928 23186 21956 23598
rect 22008 23520 22060 23526
rect 22008 23462 22060 23468
rect 22020 23361 22048 23462
rect 22006 23352 22062 23361
rect 22204 23338 22232 28358
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22296 26858 22324 28018
rect 22376 27872 22428 27878
rect 22376 27814 22428 27820
rect 22744 27872 22796 27878
rect 22744 27814 22796 27820
rect 22284 26852 22336 26858
rect 22284 26794 22336 26800
rect 22388 26314 22416 27814
rect 22468 27396 22520 27402
rect 22468 27338 22520 27344
rect 22376 26308 22428 26314
rect 22376 26250 22428 26256
rect 22284 26240 22336 26246
rect 22284 26182 22336 26188
rect 22296 26042 22324 26182
rect 22284 26036 22336 26042
rect 22284 25978 22336 25984
rect 22284 25696 22336 25702
rect 22284 25638 22336 25644
rect 22296 25362 22324 25638
rect 22480 25498 22508 27338
rect 22652 26988 22704 26994
rect 22652 26930 22704 26936
rect 22664 26586 22692 26930
rect 22652 26580 22704 26586
rect 22652 26522 22704 26528
rect 22756 26466 22784 27814
rect 22836 26988 22888 26994
rect 22836 26930 22888 26936
rect 22664 26438 22784 26466
rect 22468 25492 22520 25498
rect 22468 25434 22520 25440
rect 22284 25356 22336 25362
rect 22284 25298 22336 25304
rect 22468 25220 22520 25226
rect 22468 25162 22520 25168
rect 22480 24886 22508 25162
rect 22468 24880 22520 24886
rect 22468 24822 22520 24828
rect 22376 24812 22428 24818
rect 22376 24754 22428 24760
rect 22560 24812 22612 24818
rect 22560 24754 22612 24760
rect 22388 24070 22416 24754
rect 22572 24410 22600 24754
rect 22560 24404 22612 24410
rect 22560 24346 22612 24352
rect 22560 24268 22612 24274
rect 22560 24210 22612 24216
rect 22284 24064 22336 24070
rect 22284 24006 22336 24012
rect 22376 24064 22428 24070
rect 22376 24006 22428 24012
rect 22296 23497 22324 24006
rect 22572 23866 22600 24210
rect 22560 23860 22612 23866
rect 22560 23802 22612 23808
rect 22376 23724 22428 23730
rect 22376 23666 22428 23672
rect 22388 23633 22416 23666
rect 22374 23624 22430 23633
rect 22374 23559 22430 23568
rect 22282 23488 22338 23497
rect 22282 23423 22338 23432
rect 22204 23310 22324 23338
rect 22006 23287 22008 23296
rect 22060 23287 22062 23296
rect 22008 23258 22060 23264
rect 21916 23180 21968 23186
rect 21916 23122 21968 23128
rect 22020 22098 22048 23258
rect 22192 23180 22244 23186
rect 22192 23122 22244 23128
rect 22204 22710 22232 23122
rect 22192 22704 22244 22710
rect 22192 22646 22244 22652
rect 22190 22264 22246 22273
rect 22190 22199 22246 22208
rect 22008 22092 22060 22098
rect 21928 22052 22008 22080
rect 21824 21888 21876 21894
rect 21824 21830 21876 21836
rect 21836 21554 21864 21830
rect 21824 21548 21876 21554
rect 21824 21490 21876 21496
rect 21928 21010 21956 22052
rect 22008 22034 22060 22040
rect 22008 21616 22060 21622
rect 22008 21558 22060 21564
rect 21916 21004 21968 21010
rect 21916 20946 21968 20952
rect 21824 20936 21876 20942
rect 21824 20878 21876 20884
rect 21836 20777 21864 20878
rect 21822 20768 21878 20777
rect 21822 20703 21878 20712
rect 21928 20584 21956 20946
rect 22020 20942 22048 21558
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 22008 20936 22060 20942
rect 22008 20878 22060 20884
rect 22008 20800 22060 20806
rect 22008 20742 22060 20748
rect 21836 20556 21956 20584
rect 21836 20466 21864 20556
rect 21824 20460 21876 20466
rect 21824 20402 21876 20408
rect 21916 20460 21968 20466
rect 21916 20402 21968 20408
rect 21928 18970 21956 20402
rect 22020 19417 22048 20742
rect 22112 19922 22140 21490
rect 22204 20466 22232 22199
rect 22296 20777 22324 23310
rect 22388 23050 22416 23559
rect 22560 23520 22612 23526
rect 22560 23462 22612 23468
rect 22572 23322 22600 23462
rect 22560 23316 22612 23322
rect 22560 23258 22612 23264
rect 22376 23044 22428 23050
rect 22376 22986 22428 22992
rect 22468 22976 22520 22982
rect 22468 22918 22520 22924
rect 22376 22636 22428 22642
rect 22376 22578 22428 22584
rect 22388 21146 22416 22578
rect 22376 21140 22428 21146
rect 22376 21082 22428 21088
rect 22282 20768 22338 20777
rect 22282 20703 22338 20712
rect 22388 20584 22416 21082
rect 22296 20556 22416 20584
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 22100 19916 22152 19922
rect 22100 19858 22152 19864
rect 22006 19408 22062 19417
rect 22006 19343 22062 19352
rect 21916 18964 21968 18970
rect 21916 18906 21968 18912
rect 22112 18834 22140 19858
rect 22296 19854 22324 20556
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22388 20058 22416 20402
rect 22376 20052 22428 20058
rect 22376 19994 22428 20000
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 22192 19780 22244 19786
rect 22192 19722 22244 19728
rect 22204 19666 22232 19722
rect 22204 19638 22324 19666
rect 22190 19544 22246 19553
rect 22190 19479 22246 19488
rect 22204 19446 22232 19479
rect 22192 19440 22244 19446
rect 22192 19382 22244 19388
rect 22296 19174 22324 19638
rect 22374 19544 22430 19553
rect 22374 19479 22376 19488
rect 22428 19479 22430 19488
rect 22376 19450 22428 19456
rect 22284 19168 22336 19174
rect 22284 19110 22336 19116
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 21824 18216 21876 18222
rect 21824 18158 21876 18164
rect 21836 17882 21864 18158
rect 21916 18148 21968 18154
rect 21916 18090 21968 18096
rect 21824 17876 21876 17882
rect 21824 17818 21876 17824
rect 21928 17678 21956 18090
rect 21916 17672 21968 17678
rect 21916 17614 21968 17620
rect 21822 17096 21878 17105
rect 21822 17031 21878 17040
rect 21836 16726 21864 17031
rect 21824 16720 21876 16726
rect 21824 16662 21876 16668
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 21836 15502 21864 16186
rect 21928 16046 21956 17614
rect 22020 16794 22048 18702
rect 22284 18624 22336 18630
rect 22284 18566 22336 18572
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22100 18420 22152 18426
rect 22100 18362 22152 18368
rect 22112 18329 22140 18362
rect 22098 18320 22154 18329
rect 22098 18255 22154 18264
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 22100 17604 22152 17610
rect 22100 17546 22152 17552
rect 22112 17270 22140 17546
rect 22100 17264 22152 17270
rect 22100 17206 22152 17212
rect 22100 17128 22152 17134
rect 22100 17070 22152 17076
rect 22008 16788 22060 16794
rect 22008 16730 22060 16736
rect 22112 16726 22140 17070
rect 22100 16720 22152 16726
rect 22006 16688 22062 16697
rect 22100 16662 22152 16668
rect 22006 16623 22062 16632
rect 22020 16590 22048 16623
rect 22008 16584 22060 16590
rect 22204 16572 22232 18226
rect 22008 16526 22060 16532
rect 22112 16544 22232 16572
rect 22008 16448 22060 16454
rect 22008 16390 22060 16396
rect 21916 16040 21968 16046
rect 21916 15982 21968 15988
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21824 14816 21876 14822
rect 21824 14758 21876 14764
rect 21836 14550 21864 14758
rect 21824 14544 21876 14550
rect 21824 14486 21876 14492
rect 21928 14414 21956 15982
rect 22020 15706 22048 16390
rect 22008 15700 22060 15706
rect 22008 15642 22060 15648
rect 22112 15638 22140 16544
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22100 15632 22152 15638
rect 22100 15574 22152 15580
rect 22204 15502 22232 15642
rect 22008 15496 22060 15502
rect 22192 15496 22244 15502
rect 22008 15438 22060 15444
rect 22112 15456 22192 15484
rect 21916 14408 21968 14414
rect 21916 14350 21968 14356
rect 22020 14056 22048 15438
rect 22112 14385 22140 15456
rect 22192 15438 22244 15444
rect 22192 15360 22244 15366
rect 22190 15328 22192 15337
rect 22244 15328 22246 15337
rect 22190 15263 22246 15272
rect 22190 15056 22246 15065
rect 22190 14991 22192 15000
rect 22244 14991 22246 15000
rect 22192 14962 22244 14968
rect 22296 14618 22324 18566
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 22098 14376 22154 14385
rect 22098 14311 22154 14320
rect 22284 14340 22336 14346
rect 22284 14282 22336 14288
rect 22100 14272 22152 14278
rect 22100 14214 22152 14220
rect 22190 14240 22246 14249
rect 21928 14028 22048 14056
rect 21730 13968 21786 13977
rect 21730 13903 21786 13912
rect 21824 13932 21876 13938
rect 21824 13874 21876 13880
rect 21732 13796 21784 13802
rect 21732 13738 21784 13744
rect 21744 13530 21772 13738
rect 21732 13524 21784 13530
rect 21732 13466 21784 13472
rect 21836 13326 21864 13874
rect 21928 13870 21956 14028
rect 22006 13968 22062 13977
rect 22006 13903 22062 13912
rect 21916 13864 21968 13870
rect 21916 13806 21968 13812
rect 21824 13320 21876 13326
rect 21824 13262 21876 13268
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 21824 12980 21876 12986
rect 21824 12922 21876 12928
rect 21732 12708 21784 12714
rect 21732 12650 21784 12656
rect 21640 12640 21692 12646
rect 21640 12582 21692 12588
rect 21548 12436 21600 12442
rect 21548 12378 21600 12384
rect 21744 12152 21772 12650
rect 21560 12124 21772 12152
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21364 10668 21416 10674
rect 21192 10628 21312 10656
rect 21178 10568 21234 10577
rect 21178 10503 21234 10512
rect 20824 8894 20944 8922
rect 21088 8968 21140 8974
rect 21088 8910 21140 8916
rect 20824 8498 20852 8894
rect 20904 8832 20956 8838
rect 20904 8774 20956 8780
rect 20996 8832 21048 8838
rect 20996 8774 21048 8780
rect 20916 8498 20944 8774
rect 20812 8492 20864 8498
rect 20812 8434 20864 8440
rect 20904 8492 20956 8498
rect 20904 8434 20956 8440
rect 20824 7449 20852 8434
rect 20810 7440 20866 7449
rect 20810 7375 20866 7384
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 20812 6112 20864 6118
rect 20732 6072 20812 6100
rect 20732 5642 20760 6072
rect 20812 6054 20864 6060
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 20720 5636 20772 5642
rect 20720 5578 20772 5584
rect 20588 5528 20668 5556
rect 20536 5510 20588 5516
rect 20548 5302 20576 5510
rect 20626 5400 20682 5409
rect 20626 5335 20628 5344
rect 20680 5335 20682 5344
rect 20628 5306 20680 5312
rect 20536 5296 20588 5302
rect 20536 5238 20588 5244
rect 20536 5160 20588 5166
rect 20536 5102 20588 5108
rect 20626 5128 20682 5137
rect 20548 4758 20576 5102
rect 20626 5063 20682 5072
rect 20536 4752 20588 4758
rect 20536 4694 20588 4700
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 20444 4004 20496 4010
rect 20444 3946 20496 3952
rect 20260 3936 20312 3942
rect 20312 3896 20392 3924
rect 20260 3878 20312 3884
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 20272 3398 20300 3470
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 20128 2604 20208 2632
rect 20076 2586 20128 2592
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 20076 2508 20128 2514
rect 20076 2450 20128 2456
rect 20088 800 20116 2450
rect 20364 1970 20392 3896
rect 20456 2854 20484 3946
rect 20548 3942 20576 4558
rect 20640 4486 20668 5063
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20640 3126 20668 4422
rect 20628 3120 20680 3126
rect 20628 3062 20680 3068
rect 20444 2848 20496 2854
rect 20444 2790 20496 2796
rect 20628 2576 20680 2582
rect 20628 2518 20680 2524
rect 20352 1964 20404 1970
rect 20352 1906 20404 1912
rect 20640 800 20668 2518
rect 20732 2378 20760 5578
rect 20824 5370 20852 5850
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20824 5030 20852 5306
rect 20812 5024 20864 5030
rect 20812 4966 20864 4972
rect 20916 3738 20944 7346
rect 21008 6361 21036 8774
rect 21088 8356 21140 8362
rect 21088 8298 21140 8304
rect 20994 6352 21050 6361
rect 20994 6287 21050 6296
rect 20994 5944 21050 5953
rect 20994 5879 20996 5888
rect 21048 5879 21050 5888
rect 20996 5850 21048 5856
rect 20996 5024 21048 5030
rect 20996 4966 21048 4972
rect 20904 3732 20956 3738
rect 20904 3674 20956 3680
rect 21008 3398 21036 4966
rect 21100 3738 21128 8298
rect 21192 7002 21220 10503
rect 21284 9674 21312 10628
rect 21364 10610 21416 10616
rect 21284 9646 21496 9674
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 21180 6996 21232 7002
rect 21180 6938 21232 6944
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 21088 3732 21140 3738
rect 21088 3674 21140 3680
rect 20996 3392 21048 3398
rect 20996 3334 21048 3340
rect 21008 3126 21036 3334
rect 20996 3120 21048 3126
rect 20996 3062 21048 3068
rect 20812 2984 20864 2990
rect 21008 2961 21036 3062
rect 20812 2926 20864 2932
rect 20994 2952 21050 2961
rect 20824 2446 20852 2926
rect 20904 2916 20956 2922
rect 21100 2922 21128 3674
rect 21192 3058 21220 5646
rect 21284 3738 21312 9522
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 21376 6497 21404 9318
rect 21362 6488 21418 6497
rect 21362 6423 21418 6432
rect 21362 5808 21418 5817
rect 21362 5743 21418 5752
rect 21272 3732 21324 3738
rect 21272 3674 21324 3680
rect 21180 3052 21232 3058
rect 21180 2994 21232 3000
rect 20994 2887 21050 2896
rect 21088 2916 21140 2922
rect 20904 2858 20956 2864
rect 20916 2650 20944 2858
rect 20904 2644 20956 2650
rect 20904 2586 20956 2592
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 21008 2378 21036 2887
rect 21088 2858 21140 2864
rect 21376 2854 21404 5743
rect 21468 3754 21496 9646
rect 21560 9330 21588 12124
rect 21730 12064 21786 12073
rect 21730 11999 21786 12008
rect 21640 11688 21692 11694
rect 21640 11630 21692 11636
rect 21652 11354 21680 11630
rect 21640 11348 21692 11354
rect 21640 11290 21692 11296
rect 21560 9302 21680 9330
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 21560 8906 21588 9114
rect 21652 9110 21680 9302
rect 21640 9104 21692 9110
rect 21638 9072 21640 9081
rect 21692 9072 21694 9081
rect 21638 9007 21694 9016
rect 21548 8900 21600 8906
rect 21548 8842 21600 8848
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 21560 7478 21588 7686
rect 21548 7472 21600 7478
rect 21548 7414 21600 7420
rect 21546 7304 21602 7313
rect 21546 7239 21602 7248
rect 21560 4486 21588 7239
rect 21652 6866 21680 8570
rect 21744 7721 21772 11999
rect 21730 7712 21786 7721
rect 21730 7647 21786 7656
rect 21730 7304 21786 7313
rect 21730 7239 21786 7248
rect 21640 6860 21692 6866
rect 21640 6802 21692 6808
rect 21640 6384 21692 6390
rect 21744 6372 21772 7239
rect 21836 6730 21864 12922
rect 21928 12238 21956 13262
rect 22020 12986 22048 13903
rect 22112 13734 22140 14214
rect 22190 14175 22246 14184
rect 22204 13870 22232 14175
rect 22192 13864 22244 13870
rect 22296 13841 22324 14282
rect 22192 13806 22244 13812
rect 22282 13832 22338 13841
rect 22282 13767 22338 13776
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22112 13462 22140 13670
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22100 13456 22152 13462
rect 22100 13398 22152 13404
rect 22098 13288 22154 13297
rect 22098 13223 22154 13232
rect 22112 13190 22140 13223
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 22008 12980 22060 12986
rect 22008 12922 22060 12928
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 21916 12232 21968 12238
rect 21916 12174 21968 12180
rect 21928 11218 21956 12174
rect 22008 11892 22060 11898
rect 22008 11834 22060 11840
rect 22020 11762 22048 11834
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 22006 11656 22062 11665
rect 22006 11591 22062 11600
rect 21916 11212 21968 11218
rect 21916 11154 21968 11160
rect 21916 10668 21968 10674
rect 21916 10610 21968 10616
rect 21928 10169 21956 10610
rect 21914 10160 21970 10169
rect 21914 10095 21970 10104
rect 21916 9104 21968 9110
rect 21916 9046 21968 9052
rect 21928 8838 21956 9046
rect 21916 8832 21968 8838
rect 21916 8774 21968 8780
rect 22020 8650 22048 11591
rect 22112 9586 22140 12582
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 21928 8622 22048 8650
rect 21928 7834 21956 8622
rect 22008 8084 22060 8090
rect 22008 8026 22060 8032
rect 22020 7993 22048 8026
rect 22006 7984 22062 7993
rect 22204 7970 22232 13466
rect 22296 13190 22324 13767
rect 22284 13184 22336 13190
rect 22284 13126 22336 13132
rect 22388 12986 22416 18566
rect 22376 12980 22428 12986
rect 22376 12922 22428 12928
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 22296 12374 22324 12786
rect 22284 12368 22336 12374
rect 22284 12310 22336 12316
rect 22284 12232 22336 12238
rect 22284 12174 22336 12180
rect 22296 11762 22324 12174
rect 22284 11756 22336 11762
rect 22284 11698 22336 11704
rect 22284 11552 22336 11558
rect 22284 11494 22336 11500
rect 22006 7919 22062 7928
rect 22112 7942 22232 7970
rect 21928 7806 22048 7834
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 21824 6724 21876 6730
rect 21824 6666 21876 6672
rect 21692 6344 21772 6372
rect 21640 6326 21692 6332
rect 21652 5234 21680 6326
rect 21928 6066 21956 7686
rect 22020 6662 22048 7806
rect 22008 6656 22060 6662
rect 22008 6598 22060 6604
rect 22020 6322 22048 6598
rect 22008 6316 22060 6322
rect 22008 6258 22060 6264
rect 22112 6202 22140 7942
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 22204 6798 22232 7822
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 22204 6322 22232 6734
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 21744 6038 21956 6066
rect 22020 6174 22140 6202
rect 21640 5228 21692 5234
rect 21640 5170 21692 5176
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21744 4146 21772 6038
rect 21916 5908 21968 5914
rect 21916 5850 21968 5856
rect 21822 5672 21878 5681
rect 21822 5607 21824 5616
rect 21876 5607 21878 5616
rect 21824 5578 21876 5584
rect 21928 5409 21956 5850
rect 21914 5400 21970 5409
rect 21914 5335 21916 5344
rect 21968 5335 21970 5344
rect 21916 5306 21968 5312
rect 21928 5275 21956 5306
rect 21824 5024 21876 5030
rect 21824 4966 21876 4972
rect 21836 4554 21864 4966
rect 22020 4604 22048 6174
rect 22100 6112 22152 6118
rect 22100 6054 22152 6060
rect 22112 5642 22140 6054
rect 22100 5636 22152 5642
rect 22100 5578 22152 5584
rect 22204 5522 22232 6258
rect 22296 6089 22324 11494
rect 22480 11082 22508 22918
rect 22572 22642 22600 23258
rect 22664 23202 22692 26438
rect 22744 26240 22796 26246
rect 22744 26182 22796 26188
rect 22756 25974 22784 26182
rect 22744 25968 22796 25974
rect 22744 25910 22796 25916
rect 22744 25424 22796 25430
rect 22744 25366 22796 25372
rect 22756 25294 22784 25366
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 22756 24410 22784 25230
rect 22744 24404 22796 24410
rect 22744 24346 22796 24352
rect 22744 24268 22796 24274
rect 22744 24210 22796 24216
rect 22756 23322 22784 24210
rect 22848 24138 22876 26930
rect 22836 24132 22888 24138
rect 22836 24074 22888 24080
rect 22834 23352 22890 23361
rect 22744 23316 22796 23322
rect 22834 23287 22836 23296
rect 22744 23258 22796 23264
rect 22888 23287 22890 23296
rect 22836 23258 22888 23264
rect 22664 23174 22876 23202
rect 22744 22772 22796 22778
rect 22744 22714 22796 22720
rect 22652 22704 22704 22710
rect 22652 22646 22704 22652
rect 22560 22636 22612 22642
rect 22560 22578 22612 22584
rect 22560 22500 22612 22506
rect 22560 22442 22612 22448
rect 22572 21554 22600 22442
rect 22664 21622 22692 22646
rect 22652 21616 22704 21622
rect 22652 21558 22704 21564
rect 22560 21548 22612 21554
rect 22560 21490 22612 21496
rect 22572 20942 22600 21490
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22560 19984 22612 19990
rect 22560 19926 22612 19932
rect 22572 14958 22600 19926
rect 22652 19848 22704 19854
rect 22652 19790 22704 19796
rect 22664 19553 22692 19790
rect 22650 19544 22706 19553
rect 22650 19479 22706 19488
rect 22650 19408 22706 19417
rect 22650 19343 22652 19352
rect 22704 19343 22706 19352
rect 22652 19314 22704 19320
rect 22652 19236 22704 19242
rect 22652 19178 22704 19184
rect 22664 17202 22692 19178
rect 22652 17196 22704 17202
rect 22652 17138 22704 17144
rect 22652 16720 22704 16726
rect 22652 16662 22704 16668
rect 22560 14952 22612 14958
rect 22560 14894 22612 14900
rect 22664 14770 22692 16662
rect 22572 14742 22692 14770
rect 22468 11076 22520 11082
rect 22468 11018 22520 11024
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 22388 9625 22416 10746
rect 22468 10260 22520 10266
rect 22468 10202 22520 10208
rect 22374 9616 22430 9625
rect 22374 9551 22430 9560
rect 22376 8968 22428 8974
rect 22376 8910 22428 8916
rect 22282 6080 22338 6089
rect 22282 6015 22338 6024
rect 22284 5772 22336 5778
rect 22284 5714 22336 5720
rect 22112 5494 22232 5522
rect 22112 4758 22140 5494
rect 22296 5273 22324 5714
rect 22282 5264 22338 5273
rect 22282 5199 22338 5208
rect 22388 5114 22416 8910
rect 22480 7274 22508 10202
rect 22468 7268 22520 7274
rect 22468 7210 22520 7216
rect 22572 6458 22600 14742
rect 22650 14648 22706 14657
rect 22650 14583 22706 14592
rect 22664 14385 22692 14583
rect 22650 14376 22706 14385
rect 22650 14311 22706 14320
rect 22664 13938 22692 14311
rect 22652 13932 22704 13938
rect 22652 13874 22704 13880
rect 22650 13832 22706 13841
rect 22650 13767 22706 13776
rect 22664 12850 22692 13767
rect 22652 12844 22704 12850
rect 22652 12786 22704 12792
rect 22756 11150 22784 22714
rect 22848 19417 22876 23174
rect 22834 19408 22890 19417
rect 22834 19343 22890 19352
rect 22940 17592 22968 28494
rect 27068 28416 27120 28422
rect 27068 28358 27120 28364
rect 23296 28076 23348 28082
rect 23296 28018 23348 28024
rect 26884 28076 26936 28082
rect 26884 28018 26936 28024
rect 23308 27878 23336 28018
rect 25872 27940 25924 27946
rect 25872 27882 25924 27888
rect 23296 27872 23348 27878
rect 23296 27814 23348 27820
rect 23848 27872 23900 27878
rect 23848 27814 23900 27820
rect 23413 27772 23721 27792
rect 23413 27770 23419 27772
rect 23475 27770 23499 27772
rect 23555 27770 23579 27772
rect 23635 27770 23659 27772
rect 23715 27770 23721 27772
rect 23475 27718 23477 27770
rect 23657 27718 23659 27770
rect 23413 27716 23419 27718
rect 23475 27716 23499 27718
rect 23555 27716 23579 27718
rect 23635 27716 23659 27718
rect 23715 27716 23721 27718
rect 23413 27696 23721 27716
rect 23860 27713 23888 27814
rect 23846 27704 23902 27713
rect 23846 27639 23902 27648
rect 25228 27600 25280 27606
rect 25228 27542 25280 27548
rect 23204 27532 23256 27538
rect 23204 27474 23256 27480
rect 23020 27328 23072 27334
rect 23020 27270 23072 27276
rect 23032 25158 23060 27270
rect 23112 26784 23164 26790
rect 23112 26726 23164 26732
rect 23020 25152 23072 25158
rect 23020 25094 23072 25100
rect 23032 19666 23060 25094
rect 23124 23730 23152 26726
rect 23216 26353 23244 27474
rect 23756 27464 23808 27470
rect 23756 27406 23808 27412
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 23413 26684 23721 26704
rect 23413 26682 23419 26684
rect 23475 26682 23499 26684
rect 23555 26682 23579 26684
rect 23635 26682 23659 26684
rect 23715 26682 23721 26684
rect 23475 26630 23477 26682
rect 23657 26630 23659 26682
rect 23413 26628 23419 26630
rect 23475 26628 23499 26630
rect 23555 26628 23579 26630
rect 23635 26628 23659 26630
rect 23715 26628 23721 26630
rect 23413 26608 23721 26628
rect 23202 26344 23258 26353
rect 23202 26279 23258 26288
rect 23202 25936 23258 25945
rect 23202 25871 23204 25880
rect 23256 25871 23258 25880
rect 23296 25900 23348 25906
rect 23204 25842 23256 25848
rect 23296 25842 23348 25848
rect 23216 24886 23244 25842
rect 23204 24880 23256 24886
rect 23204 24822 23256 24828
rect 23204 24744 23256 24750
rect 23204 24686 23256 24692
rect 23216 23866 23244 24686
rect 23308 24410 23336 25842
rect 23413 25596 23721 25616
rect 23413 25594 23419 25596
rect 23475 25594 23499 25596
rect 23555 25594 23579 25596
rect 23635 25594 23659 25596
rect 23715 25594 23721 25596
rect 23475 25542 23477 25594
rect 23657 25542 23659 25594
rect 23413 25540 23419 25542
rect 23475 25540 23499 25542
rect 23555 25540 23579 25542
rect 23635 25540 23659 25542
rect 23715 25540 23721 25542
rect 23413 25520 23721 25540
rect 23413 24508 23721 24528
rect 23413 24506 23419 24508
rect 23475 24506 23499 24508
rect 23555 24506 23579 24508
rect 23635 24506 23659 24508
rect 23715 24506 23721 24508
rect 23475 24454 23477 24506
rect 23657 24454 23659 24506
rect 23413 24452 23419 24454
rect 23475 24452 23499 24454
rect 23555 24452 23579 24454
rect 23635 24452 23659 24454
rect 23715 24452 23721 24454
rect 23413 24432 23721 24452
rect 23296 24404 23348 24410
rect 23296 24346 23348 24352
rect 23388 24336 23440 24342
rect 23388 24278 23440 24284
rect 23400 24154 23428 24278
rect 23308 24126 23428 24154
rect 23204 23860 23256 23866
rect 23204 23802 23256 23808
rect 23308 23746 23336 24126
rect 23388 24064 23440 24070
rect 23388 24006 23440 24012
rect 23112 23724 23164 23730
rect 23112 23666 23164 23672
rect 23216 23718 23336 23746
rect 23400 23730 23428 24006
rect 23388 23724 23440 23730
rect 23124 23118 23152 23666
rect 23112 23112 23164 23118
rect 23112 23054 23164 23060
rect 23124 22506 23152 23054
rect 23112 22500 23164 22506
rect 23112 22442 23164 22448
rect 23112 21888 23164 21894
rect 23112 21830 23164 21836
rect 23124 21622 23152 21830
rect 23112 21616 23164 21622
rect 23112 21558 23164 21564
rect 23216 21418 23244 23718
rect 23388 23666 23440 23672
rect 23296 23656 23348 23662
rect 23296 23598 23348 23604
rect 23308 23186 23336 23598
rect 23413 23420 23721 23440
rect 23413 23418 23419 23420
rect 23475 23418 23499 23420
rect 23555 23418 23579 23420
rect 23635 23418 23659 23420
rect 23715 23418 23721 23420
rect 23475 23366 23477 23418
rect 23657 23366 23659 23418
rect 23413 23364 23419 23366
rect 23475 23364 23499 23366
rect 23555 23364 23579 23366
rect 23635 23364 23659 23366
rect 23715 23364 23721 23366
rect 23413 23344 23721 23364
rect 23386 23216 23442 23225
rect 23296 23180 23348 23186
rect 23386 23151 23442 23160
rect 23296 23122 23348 23128
rect 23308 22438 23336 23122
rect 23400 23050 23428 23151
rect 23388 23044 23440 23050
rect 23388 22986 23440 22992
rect 23400 22574 23428 22986
rect 23388 22568 23440 22574
rect 23388 22510 23440 22516
rect 23296 22432 23348 22438
rect 23296 22374 23348 22380
rect 23204 21412 23256 21418
rect 23204 21354 23256 21360
rect 23112 21072 23164 21078
rect 23112 21014 23164 21020
rect 23124 19922 23152 21014
rect 23308 21010 23336 22374
rect 23413 22332 23721 22352
rect 23413 22330 23419 22332
rect 23475 22330 23499 22332
rect 23555 22330 23579 22332
rect 23635 22330 23659 22332
rect 23715 22330 23721 22332
rect 23475 22278 23477 22330
rect 23657 22278 23659 22330
rect 23413 22276 23419 22278
rect 23475 22276 23499 22278
rect 23555 22276 23579 22278
rect 23635 22276 23659 22278
rect 23715 22276 23721 22278
rect 23413 22256 23721 22276
rect 23480 22160 23532 22166
rect 23480 22102 23532 22108
rect 23388 22092 23440 22098
rect 23388 22034 23440 22040
rect 23400 21690 23428 22034
rect 23388 21684 23440 21690
rect 23388 21626 23440 21632
rect 23388 21548 23440 21554
rect 23492 21536 23520 22102
rect 23572 22024 23624 22030
rect 23572 21966 23624 21972
rect 23440 21508 23520 21536
rect 23388 21490 23440 21496
rect 23584 21486 23612 21966
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 23676 21690 23704 21830
rect 23664 21684 23716 21690
rect 23664 21626 23716 21632
rect 23572 21480 23624 21486
rect 23572 21422 23624 21428
rect 23413 21244 23721 21264
rect 23413 21242 23419 21244
rect 23475 21242 23499 21244
rect 23555 21242 23579 21244
rect 23635 21242 23659 21244
rect 23715 21242 23721 21244
rect 23475 21190 23477 21242
rect 23657 21190 23659 21242
rect 23413 21188 23419 21190
rect 23475 21188 23499 21190
rect 23555 21188 23579 21190
rect 23635 21188 23659 21190
rect 23715 21188 23721 21190
rect 23413 21168 23721 21188
rect 23768 21146 23796 27406
rect 24216 27396 24268 27402
rect 24216 27338 24268 27344
rect 24308 27396 24360 27402
rect 24308 27338 24360 27344
rect 23940 27328 23992 27334
rect 23940 27270 23992 27276
rect 23848 26988 23900 26994
rect 23848 26930 23900 26936
rect 23860 26081 23888 26930
rect 23846 26072 23902 26081
rect 23846 26007 23902 26016
rect 23848 24744 23900 24750
rect 23848 24686 23900 24692
rect 23860 22642 23888 24686
rect 23848 22636 23900 22642
rect 23848 22578 23900 22584
rect 23860 22166 23888 22578
rect 23848 22160 23900 22166
rect 23848 22102 23900 22108
rect 23848 21344 23900 21350
rect 23848 21286 23900 21292
rect 23756 21140 23808 21146
rect 23756 21082 23808 21088
rect 23296 21004 23348 21010
rect 23296 20946 23348 20952
rect 23756 21004 23808 21010
rect 23756 20946 23808 20952
rect 23413 20156 23721 20176
rect 23413 20154 23419 20156
rect 23475 20154 23499 20156
rect 23555 20154 23579 20156
rect 23635 20154 23659 20156
rect 23715 20154 23721 20156
rect 23475 20102 23477 20154
rect 23657 20102 23659 20154
rect 23413 20100 23419 20102
rect 23475 20100 23499 20102
rect 23555 20100 23579 20102
rect 23635 20100 23659 20102
rect 23715 20100 23721 20102
rect 23413 20080 23721 20100
rect 23112 19916 23164 19922
rect 23112 19858 23164 19864
rect 23572 19916 23624 19922
rect 23572 19858 23624 19864
rect 23296 19712 23348 19718
rect 23032 19638 23152 19666
rect 23296 19654 23348 19660
rect 23020 19508 23072 19514
rect 23020 19450 23072 19456
rect 22848 17564 22968 17592
rect 22848 11558 22876 17564
rect 23032 17513 23060 19450
rect 23124 19242 23152 19638
rect 23204 19440 23256 19446
rect 23204 19382 23256 19388
rect 23112 19236 23164 19242
rect 23112 19178 23164 19184
rect 23216 19145 23244 19382
rect 23308 19378 23336 19654
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 23584 19242 23612 19858
rect 23664 19304 23716 19310
rect 23662 19272 23664 19281
rect 23716 19272 23718 19281
rect 23572 19236 23624 19242
rect 23662 19207 23718 19216
rect 23572 19178 23624 19184
rect 23202 19136 23258 19145
rect 23202 19071 23258 19080
rect 23413 19068 23721 19088
rect 23413 19066 23419 19068
rect 23475 19066 23499 19068
rect 23555 19066 23579 19068
rect 23635 19066 23659 19068
rect 23715 19066 23721 19068
rect 23475 19014 23477 19066
rect 23657 19014 23659 19066
rect 23413 19012 23419 19014
rect 23475 19012 23499 19014
rect 23555 19012 23579 19014
rect 23635 19012 23659 19014
rect 23715 19012 23721 19014
rect 23413 18992 23721 19012
rect 23204 18828 23256 18834
rect 23204 18770 23256 18776
rect 23112 18624 23164 18630
rect 23112 18566 23164 18572
rect 23124 17610 23152 18566
rect 23216 17882 23244 18770
rect 23413 17980 23721 18000
rect 23413 17978 23419 17980
rect 23475 17978 23499 17980
rect 23555 17978 23579 17980
rect 23635 17978 23659 17980
rect 23715 17978 23721 17980
rect 23475 17926 23477 17978
rect 23657 17926 23659 17978
rect 23413 17924 23419 17926
rect 23475 17924 23499 17926
rect 23555 17924 23579 17926
rect 23635 17924 23659 17926
rect 23715 17924 23721 17926
rect 23413 17904 23721 17924
rect 23204 17876 23256 17882
rect 23204 17818 23256 17824
rect 23112 17604 23164 17610
rect 23112 17546 23164 17552
rect 23296 17536 23348 17542
rect 23018 17504 23074 17513
rect 23296 17478 23348 17484
rect 23018 17439 23074 17448
rect 23020 17196 23072 17202
rect 23020 17138 23072 17144
rect 23204 17196 23256 17202
rect 23204 17138 23256 17144
rect 23032 16969 23060 17138
rect 23018 16960 23074 16969
rect 23018 16895 23074 16904
rect 23032 16658 23060 16895
rect 22928 16652 22980 16658
rect 22928 16594 22980 16600
rect 23020 16652 23072 16658
rect 23020 16594 23072 16600
rect 22940 16182 22968 16594
rect 23216 16522 23244 17138
rect 23308 17105 23336 17478
rect 23664 17196 23716 17202
rect 23768 17184 23796 20946
rect 23860 20942 23888 21286
rect 23848 20936 23900 20942
rect 23848 20878 23900 20884
rect 23848 20460 23900 20466
rect 23848 20402 23900 20408
rect 23860 19378 23888 20402
rect 23848 19372 23900 19378
rect 23848 19314 23900 19320
rect 23848 19236 23900 19242
rect 23848 19178 23900 19184
rect 23716 17156 23796 17184
rect 23860 18034 23888 19178
rect 23952 18358 23980 27270
rect 24228 26994 24256 27338
rect 24216 26988 24268 26994
rect 24216 26930 24268 26936
rect 24216 26784 24268 26790
rect 24216 26726 24268 26732
rect 24032 26240 24084 26246
rect 24032 26182 24084 26188
rect 24044 26042 24072 26182
rect 24032 26036 24084 26042
rect 24032 25978 24084 25984
rect 24044 25242 24072 25978
rect 24124 25968 24176 25974
rect 24124 25910 24176 25916
rect 24136 25362 24164 25910
rect 24228 25838 24256 26726
rect 24216 25832 24268 25838
rect 24216 25774 24268 25780
rect 24124 25356 24176 25362
rect 24124 25298 24176 25304
rect 24044 25214 24164 25242
rect 24136 24138 24164 25214
rect 24124 24132 24176 24138
rect 24124 24074 24176 24080
rect 24032 24064 24084 24070
rect 24032 24006 24084 24012
rect 24044 21978 24072 24006
rect 24136 22778 24164 24074
rect 24216 22976 24268 22982
rect 24216 22918 24268 22924
rect 24124 22772 24176 22778
rect 24124 22714 24176 22720
rect 24044 21950 24164 21978
rect 24032 21888 24084 21894
rect 24032 21830 24084 21836
rect 24044 20602 24072 21830
rect 24136 21010 24164 21950
rect 24124 21004 24176 21010
rect 24124 20946 24176 20952
rect 24228 20890 24256 22918
rect 24136 20862 24256 20890
rect 24032 20596 24084 20602
rect 24032 20538 24084 20544
rect 24136 20482 24164 20862
rect 24216 20800 24268 20806
rect 24216 20742 24268 20748
rect 24044 20454 24164 20482
rect 24044 19258 24072 20454
rect 24228 20398 24256 20742
rect 24216 20392 24268 20398
rect 24216 20334 24268 20340
rect 24124 20256 24176 20262
rect 24124 20198 24176 20204
rect 24136 19446 24164 20198
rect 24320 20058 24348 27338
rect 24492 27328 24544 27334
rect 24492 27270 24544 27276
rect 24504 26314 24532 27270
rect 24492 26308 24544 26314
rect 24492 26250 24544 26256
rect 24596 26042 24624 27406
rect 25136 27328 25188 27334
rect 25136 27270 25188 27276
rect 24584 26036 24636 26042
rect 24584 25978 24636 25984
rect 24952 25900 25004 25906
rect 24952 25842 25004 25848
rect 24860 25696 24912 25702
rect 24860 25638 24912 25644
rect 24400 25288 24452 25294
rect 24400 25230 24452 25236
rect 24584 25288 24636 25294
rect 24584 25230 24636 25236
rect 24412 24818 24440 25230
rect 24400 24812 24452 24818
rect 24400 24754 24452 24760
rect 24492 24200 24544 24206
rect 24492 24142 24544 24148
rect 24400 23656 24452 23662
rect 24400 23598 24452 23604
rect 24412 22953 24440 23598
rect 24398 22944 24454 22953
rect 24398 22879 24454 22888
rect 24400 22772 24452 22778
rect 24400 22714 24452 22720
rect 24412 21146 24440 22714
rect 24400 21140 24452 21146
rect 24400 21082 24452 21088
rect 24400 21004 24452 21010
rect 24400 20946 24452 20952
rect 24308 20052 24360 20058
rect 24308 19994 24360 20000
rect 24216 19848 24268 19854
rect 24216 19790 24268 19796
rect 24308 19848 24360 19854
rect 24308 19790 24360 19796
rect 24124 19440 24176 19446
rect 24124 19382 24176 19388
rect 24044 19230 24164 19258
rect 24032 19168 24084 19174
rect 24032 19110 24084 19116
rect 23940 18352 23992 18358
rect 23940 18294 23992 18300
rect 23940 18080 23992 18086
rect 23860 18028 23940 18034
rect 23860 18022 23992 18028
rect 23860 18006 23980 18022
rect 23664 17138 23716 17144
rect 23294 17096 23350 17105
rect 23294 17031 23350 17040
rect 23296 16992 23348 16998
rect 23296 16934 23348 16940
rect 23204 16516 23256 16522
rect 23204 16458 23256 16464
rect 23018 16416 23074 16425
rect 23018 16351 23074 16360
rect 22928 16176 22980 16182
rect 22928 16118 22980 16124
rect 22940 15638 22968 16118
rect 22928 15632 22980 15638
rect 22928 15574 22980 15580
rect 22928 14816 22980 14822
rect 22928 14758 22980 14764
rect 22940 14278 22968 14758
rect 22928 14272 22980 14278
rect 22928 14214 22980 14220
rect 23032 13530 23060 16351
rect 23204 16108 23256 16114
rect 23204 16050 23256 16056
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 23124 15201 23152 15846
rect 23216 15706 23244 16050
rect 23204 15700 23256 15706
rect 23204 15642 23256 15648
rect 23204 15564 23256 15570
rect 23204 15506 23256 15512
rect 23216 15473 23244 15506
rect 23308 15502 23336 16934
rect 23413 16892 23721 16912
rect 23413 16890 23419 16892
rect 23475 16890 23499 16892
rect 23555 16890 23579 16892
rect 23635 16890 23659 16892
rect 23715 16890 23721 16892
rect 23475 16838 23477 16890
rect 23657 16838 23659 16890
rect 23413 16836 23419 16838
rect 23475 16836 23499 16838
rect 23555 16836 23579 16838
rect 23635 16836 23659 16838
rect 23715 16836 23721 16838
rect 23413 16816 23721 16836
rect 23756 16244 23808 16250
rect 23756 16186 23808 16192
rect 23768 16046 23796 16186
rect 23756 16040 23808 16046
rect 23756 15982 23808 15988
rect 23413 15804 23721 15824
rect 23413 15802 23419 15804
rect 23475 15802 23499 15804
rect 23555 15802 23579 15804
rect 23635 15802 23659 15804
rect 23715 15802 23721 15804
rect 23475 15750 23477 15802
rect 23657 15750 23659 15802
rect 23413 15748 23419 15750
rect 23475 15748 23499 15750
rect 23555 15748 23579 15750
rect 23635 15748 23659 15750
rect 23715 15748 23721 15750
rect 23413 15728 23721 15748
rect 23664 15564 23716 15570
rect 23664 15506 23716 15512
rect 23296 15496 23348 15502
rect 23202 15464 23258 15473
rect 23296 15438 23348 15444
rect 23202 15399 23258 15408
rect 23676 15201 23704 15506
rect 23110 15192 23166 15201
rect 23110 15127 23166 15136
rect 23662 15192 23718 15201
rect 23662 15127 23718 15136
rect 23112 15020 23164 15026
rect 23112 14962 23164 14968
rect 23124 14618 23152 14962
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 23478 14920 23534 14929
rect 23204 14884 23256 14890
rect 23204 14826 23256 14832
rect 23216 14657 23244 14826
rect 23202 14648 23258 14657
rect 23112 14612 23164 14618
rect 23202 14583 23258 14592
rect 23112 14554 23164 14560
rect 23308 14482 23336 14894
rect 23478 14855 23480 14864
rect 23532 14855 23534 14864
rect 23480 14826 23532 14832
rect 23413 14716 23721 14736
rect 23413 14714 23419 14716
rect 23475 14714 23499 14716
rect 23555 14714 23579 14716
rect 23635 14714 23659 14716
rect 23715 14714 23721 14716
rect 23475 14662 23477 14714
rect 23657 14662 23659 14714
rect 23413 14660 23419 14662
rect 23475 14660 23499 14662
rect 23555 14660 23579 14662
rect 23635 14660 23659 14662
rect 23715 14660 23721 14662
rect 23413 14640 23721 14660
rect 23662 14512 23718 14521
rect 23296 14476 23348 14482
rect 23768 14482 23796 15982
rect 23860 15502 23888 18006
rect 24044 17898 24072 19110
rect 23952 17882 24072 17898
rect 23952 17876 24084 17882
rect 23952 17870 24032 17876
rect 23952 16130 23980 17870
rect 24032 17818 24084 17824
rect 24044 17787 24072 17818
rect 24032 17128 24084 17134
rect 24032 17070 24084 17076
rect 24044 16726 24072 17070
rect 24032 16720 24084 16726
rect 24032 16662 24084 16668
rect 24044 16250 24072 16662
rect 24136 16454 24164 19230
rect 24228 19174 24256 19790
rect 24216 19168 24268 19174
rect 24216 19110 24268 19116
rect 24320 18850 24348 19790
rect 24412 19334 24440 20946
rect 24504 19854 24532 24142
rect 24596 23322 24624 25230
rect 24676 25220 24728 25226
rect 24676 25162 24728 25168
rect 24584 23316 24636 23322
rect 24584 23258 24636 23264
rect 24688 23168 24716 25162
rect 24768 24812 24820 24818
rect 24768 24754 24820 24760
rect 24780 23866 24808 24754
rect 24768 23860 24820 23866
rect 24768 23802 24820 23808
rect 24768 23724 24820 23730
rect 24768 23666 24820 23672
rect 24596 23140 24716 23168
rect 24596 22982 24624 23140
rect 24780 23118 24808 23666
rect 24768 23112 24820 23118
rect 24688 23072 24768 23100
rect 24584 22976 24636 22982
rect 24584 22918 24636 22924
rect 24688 21962 24716 23072
rect 24768 23054 24820 23060
rect 24676 21956 24728 21962
rect 24676 21898 24728 21904
rect 24768 21888 24820 21894
rect 24768 21830 24820 21836
rect 24780 21690 24808 21830
rect 24768 21684 24820 21690
rect 24768 21626 24820 21632
rect 24872 21622 24900 25638
rect 24964 25498 24992 25842
rect 24952 25492 25004 25498
rect 24952 25434 25004 25440
rect 24952 25288 25004 25294
rect 24952 25230 25004 25236
rect 24964 24818 24992 25230
rect 24952 24812 25004 24818
rect 24952 24754 25004 24760
rect 25044 24744 25096 24750
rect 25044 24686 25096 24692
rect 24952 24608 25004 24614
rect 24952 24550 25004 24556
rect 24584 21616 24636 21622
rect 24584 21558 24636 21564
rect 24860 21616 24912 21622
rect 24860 21558 24912 21564
rect 24492 19848 24544 19854
rect 24492 19790 24544 19796
rect 24490 19544 24546 19553
rect 24490 19479 24546 19488
rect 24504 19446 24532 19479
rect 24492 19440 24544 19446
rect 24492 19382 24544 19388
rect 24412 19306 24532 19334
rect 24228 18822 24348 18850
rect 24228 17785 24256 18822
rect 24308 18760 24360 18766
rect 24308 18702 24360 18708
rect 24214 17776 24270 17785
rect 24214 17711 24270 17720
rect 24216 17604 24268 17610
rect 24216 17546 24268 17552
rect 24228 17338 24256 17546
rect 24216 17332 24268 17338
rect 24216 17274 24268 17280
rect 24320 17134 24348 18702
rect 24308 17128 24360 17134
rect 24308 17070 24360 17076
rect 24216 16652 24268 16658
rect 24216 16594 24268 16600
rect 24124 16448 24176 16454
rect 24124 16390 24176 16396
rect 24032 16244 24084 16250
rect 24032 16186 24084 16192
rect 23952 16102 24072 16130
rect 23848 15496 23900 15502
rect 23848 15438 23900 15444
rect 23848 15360 23900 15366
rect 23848 15302 23900 15308
rect 23662 14447 23718 14456
rect 23756 14476 23808 14482
rect 23296 14418 23348 14424
rect 23110 14376 23166 14385
rect 23676 14346 23704 14447
rect 23756 14418 23808 14424
rect 23110 14311 23166 14320
rect 23664 14340 23716 14346
rect 23124 13938 23152 14311
rect 23664 14282 23716 14288
rect 23478 13968 23534 13977
rect 23112 13932 23164 13938
rect 23112 13874 23164 13880
rect 23204 13932 23256 13938
rect 23478 13903 23534 13912
rect 23204 13874 23256 13880
rect 23112 13796 23164 13802
rect 23112 13738 23164 13744
rect 23020 13524 23072 13530
rect 23020 13466 23072 13472
rect 22928 12776 22980 12782
rect 22928 12718 22980 12724
rect 22940 12374 22968 12718
rect 23124 12434 23152 13738
rect 23032 12406 23152 12434
rect 22928 12368 22980 12374
rect 22928 12310 22980 12316
rect 22836 11552 22888 11558
rect 22836 11494 22888 11500
rect 22744 11144 22796 11150
rect 22744 11086 22796 11092
rect 22756 9994 22784 11086
rect 22940 10674 22968 12310
rect 22928 10668 22980 10674
rect 22928 10610 22980 10616
rect 22836 10464 22888 10470
rect 22836 10406 22888 10412
rect 22744 9988 22796 9994
rect 22744 9930 22796 9936
rect 22652 9920 22704 9926
rect 22652 9862 22704 9868
rect 22664 6934 22692 9862
rect 22756 8566 22784 9930
rect 22744 8560 22796 8566
rect 22744 8502 22796 8508
rect 22744 8356 22796 8362
rect 22744 8298 22796 8304
rect 22652 6928 22704 6934
rect 22652 6870 22704 6876
rect 22560 6452 22612 6458
rect 22560 6394 22612 6400
rect 22650 6352 22706 6361
rect 22650 6287 22652 6296
rect 22704 6287 22706 6296
rect 22652 6258 22704 6264
rect 22466 5944 22522 5953
rect 22466 5879 22468 5888
rect 22520 5879 22522 5888
rect 22468 5850 22520 5856
rect 22652 5568 22704 5574
rect 22652 5510 22704 5516
rect 22468 5296 22520 5302
rect 22468 5238 22520 5244
rect 22204 5086 22416 5114
rect 22100 4752 22152 4758
rect 22100 4694 22152 4700
rect 22020 4576 22094 4604
rect 21824 4548 21876 4554
rect 22066 4536 22094 4576
rect 22066 4508 22140 4536
rect 21824 4490 21876 4496
rect 22112 4214 22140 4508
rect 22100 4208 22152 4214
rect 22100 4150 22152 4156
rect 21732 4140 21784 4146
rect 21732 4082 21784 4088
rect 22100 4072 22152 4078
rect 22100 4014 22152 4020
rect 21468 3726 21680 3754
rect 21456 3664 21508 3670
rect 21456 3606 21508 3612
rect 21468 2990 21496 3606
rect 21652 3194 21680 3726
rect 21732 3528 21784 3534
rect 21732 3470 21784 3476
rect 21640 3188 21692 3194
rect 21640 3130 21692 3136
rect 21456 2984 21508 2990
rect 21456 2926 21508 2932
rect 21364 2848 21416 2854
rect 21364 2790 21416 2796
rect 21744 2650 21772 3470
rect 22112 3058 22140 4014
rect 22100 3052 22152 3058
rect 22100 2994 22152 3000
rect 22204 2650 22232 5086
rect 22284 4684 22336 4690
rect 22284 4626 22336 4632
rect 22296 4078 22324 4626
rect 22480 4486 22508 5238
rect 22560 5228 22612 5234
rect 22560 5170 22612 5176
rect 22572 4729 22600 5170
rect 22558 4720 22614 4729
rect 22558 4655 22614 4664
rect 22560 4548 22612 4554
rect 22560 4490 22612 4496
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 22284 4072 22336 4078
rect 22284 4014 22336 4020
rect 22388 3482 22416 4082
rect 22296 3454 22416 3482
rect 22480 3466 22508 4422
rect 22572 4146 22600 4490
rect 22560 4140 22612 4146
rect 22560 4082 22612 4088
rect 22468 3460 22520 3466
rect 22296 2854 22324 3454
rect 22468 3402 22520 3408
rect 22376 3392 22428 3398
rect 22376 3334 22428 3340
rect 22388 3058 22416 3334
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 22284 2848 22336 2854
rect 22284 2790 22336 2796
rect 21732 2644 21784 2650
rect 21732 2586 21784 2592
rect 22192 2644 22244 2650
rect 22192 2586 22244 2592
rect 22664 2446 22692 5510
rect 22756 5166 22784 8298
rect 22848 5778 22876 10406
rect 22928 10260 22980 10266
rect 22928 10202 22980 10208
rect 22836 5772 22888 5778
rect 22836 5714 22888 5720
rect 22940 5302 22968 10202
rect 23032 8072 23060 12406
rect 23112 12096 23164 12102
rect 23112 12038 23164 12044
rect 23124 11762 23152 12038
rect 23112 11756 23164 11762
rect 23112 11698 23164 11704
rect 23216 11354 23244 13874
rect 23492 13870 23520 13903
rect 23480 13864 23532 13870
rect 23480 13806 23532 13812
rect 23413 13628 23721 13648
rect 23413 13626 23419 13628
rect 23475 13626 23499 13628
rect 23555 13626 23579 13628
rect 23635 13626 23659 13628
rect 23715 13626 23721 13628
rect 23475 13574 23477 13626
rect 23657 13574 23659 13626
rect 23413 13572 23419 13574
rect 23475 13572 23499 13574
rect 23555 13572 23579 13574
rect 23635 13572 23659 13574
rect 23715 13572 23721 13574
rect 23413 13552 23721 13572
rect 23480 13456 23532 13462
rect 23480 13398 23532 13404
rect 23296 13252 23348 13258
rect 23296 13194 23348 13200
rect 23308 12442 23336 13194
rect 23386 13152 23442 13161
rect 23386 13087 23442 13096
rect 23400 12782 23428 13087
rect 23492 12918 23520 13398
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23480 12912 23532 12918
rect 23480 12854 23532 12860
rect 23388 12776 23440 12782
rect 23388 12718 23440 12724
rect 23584 12714 23612 13330
rect 23756 13320 23808 13326
rect 23756 13262 23808 13268
rect 23768 12918 23796 13262
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 23572 12708 23624 12714
rect 23572 12650 23624 12656
rect 23413 12540 23721 12560
rect 23413 12538 23419 12540
rect 23475 12538 23499 12540
rect 23555 12538 23579 12540
rect 23635 12538 23659 12540
rect 23715 12538 23721 12540
rect 23475 12486 23477 12538
rect 23657 12486 23659 12538
rect 23413 12484 23419 12486
rect 23475 12484 23499 12486
rect 23555 12484 23579 12486
rect 23635 12484 23659 12486
rect 23715 12484 23721 12486
rect 23413 12464 23721 12484
rect 23296 12436 23348 12442
rect 23296 12378 23348 12384
rect 23296 11892 23348 11898
rect 23296 11834 23348 11840
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23308 11082 23336 11834
rect 23768 11830 23796 12854
rect 23860 12238 23888 15302
rect 24044 13297 24072 16102
rect 24228 15042 24256 16594
rect 24320 15706 24348 17070
rect 24400 16584 24452 16590
rect 24400 16526 24452 16532
rect 24412 16114 24440 16526
rect 24400 16108 24452 16114
rect 24400 16050 24452 16056
rect 24308 15700 24360 15706
rect 24308 15642 24360 15648
rect 24136 15014 24256 15042
rect 24400 15020 24452 15026
rect 24030 13288 24086 13297
rect 24030 13223 24086 13232
rect 24032 13184 24084 13190
rect 24032 13126 24084 13132
rect 23940 12844 23992 12850
rect 23940 12786 23992 12792
rect 23848 12232 23900 12238
rect 23848 12174 23900 12180
rect 23952 11898 23980 12786
rect 24044 12306 24072 13126
rect 24136 12753 24164 15014
rect 24400 14962 24452 14968
rect 24216 14816 24268 14822
rect 24216 14758 24268 14764
rect 24228 14414 24256 14758
rect 24216 14408 24268 14414
rect 24216 14350 24268 14356
rect 24308 14340 24360 14346
rect 24308 14282 24360 14288
rect 24216 14272 24268 14278
rect 24216 14214 24268 14220
rect 24228 14006 24256 14214
rect 24216 14000 24268 14006
rect 24214 13968 24216 13977
rect 24268 13968 24270 13977
rect 24214 13903 24270 13912
rect 24216 13864 24268 13870
rect 24216 13806 24268 13812
rect 24122 12744 24178 12753
rect 24122 12679 24178 12688
rect 24122 12472 24178 12481
rect 24122 12407 24178 12416
rect 24136 12374 24164 12407
rect 24124 12368 24176 12374
rect 24124 12310 24176 12316
rect 24032 12300 24084 12306
rect 24032 12242 24084 12248
rect 24032 12096 24084 12102
rect 24032 12038 24084 12044
rect 23940 11892 23992 11898
rect 23940 11834 23992 11840
rect 23756 11824 23808 11830
rect 23756 11766 23808 11772
rect 23754 11656 23810 11665
rect 23754 11591 23810 11600
rect 23413 11452 23721 11472
rect 23413 11450 23419 11452
rect 23475 11450 23499 11452
rect 23555 11450 23579 11452
rect 23635 11450 23659 11452
rect 23715 11450 23721 11452
rect 23475 11398 23477 11450
rect 23657 11398 23659 11450
rect 23413 11396 23419 11398
rect 23475 11396 23499 11398
rect 23555 11396 23579 11398
rect 23635 11396 23659 11398
rect 23715 11396 23721 11398
rect 23413 11376 23721 11396
rect 23296 11076 23348 11082
rect 23296 11018 23348 11024
rect 23308 10674 23336 11018
rect 23296 10668 23348 10674
rect 23216 10628 23296 10656
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 23124 8566 23152 9998
rect 23216 8974 23244 10628
rect 23296 10610 23348 10616
rect 23413 10364 23721 10384
rect 23413 10362 23419 10364
rect 23475 10362 23499 10364
rect 23555 10362 23579 10364
rect 23635 10362 23659 10364
rect 23715 10362 23721 10364
rect 23475 10310 23477 10362
rect 23657 10310 23659 10362
rect 23413 10308 23419 10310
rect 23475 10308 23499 10310
rect 23555 10308 23579 10310
rect 23635 10308 23659 10310
rect 23715 10308 23721 10310
rect 23413 10288 23721 10308
rect 23664 10192 23716 10198
rect 23664 10134 23716 10140
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 23308 9722 23336 9862
rect 23296 9716 23348 9722
rect 23296 9658 23348 9664
rect 23294 9616 23350 9625
rect 23676 9586 23704 10134
rect 23294 9551 23350 9560
rect 23664 9580 23716 9586
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 23112 8560 23164 8566
rect 23112 8502 23164 8508
rect 23204 8424 23256 8430
rect 23204 8366 23256 8372
rect 23216 8294 23244 8366
rect 23204 8288 23256 8294
rect 23204 8230 23256 8236
rect 23112 8084 23164 8090
rect 23032 8044 23112 8072
rect 23112 8026 23164 8032
rect 23216 7886 23244 8230
rect 23204 7880 23256 7886
rect 23204 7822 23256 7828
rect 23308 7818 23336 9551
rect 23664 9522 23716 9528
rect 23676 9450 23704 9522
rect 23768 9489 23796 11591
rect 23848 11008 23900 11014
rect 23848 10950 23900 10956
rect 23860 10674 23888 10950
rect 23848 10668 23900 10674
rect 23848 10610 23900 10616
rect 23940 10600 23992 10606
rect 23940 10542 23992 10548
rect 23754 9480 23810 9489
rect 23664 9444 23716 9450
rect 23754 9415 23810 9424
rect 23664 9386 23716 9392
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 23413 9276 23721 9296
rect 23413 9274 23419 9276
rect 23475 9274 23499 9276
rect 23555 9274 23579 9276
rect 23635 9274 23659 9276
rect 23715 9274 23721 9276
rect 23475 9222 23477 9274
rect 23657 9222 23659 9274
rect 23413 9220 23419 9222
rect 23475 9220 23499 9222
rect 23555 9220 23579 9222
rect 23635 9220 23659 9222
rect 23715 9220 23721 9222
rect 23413 9200 23721 9220
rect 23860 9042 23888 9318
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23952 8922 23980 10542
rect 23388 8900 23440 8906
rect 23388 8842 23440 8848
rect 23860 8894 23980 8922
rect 23400 8401 23428 8842
rect 23662 8664 23718 8673
rect 23662 8599 23664 8608
rect 23716 8599 23718 8608
rect 23664 8570 23716 8576
rect 23386 8392 23442 8401
rect 23386 8327 23442 8336
rect 23413 8188 23721 8208
rect 23413 8186 23419 8188
rect 23475 8186 23499 8188
rect 23555 8186 23579 8188
rect 23635 8186 23659 8188
rect 23715 8186 23721 8188
rect 23475 8134 23477 8186
rect 23657 8134 23659 8186
rect 23413 8132 23419 8134
rect 23475 8132 23499 8134
rect 23555 8132 23579 8134
rect 23635 8132 23659 8134
rect 23715 8132 23721 8134
rect 23413 8112 23721 8132
rect 23662 7984 23718 7993
rect 23662 7919 23718 7928
rect 23296 7812 23348 7818
rect 23296 7754 23348 7760
rect 23676 7546 23704 7919
rect 23756 7744 23808 7750
rect 23756 7686 23808 7692
rect 23664 7540 23716 7546
rect 23664 7482 23716 7488
rect 23768 7478 23796 7686
rect 23756 7472 23808 7478
rect 23756 7414 23808 7420
rect 23112 7404 23164 7410
rect 23112 7346 23164 7352
rect 23020 6656 23072 6662
rect 23020 6598 23072 6604
rect 23032 5914 23060 6598
rect 23020 5908 23072 5914
rect 23020 5850 23072 5856
rect 23124 5817 23152 7346
rect 23204 7200 23256 7206
rect 23204 7142 23256 7148
rect 23110 5808 23166 5817
rect 23110 5743 23166 5752
rect 23112 5704 23164 5710
rect 23112 5646 23164 5652
rect 22928 5296 22980 5302
rect 22928 5238 22980 5244
rect 22744 5160 22796 5166
rect 23020 5160 23072 5166
rect 22796 5120 22876 5148
rect 22744 5102 22796 5108
rect 22744 5024 22796 5030
rect 22744 4966 22796 4972
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 20720 2372 20772 2378
rect 20720 2314 20772 2320
rect 20996 2372 21048 2378
rect 20996 2314 21048 2320
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 21284 1970 21312 2246
rect 21272 1964 21324 1970
rect 21272 1906 21324 1912
rect 21088 1488 21140 1494
rect 21088 1430 21140 1436
rect 21100 800 21128 1430
rect 21640 1420 21692 1426
rect 21640 1362 21692 1368
rect 21652 800 21680 1362
rect 22204 800 22232 2246
rect 22756 800 22784 4966
rect 22848 4758 22876 5120
rect 23020 5102 23072 5108
rect 22836 4752 22888 4758
rect 22836 4694 22888 4700
rect 22848 3754 22876 4694
rect 23032 4622 23060 5102
rect 23020 4616 23072 4622
rect 23020 4558 23072 4564
rect 22928 4480 22980 4486
rect 22928 4422 22980 4428
rect 22940 4214 22968 4422
rect 22928 4208 22980 4214
rect 22928 4150 22980 4156
rect 23020 4140 23072 4146
rect 23020 4082 23072 4088
rect 23032 3754 23060 4082
rect 22848 3726 23060 3754
rect 23124 3738 23152 5646
rect 23032 3516 23060 3726
rect 23112 3732 23164 3738
rect 23112 3674 23164 3680
rect 23112 3528 23164 3534
rect 23032 3488 23112 3516
rect 23112 3470 23164 3476
rect 23112 3052 23164 3058
rect 23112 2994 23164 3000
rect 23020 2576 23072 2582
rect 23020 2518 23072 2524
rect 23032 1426 23060 2518
rect 23124 1442 23152 2994
rect 23216 2446 23244 7142
rect 23413 7100 23721 7120
rect 23413 7098 23419 7100
rect 23475 7098 23499 7100
rect 23555 7098 23579 7100
rect 23635 7098 23659 7100
rect 23715 7098 23721 7100
rect 23475 7046 23477 7098
rect 23657 7046 23659 7098
rect 23413 7044 23419 7046
rect 23475 7044 23499 7046
rect 23555 7044 23579 7046
rect 23635 7044 23659 7046
rect 23715 7044 23721 7046
rect 23413 7024 23721 7044
rect 23294 6488 23350 6497
rect 23294 6423 23350 6432
rect 23308 4758 23336 6423
rect 23413 6012 23721 6032
rect 23413 6010 23419 6012
rect 23475 6010 23499 6012
rect 23555 6010 23579 6012
rect 23635 6010 23659 6012
rect 23715 6010 23721 6012
rect 23475 5958 23477 6010
rect 23657 5958 23659 6010
rect 23413 5956 23419 5958
rect 23475 5956 23499 5958
rect 23555 5956 23579 5958
rect 23635 5956 23659 5958
rect 23715 5956 23721 5958
rect 23413 5936 23721 5956
rect 23768 5710 23796 7414
rect 23860 5846 23888 8894
rect 23940 8832 23992 8838
rect 23940 8774 23992 8780
rect 23848 5840 23900 5846
rect 23848 5782 23900 5788
rect 23756 5704 23808 5710
rect 23756 5646 23808 5652
rect 23848 5568 23900 5574
rect 23478 5536 23534 5545
rect 23848 5510 23900 5516
rect 23478 5471 23534 5480
rect 23492 5370 23520 5471
rect 23480 5364 23532 5370
rect 23480 5306 23532 5312
rect 23664 5296 23716 5302
rect 23716 5256 23796 5284
rect 23664 5238 23716 5244
rect 23413 4924 23721 4944
rect 23413 4922 23419 4924
rect 23475 4922 23499 4924
rect 23555 4922 23579 4924
rect 23635 4922 23659 4924
rect 23715 4922 23721 4924
rect 23475 4870 23477 4922
rect 23657 4870 23659 4922
rect 23413 4868 23419 4870
rect 23475 4868 23499 4870
rect 23555 4868 23579 4870
rect 23635 4868 23659 4870
rect 23715 4868 23721 4870
rect 23413 4848 23721 4868
rect 23296 4752 23348 4758
rect 23296 4694 23348 4700
rect 23386 4720 23442 4729
rect 23386 4655 23442 4664
rect 23400 4622 23428 4655
rect 23388 4616 23440 4622
rect 23308 4576 23388 4604
rect 23308 3534 23336 4576
rect 23388 4558 23440 4564
rect 23480 4480 23532 4486
rect 23480 4422 23532 4428
rect 23492 4282 23520 4422
rect 23768 4282 23796 5256
rect 23480 4276 23532 4282
rect 23480 4218 23532 4224
rect 23756 4276 23808 4282
rect 23756 4218 23808 4224
rect 23756 4072 23808 4078
rect 23756 4014 23808 4020
rect 23413 3836 23721 3856
rect 23413 3834 23419 3836
rect 23475 3834 23499 3836
rect 23555 3834 23579 3836
rect 23635 3834 23659 3836
rect 23715 3834 23721 3836
rect 23475 3782 23477 3834
rect 23657 3782 23659 3834
rect 23413 3780 23419 3782
rect 23475 3780 23499 3782
rect 23555 3780 23579 3782
rect 23635 3780 23659 3782
rect 23715 3780 23721 3782
rect 23413 3760 23721 3780
rect 23296 3528 23348 3534
rect 23296 3470 23348 3476
rect 23296 3392 23348 3398
rect 23296 3334 23348 3340
rect 23308 2854 23336 3334
rect 23768 3058 23796 4014
rect 23756 3052 23808 3058
rect 23756 2994 23808 3000
rect 23296 2848 23348 2854
rect 23296 2790 23348 2796
rect 23308 2514 23336 2790
rect 23413 2748 23721 2768
rect 23413 2746 23419 2748
rect 23475 2746 23499 2748
rect 23555 2746 23579 2748
rect 23635 2746 23659 2748
rect 23715 2746 23721 2748
rect 23475 2694 23477 2746
rect 23657 2694 23659 2746
rect 23413 2692 23419 2694
rect 23475 2692 23499 2694
rect 23555 2692 23579 2694
rect 23635 2692 23659 2694
rect 23715 2692 23721 2694
rect 23413 2672 23721 2692
rect 23296 2508 23348 2514
rect 23296 2450 23348 2456
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 23388 2304 23440 2310
rect 23388 2246 23440 2252
rect 23400 1494 23428 2246
rect 23388 1488 23440 1494
rect 23020 1420 23072 1426
rect 23124 1414 23336 1442
rect 23388 1430 23440 1436
rect 23020 1362 23072 1368
rect 23308 800 23336 1414
rect 23860 800 23888 5510
rect 23952 2514 23980 8774
rect 24044 6798 24072 12038
rect 24228 11762 24256 13806
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 24320 11558 24348 14282
rect 24412 12238 24440 14962
rect 24400 12232 24452 12238
rect 24400 12174 24452 12180
rect 24216 11552 24268 11558
rect 24216 11494 24268 11500
rect 24308 11552 24360 11558
rect 24308 11494 24360 11500
rect 24228 11286 24256 11494
rect 24216 11280 24268 11286
rect 24216 11222 24268 11228
rect 24124 11008 24176 11014
rect 24124 10950 24176 10956
rect 24136 8809 24164 10950
rect 24228 10674 24256 11222
rect 24308 11212 24360 11218
rect 24308 11154 24360 11160
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 24228 10062 24256 10610
rect 24216 10056 24268 10062
rect 24216 9998 24268 10004
rect 24228 8974 24256 9998
rect 24216 8968 24268 8974
rect 24216 8910 24268 8916
rect 24122 8800 24178 8809
rect 24122 8735 24178 8744
rect 24228 8498 24256 8910
rect 24124 8492 24176 8498
rect 24124 8434 24176 8440
rect 24216 8492 24268 8498
rect 24216 8434 24268 8440
rect 24032 6792 24084 6798
rect 24032 6734 24084 6740
rect 24032 6656 24084 6662
rect 24032 6598 24084 6604
rect 24044 2854 24072 6598
rect 24032 2848 24084 2854
rect 24032 2790 24084 2796
rect 23940 2508 23992 2514
rect 23940 2450 23992 2456
rect 24136 1970 24164 8434
rect 24320 7886 24348 11154
rect 24412 11150 24440 12174
rect 24400 11144 24452 11150
rect 24400 11086 24452 11092
rect 24504 11014 24532 19306
rect 24492 11008 24544 11014
rect 24492 10950 24544 10956
rect 24490 10160 24546 10169
rect 24490 10095 24546 10104
rect 24400 8288 24452 8294
rect 24400 8230 24452 8236
rect 24308 7880 24360 7886
rect 24308 7822 24360 7828
rect 24216 7812 24268 7818
rect 24216 7754 24268 7760
rect 24228 7546 24256 7754
rect 24216 7540 24268 7546
rect 24216 7482 24268 7488
rect 24308 7472 24360 7478
rect 24308 7414 24360 7420
rect 24320 7342 24348 7414
rect 24308 7336 24360 7342
rect 24308 7278 24360 7284
rect 24216 7268 24268 7274
rect 24216 7210 24268 7216
rect 24228 6798 24256 7210
rect 24306 7168 24362 7177
rect 24306 7103 24362 7112
rect 24216 6792 24268 6798
rect 24216 6734 24268 6740
rect 24320 6458 24348 7103
rect 24412 7002 24440 8230
rect 24400 6996 24452 7002
rect 24400 6938 24452 6944
rect 24398 6896 24454 6905
rect 24398 6831 24454 6840
rect 24412 6730 24440 6831
rect 24400 6724 24452 6730
rect 24400 6666 24452 6672
rect 24398 6624 24454 6633
rect 24398 6559 24454 6568
rect 24308 6452 24360 6458
rect 24308 6394 24360 6400
rect 24216 6384 24268 6390
rect 24216 6326 24268 6332
rect 24228 5574 24256 6326
rect 24308 6112 24360 6118
rect 24308 6054 24360 6060
rect 24320 5642 24348 6054
rect 24308 5636 24360 5642
rect 24308 5578 24360 5584
rect 24216 5568 24268 5574
rect 24216 5510 24268 5516
rect 24228 5302 24256 5510
rect 24412 5386 24440 6559
rect 24504 5930 24532 10095
rect 24596 7886 24624 21558
rect 24768 21548 24820 21554
rect 24768 21490 24820 21496
rect 24676 21412 24728 21418
rect 24676 21354 24728 21360
rect 24688 19553 24716 21354
rect 24780 19922 24808 21490
rect 24964 21010 24992 24550
rect 25056 24070 25084 24686
rect 25044 24064 25096 24070
rect 25044 24006 25096 24012
rect 25044 22568 25096 22574
rect 25044 22510 25096 22516
rect 25056 21962 25084 22510
rect 25044 21956 25096 21962
rect 25044 21898 25096 21904
rect 25056 21554 25084 21898
rect 25044 21548 25096 21554
rect 25044 21490 25096 21496
rect 24952 21004 25004 21010
rect 24952 20946 25004 20952
rect 25056 20890 25084 21490
rect 24964 20862 25084 20890
rect 24860 20528 24912 20534
rect 24860 20470 24912 20476
rect 24768 19916 24820 19922
rect 24768 19858 24820 19864
rect 24768 19712 24820 19718
rect 24768 19654 24820 19660
rect 24674 19544 24730 19553
rect 24674 19479 24730 19488
rect 24780 19446 24808 19654
rect 24768 19440 24820 19446
rect 24768 19382 24820 19388
rect 24872 19258 24900 20470
rect 24964 20466 24992 20862
rect 25044 20800 25096 20806
rect 25044 20742 25096 20748
rect 25056 20534 25084 20742
rect 25044 20528 25096 20534
rect 25044 20470 25096 20476
rect 24952 20460 25004 20466
rect 24952 20402 25004 20408
rect 24952 20324 25004 20330
rect 24952 20266 25004 20272
rect 24780 19230 24900 19258
rect 24676 18420 24728 18426
rect 24676 18362 24728 18368
rect 24688 17202 24716 18362
rect 24676 17196 24728 17202
rect 24676 17138 24728 17144
rect 24676 16516 24728 16522
rect 24676 16458 24728 16464
rect 24688 16250 24716 16458
rect 24676 16244 24728 16250
rect 24676 16186 24728 16192
rect 24676 16108 24728 16114
rect 24676 16050 24728 16056
rect 24688 15570 24716 16050
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24688 15026 24716 15506
rect 24676 15020 24728 15026
rect 24676 14962 24728 14968
rect 24688 13938 24716 14962
rect 24676 13932 24728 13938
rect 24676 13874 24728 13880
rect 24688 13326 24716 13874
rect 24676 13320 24728 13326
rect 24676 13262 24728 13268
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24688 11694 24716 12922
rect 24780 12782 24808 19230
rect 24964 19174 24992 20266
rect 25044 19712 25096 19718
rect 25044 19654 25096 19660
rect 25056 19174 25084 19654
rect 24952 19168 25004 19174
rect 24952 19110 25004 19116
rect 25044 19168 25096 19174
rect 25044 19110 25096 19116
rect 24860 18760 24912 18766
rect 24860 18702 24912 18708
rect 24872 18222 24900 18702
rect 24964 18630 24992 19110
rect 25148 18698 25176 27270
rect 25240 19922 25268 27542
rect 25780 27328 25832 27334
rect 25780 27270 25832 27276
rect 25688 26784 25740 26790
rect 25688 26726 25740 26732
rect 25412 26376 25464 26382
rect 25412 26318 25464 26324
rect 25424 25362 25452 26318
rect 25504 26308 25556 26314
rect 25504 26250 25556 26256
rect 25412 25356 25464 25362
rect 25412 25298 25464 25304
rect 25320 24608 25372 24614
rect 25320 24550 25372 24556
rect 25332 24206 25360 24550
rect 25424 24274 25452 25298
rect 25516 24410 25544 26250
rect 25596 24608 25648 24614
rect 25596 24550 25648 24556
rect 25504 24404 25556 24410
rect 25504 24346 25556 24352
rect 25412 24268 25464 24274
rect 25412 24210 25464 24216
rect 25320 24200 25372 24206
rect 25320 24142 25372 24148
rect 25504 24064 25556 24070
rect 25504 24006 25556 24012
rect 25516 23798 25544 24006
rect 25320 23792 25372 23798
rect 25320 23734 25372 23740
rect 25504 23792 25556 23798
rect 25608 23769 25636 24550
rect 25700 23866 25728 26726
rect 25688 23860 25740 23866
rect 25688 23802 25740 23808
rect 25504 23734 25556 23740
rect 25594 23760 25650 23769
rect 25332 23526 25360 23734
rect 25516 23644 25544 23734
rect 25594 23695 25650 23704
rect 25424 23616 25544 23644
rect 25596 23656 25648 23662
rect 25320 23520 25372 23526
rect 25320 23462 25372 23468
rect 25332 22710 25360 23462
rect 25320 22704 25372 22710
rect 25320 22646 25372 22652
rect 25332 20874 25360 22646
rect 25320 20868 25372 20874
rect 25320 20810 25372 20816
rect 25228 19916 25280 19922
rect 25228 19858 25280 19864
rect 25228 19712 25280 19718
rect 25228 19654 25280 19660
rect 25136 18692 25188 18698
rect 25136 18634 25188 18640
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24860 18216 24912 18222
rect 24860 18158 24912 18164
rect 24860 17536 24912 17542
rect 24860 17478 24912 17484
rect 24872 17202 24900 17478
rect 24860 17196 24912 17202
rect 24860 17138 24912 17144
rect 24964 17082 24992 18566
rect 25044 18216 25096 18222
rect 25044 18158 25096 18164
rect 25056 17678 25084 18158
rect 25044 17672 25096 17678
rect 25044 17614 25096 17620
rect 24872 17054 24992 17082
rect 24872 14006 24900 17054
rect 25056 16658 25084 17614
rect 25136 17196 25188 17202
rect 25136 17138 25188 17144
rect 25148 16794 25176 17138
rect 25136 16788 25188 16794
rect 25136 16730 25188 16736
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 25240 16538 25268 19654
rect 25320 19304 25372 19310
rect 25320 19246 25372 19252
rect 25332 19174 25360 19246
rect 25320 19168 25372 19174
rect 25320 19110 25372 19116
rect 25332 18086 25360 19110
rect 25320 18080 25372 18086
rect 25320 18022 25372 18028
rect 24964 16510 25268 16538
rect 24860 14000 24912 14006
rect 24860 13942 24912 13948
rect 24964 13716 24992 16510
rect 25228 16448 25280 16454
rect 25228 16390 25280 16396
rect 25136 16176 25188 16182
rect 25136 16118 25188 16124
rect 25148 15065 25176 16118
rect 25240 15706 25268 16390
rect 25228 15700 25280 15706
rect 25228 15642 25280 15648
rect 25228 15360 25280 15366
rect 25228 15302 25280 15308
rect 25134 15056 25190 15065
rect 25134 14991 25190 15000
rect 25136 14952 25188 14958
rect 25136 14894 25188 14900
rect 25148 14074 25176 14894
rect 25136 14068 25188 14074
rect 25136 14010 25188 14016
rect 25148 13938 25176 14010
rect 25136 13932 25188 13938
rect 24872 13688 24992 13716
rect 25056 13892 25136 13920
rect 24872 13138 24900 13688
rect 24952 13320 25004 13326
rect 25056 13308 25084 13892
rect 25136 13874 25188 13880
rect 25240 13841 25268 15302
rect 25332 14385 25360 18022
rect 25424 16182 25452 23616
rect 25596 23598 25648 23604
rect 25608 23254 25636 23598
rect 25688 23588 25740 23594
rect 25688 23530 25740 23536
rect 25596 23248 25648 23254
rect 25596 23190 25648 23196
rect 25504 22976 25556 22982
rect 25504 22918 25556 22924
rect 25516 22778 25544 22918
rect 25504 22772 25556 22778
rect 25504 22714 25556 22720
rect 25516 21962 25544 22714
rect 25700 22234 25728 23530
rect 25688 22228 25740 22234
rect 25688 22170 25740 22176
rect 25504 21956 25556 21962
rect 25504 21898 25556 21904
rect 25412 16176 25464 16182
rect 25412 16118 25464 16124
rect 25412 15700 25464 15706
rect 25412 15642 25464 15648
rect 25318 14376 25374 14385
rect 25318 14311 25374 14320
rect 25424 13954 25452 15642
rect 25332 13926 25452 13954
rect 25516 13938 25544 21898
rect 25596 21888 25648 21894
rect 25596 21830 25648 21836
rect 25688 21888 25740 21894
rect 25688 21830 25740 21836
rect 25608 21622 25636 21830
rect 25700 21690 25728 21830
rect 25688 21684 25740 21690
rect 25688 21626 25740 21632
rect 25596 21616 25648 21622
rect 25596 21558 25648 21564
rect 25688 21344 25740 21350
rect 25688 21286 25740 21292
rect 25596 20800 25648 20806
rect 25596 20742 25648 20748
rect 25608 20466 25636 20742
rect 25596 20460 25648 20466
rect 25596 20402 25648 20408
rect 25608 19718 25636 20402
rect 25596 19712 25648 19718
rect 25596 19654 25648 19660
rect 25504 13932 25556 13938
rect 25226 13832 25282 13841
rect 25136 13796 25188 13802
rect 25226 13767 25282 13776
rect 25136 13738 25188 13744
rect 25004 13280 25084 13308
rect 24952 13262 25004 13268
rect 24872 13110 24992 13138
rect 24860 12844 24912 12850
rect 24860 12786 24912 12792
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 24768 11824 24820 11830
rect 24768 11766 24820 11772
rect 24676 11688 24728 11694
rect 24676 11630 24728 11636
rect 24780 10674 24808 11766
rect 24872 10742 24900 12786
rect 24860 10736 24912 10742
rect 24860 10678 24912 10684
rect 24768 10668 24820 10674
rect 24768 10610 24820 10616
rect 24780 10198 24808 10610
rect 24768 10192 24820 10198
rect 24768 10134 24820 10140
rect 24676 10056 24728 10062
rect 24676 9998 24728 10004
rect 24584 7880 24636 7886
rect 24584 7822 24636 7828
rect 24584 7744 24636 7750
rect 24584 7686 24636 7692
rect 24596 7478 24624 7686
rect 24584 7472 24636 7478
rect 24584 7414 24636 7420
rect 24596 7041 24624 7414
rect 24688 7177 24716 9998
rect 24780 9042 24808 10134
rect 24860 9444 24912 9450
rect 24860 9386 24912 9392
rect 24768 9036 24820 9042
rect 24768 8978 24820 8984
rect 24872 8906 24900 9386
rect 24860 8900 24912 8906
rect 24860 8842 24912 8848
rect 24964 8786 24992 13110
rect 25044 12232 25096 12238
rect 25044 12174 25096 12180
rect 25148 12186 25176 13738
rect 25056 11082 25084 12174
rect 25148 12158 25268 12186
rect 25136 12096 25188 12102
rect 25136 12038 25188 12044
rect 25148 11762 25176 12038
rect 25136 11756 25188 11762
rect 25136 11698 25188 11704
rect 25044 11076 25096 11082
rect 25044 11018 25096 11024
rect 25240 9654 25268 12158
rect 25228 9648 25280 9654
rect 25228 9590 25280 9596
rect 25332 9450 25360 13926
rect 25504 13874 25556 13880
rect 25412 13864 25464 13870
rect 25412 13806 25464 13812
rect 25424 13394 25452 13806
rect 25412 13388 25464 13394
rect 25412 13330 25464 13336
rect 25608 13326 25636 19654
rect 25700 16130 25728 21286
rect 25792 20942 25820 27270
rect 25884 22574 25912 27882
rect 26608 27872 26660 27878
rect 26608 27814 26660 27820
rect 26056 27464 26108 27470
rect 26056 27406 26108 27412
rect 25964 26988 26016 26994
rect 25964 26930 26016 26936
rect 25976 24410 26004 26930
rect 25964 24404 26016 24410
rect 25964 24346 26016 24352
rect 25964 24268 26016 24274
rect 25964 24210 26016 24216
rect 25976 23186 26004 24210
rect 25964 23180 26016 23186
rect 25964 23122 26016 23128
rect 25872 22568 25924 22574
rect 25872 22510 25924 22516
rect 25872 22432 25924 22438
rect 25872 22374 25924 22380
rect 25884 22030 25912 22374
rect 25872 22024 25924 22030
rect 25872 21966 25924 21972
rect 25870 21720 25926 21729
rect 25976 21690 26004 23122
rect 26068 22166 26096 27406
rect 26332 27328 26384 27334
rect 26332 27270 26384 27276
rect 26240 26784 26292 26790
rect 26240 26726 26292 26732
rect 26148 25832 26200 25838
rect 26148 25774 26200 25780
rect 26160 24138 26188 25774
rect 26252 25294 26280 26726
rect 26240 25288 26292 25294
rect 26240 25230 26292 25236
rect 26240 24812 26292 24818
rect 26240 24754 26292 24760
rect 26148 24132 26200 24138
rect 26148 24074 26200 24080
rect 26160 22574 26188 24074
rect 26148 22568 26200 22574
rect 26148 22510 26200 22516
rect 26148 22228 26200 22234
rect 26148 22170 26200 22176
rect 26056 22160 26108 22166
rect 26056 22102 26108 22108
rect 26056 22024 26108 22030
rect 26056 21966 26108 21972
rect 25870 21655 25926 21664
rect 25964 21684 26016 21690
rect 25780 20936 25832 20942
rect 25780 20878 25832 20884
rect 25780 20460 25832 20466
rect 25780 20402 25832 20408
rect 25792 19553 25820 20402
rect 25884 19786 25912 21655
rect 25964 21626 26016 21632
rect 25976 21010 26004 21626
rect 26068 21554 26096 21966
rect 26160 21729 26188 22170
rect 26252 21962 26280 24754
rect 26344 23050 26372 27270
rect 26424 26988 26476 26994
rect 26424 26930 26476 26936
rect 26436 26042 26464 26930
rect 26516 26512 26568 26518
rect 26516 26454 26568 26460
rect 26424 26036 26476 26042
rect 26424 25978 26476 25984
rect 26424 25900 26476 25906
rect 26424 25842 26476 25848
rect 26436 24993 26464 25842
rect 26422 24984 26478 24993
rect 26422 24919 26478 24928
rect 26528 24206 26556 26454
rect 26516 24200 26568 24206
rect 26516 24142 26568 24148
rect 26332 23044 26384 23050
rect 26332 22986 26384 22992
rect 26620 22094 26648 27814
rect 26700 26376 26752 26382
rect 26700 26318 26752 26324
rect 26528 22066 26648 22094
rect 26240 21956 26292 21962
rect 26240 21898 26292 21904
rect 26146 21720 26202 21729
rect 26146 21655 26202 21664
rect 26148 21616 26200 21622
rect 26148 21558 26200 21564
rect 26056 21548 26108 21554
rect 26056 21490 26108 21496
rect 25964 21004 26016 21010
rect 25964 20946 26016 20952
rect 25976 19922 26004 20946
rect 26160 20806 26188 21558
rect 26240 21548 26292 21554
rect 26240 21490 26292 21496
rect 26148 20800 26200 20806
rect 26148 20742 26200 20748
rect 25964 19916 26016 19922
rect 25964 19858 26016 19864
rect 25872 19780 25924 19786
rect 25872 19722 25924 19728
rect 25962 19680 26018 19689
rect 25962 19615 26018 19624
rect 25778 19544 25834 19553
rect 25778 19479 25834 19488
rect 25792 19378 25820 19479
rect 25780 19372 25832 19378
rect 25780 19314 25832 19320
rect 25780 17672 25832 17678
rect 25780 17614 25832 17620
rect 25792 16250 25820 17614
rect 25976 17202 26004 19615
rect 26056 19372 26108 19378
rect 26056 19314 26108 19320
rect 25964 17196 26016 17202
rect 25884 17156 25964 17184
rect 25884 16454 25912 17156
rect 25964 17138 26016 17144
rect 25964 17060 26016 17066
rect 25964 17002 26016 17008
rect 25976 16658 26004 17002
rect 25964 16652 26016 16658
rect 25964 16594 26016 16600
rect 25872 16448 25924 16454
rect 25872 16390 25924 16396
rect 25780 16244 25832 16250
rect 25780 16186 25832 16192
rect 25700 16102 25820 16130
rect 25688 15972 25740 15978
rect 25688 15914 25740 15920
rect 25700 15026 25728 15914
rect 25688 15020 25740 15026
rect 25688 14962 25740 14968
rect 25688 14000 25740 14006
rect 25688 13942 25740 13948
rect 25596 13320 25648 13326
rect 25596 13262 25648 13268
rect 25412 13184 25464 13190
rect 25412 13126 25464 13132
rect 25424 12238 25452 13126
rect 25504 12300 25556 12306
rect 25504 12242 25556 12248
rect 25412 12232 25464 12238
rect 25412 12174 25464 12180
rect 25516 11898 25544 12242
rect 25504 11892 25556 11898
rect 25504 11834 25556 11840
rect 25596 11756 25648 11762
rect 25516 11716 25596 11744
rect 25516 11218 25544 11716
rect 25596 11698 25648 11704
rect 25504 11212 25556 11218
rect 25504 11154 25556 11160
rect 25596 11008 25648 11014
rect 25596 10950 25648 10956
rect 25504 10668 25556 10674
rect 25504 10610 25556 10616
rect 25516 9674 25544 10610
rect 25424 9646 25544 9674
rect 25320 9444 25372 9450
rect 25320 9386 25372 9392
rect 24964 8758 25268 8786
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25044 7880 25096 7886
rect 25044 7822 25096 7828
rect 24950 7440 25006 7449
rect 24950 7375 24952 7384
rect 25004 7375 25006 7384
rect 24952 7346 25004 7352
rect 25056 7290 25084 7822
rect 24964 7262 25084 7290
rect 24860 7200 24912 7206
rect 24674 7168 24730 7177
rect 24860 7142 24912 7148
rect 24674 7103 24730 7112
rect 24582 7032 24638 7041
rect 24872 7002 24900 7142
rect 24582 6967 24638 6976
rect 24676 6996 24728 7002
rect 24676 6938 24728 6944
rect 24860 6996 24912 7002
rect 24860 6938 24912 6944
rect 24688 6186 24716 6938
rect 24766 6760 24822 6769
rect 24964 6746 24992 7262
rect 25044 7200 25096 7206
rect 25044 7142 25096 7148
rect 25056 6769 25084 7142
rect 24766 6695 24822 6704
rect 24872 6718 24992 6746
rect 25042 6760 25098 6769
rect 24780 6662 24808 6695
rect 24768 6656 24820 6662
rect 24768 6598 24820 6604
rect 24780 6458 24808 6598
rect 24768 6452 24820 6458
rect 24768 6394 24820 6400
rect 24768 6316 24820 6322
rect 24768 6258 24820 6264
rect 24676 6180 24728 6186
rect 24676 6122 24728 6128
rect 24504 5902 24624 5930
rect 24688 5914 24716 6122
rect 24492 5840 24544 5846
rect 24492 5782 24544 5788
rect 24320 5358 24440 5386
rect 24216 5296 24268 5302
rect 24216 5238 24268 5244
rect 24214 5128 24270 5137
rect 24214 5063 24270 5072
rect 24228 5030 24256 5063
rect 24216 5024 24268 5030
rect 24216 4966 24268 4972
rect 24320 4826 24348 5358
rect 24400 5296 24452 5302
rect 24400 5238 24452 5244
rect 24308 4820 24360 4826
rect 24308 4762 24360 4768
rect 24308 4616 24360 4622
rect 24308 4558 24360 4564
rect 24320 2446 24348 4558
rect 24412 4486 24440 5238
rect 24400 4480 24452 4486
rect 24400 4422 24452 4428
rect 24412 4282 24440 4422
rect 24400 4276 24452 4282
rect 24400 4218 24452 4224
rect 24400 3392 24452 3398
rect 24400 3334 24452 3340
rect 24412 3126 24440 3334
rect 24400 3120 24452 3126
rect 24400 3062 24452 3068
rect 24504 2774 24532 5782
rect 24596 5710 24624 5902
rect 24676 5908 24728 5914
rect 24676 5850 24728 5856
rect 24584 5704 24636 5710
rect 24584 5646 24636 5652
rect 24584 5568 24636 5574
rect 24584 5510 24636 5516
rect 24596 5302 24624 5510
rect 24584 5296 24636 5302
rect 24584 5238 24636 5244
rect 24688 5137 24716 5850
rect 24780 5778 24808 6258
rect 24768 5772 24820 5778
rect 24768 5714 24820 5720
rect 24872 5302 24900 6718
rect 25042 6695 25098 6704
rect 24952 6656 25004 6662
rect 24952 6598 25004 6604
rect 24860 5296 24912 5302
rect 24860 5238 24912 5244
rect 24674 5128 24730 5137
rect 24674 5063 24730 5072
rect 24575 5024 24627 5030
rect 24688 5012 24716 5063
rect 24627 4984 24716 5012
rect 24575 4966 24627 4972
rect 24860 4548 24912 4554
rect 24860 4490 24912 4496
rect 24584 4140 24636 4146
rect 24584 4082 24636 4088
rect 24768 4140 24820 4146
rect 24768 4082 24820 4088
rect 24596 3534 24624 4082
rect 24780 3534 24808 4082
rect 24872 4010 24900 4490
rect 24860 4004 24912 4010
rect 24860 3946 24912 3952
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24780 3194 24808 3334
rect 24768 3188 24820 3194
rect 24768 3130 24820 3136
rect 24412 2746 24532 2774
rect 24308 2440 24360 2446
rect 24308 2382 24360 2388
rect 24124 1964 24176 1970
rect 24124 1906 24176 1912
rect 24412 800 24440 2746
rect 24964 800 24992 6598
rect 25042 6488 25098 6497
rect 25042 6423 25098 6432
rect 25056 6390 25084 6423
rect 25044 6384 25096 6390
rect 25044 6326 25096 6332
rect 25148 2446 25176 8570
rect 25240 6458 25268 8758
rect 25318 8664 25374 8673
rect 25318 8599 25320 8608
rect 25372 8599 25374 8608
rect 25320 8570 25372 8576
rect 25318 8392 25374 8401
rect 25318 8327 25374 8336
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 25332 3398 25360 8327
rect 25424 5545 25452 9646
rect 25504 9376 25556 9382
rect 25504 9318 25556 9324
rect 25516 8974 25544 9318
rect 25504 8968 25556 8974
rect 25504 8910 25556 8916
rect 25504 7404 25556 7410
rect 25504 7346 25556 7352
rect 25516 7313 25544 7346
rect 25502 7304 25558 7313
rect 25502 7239 25558 7248
rect 25504 6860 25556 6866
rect 25504 6802 25556 6808
rect 25516 5778 25544 6802
rect 25504 5772 25556 5778
rect 25504 5714 25556 5720
rect 25410 5536 25466 5545
rect 25410 5471 25466 5480
rect 25412 3936 25464 3942
rect 25412 3878 25464 3884
rect 25320 3392 25372 3398
rect 25320 3334 25372 3340
rect 25136 2440 25188 2446
rect 25136 2382 25188 2388
rect 25424 800 25452 3878
rect 25608 3670 25636 10950
rect 25700 5710 25728 13942
rect 25792 12850 25820 16102
rect 25872 16108 25924 16114
rect 25872 16050 25924 16056
rect 25884 15366 25912 16050
rect 25976 15570 26004 16594
rect 25964 15564 26016 15570
rect 25964 15506 26016 15512
rect 25872 15360 25924 15366
rect 25872 15302 25924 15308
rect 25872 14952 25924 14958
rect 25872 14894 25924 14900
rect 25884 14346 25912 14894
rect 25976 14482 26004 15506
rect 25964 14476 26016 14482
rect 25964 14418 26016 14424
rect 25872 14340 25924 14346
rect 25872 14282 25924 14288
rect 25884 13870 25912 14282
rect 26068 13954 26096 19314
rect 26160 15026 26188 20742
rect 26252 19281 26280 21490
rect 26332 20392 26384 20398
rect 26332 20334 26384 20340
rect 26344 20058 26372 20334
rect 26332 20052 26384 20058
rect 26332 19994 26384 20000
rect 26344 19310 26372 19994
rect 26424 19508 26476 19514
rect 26424 19450 26476 19456
rect 26332 19304 26384 19310
rect 26238 19272 26294 19281
rect 26332 19246 26384 19252
rect 26238 19207 26294 19216
rect 26252 17338 26280 19207
rect 26332 17536 26384 17542
rect 26332 17478 26384 17484
rect 26240 17332 26292 17338
rect 26240 17274 26292 17280
rect 26240 17128 26292 17134
rect 26240 17070 26292 17076
rect 26252 16590 26280 17070
rect 26240 16584 26292 16590
rect 26240 16526 26292 16532
rect 26240 15904 26292 15910
rect 26240 15846 26292 15852
rect 26148 15020 26200 15026
rect 26148 14962 26200 14968
rect 25976 13926 26096 13954
rect 25872 13864 25924 13870
rect 25872 13806 25924 13812
rect 25976 13410 26004 13926
rect 26056 13864 26108 13870
rect 26056 13806 26108 13812
rect 25884 13382 26004 13410
rect 25780 12844 25832 12850
rect 25780 12786 25832 12792
rect 25884 12345 25912 13382
rect 25964 13320 26016 13326
rect 25964 13262 26016 13268
rect 25976 12918 26004 13262
rect 25964 12912 26016 12918
rect 25964 12854 26016 12860
rect 25870 12336 25926 12345
rect 25976 12306 26004 12854
rect 25870 12271 25926 12280
rect 25964 12300 26016 12306
rect 25964 12242 26016 12248
rect 25780 9920 25832 9926
rect 25780 9862 25832 9868
rect 25792 9586 25820 9862
rect 25870 9752 25926 9761
rect 26068 9738 26096 13806
rect 26148 13728 26200 13734
rect 26148 13670 26200 13676
rect 26160 12850 26188 13670
rect 26252 13530 26280 15846
rect 26344 15434 26372 17478
rect 26332 15428 26384 15434
rect 26332 15370 26384 15376
rect 26240 13524 26292 13530
rect 26240 13466 26292 13472
rect 26436 13433 26464 19450
rect 26528 18358 26556 22066
rect 26608 21480 26660 21486
rect 26608 21422 26660 21428
rect 26516 18352 26568 18358
rect 26516 18294 26568 18300
rect 26516 17672 26568 17678
rect 26516 17614 26568 17620
rect 26528 16998 26556 17614
rect 26516 16992 26568 16998
rect 26516 16934 26568 16940
rect 26620 16946 26648 21422
rect 26712 17338 26740 26318
rect 26792 25696 26844 25702
rect 26792 25638 26844 25644
rect 26804 25129 26832 25638
rect 26790 25120 26846 25129
rect 26790 25055 26846 25064
rect 26792 22568 26844 22574
rect 26792 22510 26844 22516
rect 26804 22098 26832 22510
rect 26792 22092 26844 22098
rect 26792 22034 26844 22040
rect 26792 21956 26844 21962
rect 26792 21898 26844 21904
rect 26804 18970 26832 21898
rect 26896 19514 26924 28018
rect 26976 27464 27028 27470
rect 26976 27406 27028 27412
rect 26988 22778 27016 27406
rect 27080 25242 27108 28358
rect 27160 28076 27212 28082
rect 27160 28018 27212 28024
rect 27172 27606 27200 28018
rect 27160 27600 27212 27606
rect 27160 27542 27212 27548
rect 27160 27464 27212 27470
rect 27160 27406 27212 27412
rect 27172 27130 27200 27406
rect 27252 27328 27304 27334
rect 27250 27296 27252 27305
rect 27304 27296 27306 27305
rect 27250 27231 27306 27240
rect 27160 27124 27212 27130
rect 27160 27066 27212 27072
rect 27160 25900 27212 25906
rect 27160 25842 27212 25848
rect 27172 25401 27200 25842
rect 27158 25392 27214 25401
rect 27158 25327 27214 25336
rect 27080 25214 27292 25242
rect 27068 24608 27120 24614
rect 27068 24550 27120 24556
rect 26976 22772 27028 22778
rect 26976 22714 27028 22720
rect 26976 21548 27028 21554
rect 26976 21490 27028 21496
rect 26884 19508 26936 19514
rect 26884 19450 26936 19456
rect 26792 18964 26844 18970
rect 26792 18906 26844 18912
rect 26804 17649 26832 18906
rect 26988 18290 27016 21490
rect 26976 18284 27028 18290
rect 26976 18226 27028 18232
rect 26884 17740 26936 17746
rect 26884 17682 26936 17688
rect 26790 17640 26846 17649
rect 26790 17575 26846 17584
rect 26792 17536 26844 17542
rect 26792 17478 26844 17484
rect 26700 17332 26752 17338
rect 26700 17274 26752 17280
rect 26528 16250 26556 16934
rect 26620 16918 26740 16946
rect 26606 16824 26662 16833
rect 26606 16759 26662 16768
rect 26516 16244 26568 16250
rect 26516 16186 26568 16192
rect 26516 16108 26568 16114
rect 26516 16050 26568 16056
rect 26528 14521 26556 16050
rect 26514 14512 26570 14521
rect 26514 14447 26570 14456
rect 26516 13932 26568 13938
rect 26516 13874 26568 13880
rect 26422 13424 26478 13433
rect 26422 13359 26478 13368
rect 26424 13252 26476 13258
rect 26424 13194 26476 13200
rect 26148 12844 26200 12850
rect 26148 12786 26200 12792
rect 26146 12744 26202 12753
rect 26146 12679 26202 12688
rect 26240 12708 26292 12714
rect 26160 12050 26188 12679
rect 26240 12650 26292 12656
rect 26252 12238 26280 12650
rect 26332 12640 26384 12646
rect 26332 12582 26384 12588
rect 26344 12442 26372 12582
rect 26332 12436 26384 12442
rect 26332 12378 26384 12384
rect 26240 12232 26292 12238
rect 26240 12174 26292 12180
rect 26160 12022 26280 12050
rect 25870 9687 25926 9696
rect 25976 9710 26096 9738
rect 25780 9580 25832 9586
rect 25780 9522 25832 9528
rect 25780 8560 25832 8566
rect 25780 8502 25832 8508
rect 25688 5704 25740 5710
rect 25688 5646 25740 5652
rect 25686 5400 25742 5409
rect 25686 5335 25742 5344
rect 25700 5166 25728 5335
rect 25688 5160 25740 5166
rect 25688 5102 25740 5108
rect 25792 4758 25820 8502
rect 25780 4752 25832 4758
rect 25780 4694 25832 4700
rect 25884 3942 25912 9687
rect 25976 7886 26004 9710
rect 26056 9580 26108 9586
rect 26056 9522 26108 9528
rect 26068 9178 26096 9522
rect 26056 9172 26108 9178
rect 26056 9114 26108 9120
rect 26056 8560 26108 8566
rect 26056 8502 26108 8508
rect 25964 7880 26016 7886
rect 25964 7822 26016 7828
rect 25962 7712 26018 7721
rect 25962 7647 26018 7656
rect 25976 7546 26004 7647
rect 25964 7540 26016 7546
rect 25964 7482 26016 7488
rect 25964 6384 26016 6390
rect 26068 6361 26096 8502
rect 26148 8492 26200 8498
rect 26148 8434 26200 8440
rect 26160 8090 26188 8434
rect 26148 8084 26200 8090
rect 26148 8026 26200 8032
rect 26252 7993 26280 12022
rect 26344 11558 26372 12378
rect 26332 11552 26384 11558
rect 26332 11494 26384 11500
rect 26344 11218 26372 11494
rect 26436 11354 26464 13194
rect 26424 11348 26476 11354
rect 26424 11290 26476 11296
rect 26332 11212 26384 11218
rect 26332 11154 26384 11160
rect 26332 11076 26384 11082
rect 26332 11018 26384 11024
rect 26344 10810 26372 11018
rect 26332 10804 26384 10810
rect 26332 10746 26384 10752
rect 26332 10464 26384 10470
rect 26332 10406 26384 10412
rect 26238 7984 26294 7993
rect 26238 7919 26294 7928
rect 26148 7472 26200 7478
rect 26148 7414 26200 7420
rect 26160 7342 26188 7414
rect 26148 7336 26200 7342
rect 26148 7278 26200 7284
rect 26240 7200 26292 7206
rect 26240 7142 26292 7148
rect 26252 7002 26280 7142
rect 26240 6996 26292 7002
rect 26240 6938 26292 6944
rect 26240 6452 26292 6458
rect 26240 6394 26292 6400
rect 25964 6326 26016 6332
rect 26054 6352 26110 6361
rect 25976 6118 26004 6326
rect 26054 6287 26110 6296
rect 25964 6112 26016 6118
rect 25964 6054 26016 6060
rect 25872 3936 25924 3942
rect 25872 3878 25924 3884
rect 25884 3738 25912 3878
rect 25872 3732 25924 3738
rect 25872 3674 25924 3680
rect 25596 3664 25648 3670
rect 25596 3606 25648 3612
rect 25976 3466 26004 6054
rect 26148 5092 26200 5098
rect 26148 5034 26200 5040
rect 26160 4826 26188 5034
rect 26148 4820 26200 4826
rect 26148 4762 26200 4768
rect 26252 4298 26280 6394
rect 26160 4282 26280 4298
rect 26148 4276 26280 4282
rect 26200 4270 26280 4276
rect 26148 4218 26200 4224
rect 26240 4208 26292 4214
rect 26240 4150 26292 4156
rect 26252 3913 26280 4150
rect 26344 4146 26372 10406
rect 26424 9648 26476 9654
rect 26424 9590 26476 9596
rect 26436 8838 26464 9590
rect 26424 8832 26476 8838
rect 26424 8774 26476 8780
rect 26332 4140 26384 4146
rect 26332 4082 26384 4088
rect 26238 3904 26294 3913
rect 26238 3839 26294 3848
rect 26148 3732 26200 3738
rect 26148 3674 26200 3680
rect 25964 3460 26016 3466
rect 25964 3402 26016 3408
rect 26160 2854 26188 3674
rect 26436 3466 26464 8774
rect 26528 8514 26556 13874
rect 26620 12889 26648 16759
rect 26606 12880 26662 12889
rect 26606 12815 26662 12824
rect 26608 12776 26660 12782
rect 26608 12718 26660 12724
rect 26620 12170 26648 12718
rect 26608 12164 26660 12170
rect 26608 12106 26660 12112
rect 26608 11892 26660 11898
rect 26608 11834 26660 11840
rect 26620 8906 26648 11834
rect 26712 11762 26740 16918
rect 26804 15609 26832 17478
rect 26896 15706 26924 17682
rect 26976 17332 27028 17338
rect 26976 17274 27028 17280
rect 26884 15700 26936 15706
rect 26884 15642 26936 15648
rect 26790 15600 26846 15609
rect 26790 15535 26846 15544
rect 26792 14068 26844 14074
rect 26792 14010 26844 14016
rect 26700 11756 26752 11762
rect 26700 11698 26752 11704
rect 26700 9988 26752 9994
rect 26700 9930 26752 9936
rect 26712 9178 26740 9930
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26700 8968 26752 8974
rect 26700 8910 26752 8916
rect 26608 8900 26660 8906
rect 26608 8842 26660 8848
rect 26528 8486 26648 8514
rect 26516 8356 26568 8362
rect 26516 8298 26568 8304
rect 26424 3460 26476 3466
rect 26424 3402 26476 3408
rect 25964 2848 26016 2854
rect 25964 2790 26016 2796
rect 26148 2848 26200 2854
rect 26148 2790 26200 2796
rect 25976 800 26004 2790
rect 26528 800 26556 8298
rect 26620 3670 26648 8486
rect 26712 7886 26740 8910
rect 26804 8498 26832 14010
rect 26884 13796 26936 13802
rect 26884 13738 26936 13744
rect 26896 13530 26924 13738
rect 26884 13524 26936 13530
rect 26884 13466 26936 13472
rect 26896 11218 26924 13466
rect 26884 11212 26936 11218
rect 26884 11154 26936 11160
rect 26884 9920 26936 9926
rect 26884 9862 26936 9868
rect 26896 8838 26924 9862
rect 26884 8832 26936 8838
rect 26884 8774 26936 8780
rect 26792 8492 26844 8498
rect 26792 8434 26844 8440
rect 26896 8378 26924 8774
rect 26804 8350 26924 8378
rect 26988 8378 27016 17274
rect 27080 12753 27108 24550
rect 27160 24404 27212 24410
rect 27160 24346 27212 24352
rect 27172 23798 27200 24346
rect 27160 23792 27212 23798
rect 27160 23734 27212 23740
rect 27160 22636 27212 22642
rect 27160 22578 27212 22584
rect 27172 22234 27200 22578
rect 27160 22228 27212 22234
rect 27160 22170 27212 22176
rect 27264 19854 27292 25214
rect 27356 20602 27384 28494
rect 27804 28008 27856 28014
rect 27804 27950 27856 27956
rect 27620 27668 27672 27674
rect 27620 27610 27672 27616
rect 27528 24608 27580 24614
rect 27528 24550 27580 24556
rect 27436 23588 27488 23594
rect 27436 23530 27488 23536
rect 27344 20596 27396 20602
rect 27344 20538 27396 20544
rect 27252 19848 27304 19854
rect 27252 19790 27304 19796
rect 27250 19544 27306 19553
rect 27250 19479 27306 19488
rect 27264 18970 27292 19479
rect 27252 18964 27304 18970
rect 27252 18906 27304 18912
rect 27344 18284 27396 18290
rect 27344 18226 27396 18232
rect 27252 18216 27304 18222
rect 27252 18158 27304 18164
rect 27160 18080 27212 18086
rect 27160 18022 27212 18028
rect 27066 12744 27122 12753
rect 27066 12679 27122 12688
rect 27068 12640 27120 12646
rect 27068 12582 27120 12588
rect 27080 11762 27108 12582
rect 27068 11756 27120 11762
rect 27068 11698 27120 11704
rect 27172 9602 27200 18022
rect 27264 11744 27292 18158
rect 27356 11898 27384 18226
rect 27448 12306 27476 23530
rect 27540 12646 27568 24550
rect 27528 12640 27580 12646
rect 27528 12582 27580 12588
rect 27526 12472 27582 12481
rect 27632 12442 27660 27610
rect 27712 26580 27764 26586
rect 27712 26522 27764 26528
rect 27526 12407 27582 12416
rect 27620 12436 27672 12442
rect 27436 12300 27488 12306
rect 27436 12242 27488 12248
rect 27436 12096 27488 12102
rect 27436 12038 27488 12044
rect 27344 11892 27396 11898
rect 27344 11834 27396 11840
rect 27264 11716 27384 11744
rect 27250 11656 27306 11665
rect 27250 11591 27252 11600
rect 27304 11591 27306 11600
rect 27252 11562 27304 11568
rect 27252 11348 27304 11354
rect 27252 11290 27304 11296
rect 27080 9574 27200 9602
rect 27080 9450 27108 9574
rect 27160 9512 27212 9518
rect 27160 9454 27212 9460
rect 27068 9444 27120 9450
rect 27068 9386 27120 9392
rect 27172 8974 27200 9454
rect 27160 8968 27212 8974
rect 27160 8910 27212 8916
rect 26988 8350 27108 8378
rect 26700 7880 26752 7886
rect 26700 7822 26752 7828
rect 26700 7404 26752 7410
rect 26700 7346 26752 7352
rect 26712 4554 26740 7346
rect 26700 4548 26752 4554
rect 26700 4490 26752 4496
rect 26804 4214 26832 8350
rect 26976 8288 27028 8294
rect 26976 8230 27028 8236
rect 26988 7750 27016 8230
rect 26976 7744 27028 7750
rect 26976 7686 27028 7692
rect 26884 7472 26936 7478
rect 26884 7414 26936 7420
rect 26896 5574 26924 7414
rect 26884 5568 26936 5574
rect 26884 5510 26936 5516
rect 26988 5302 27016 7686
rect 27080 7274 27108 8350
rect 27172 7886 27200 8910
rect 27264 8566 27292 11290
rect 27356 9722 27384 11716
rect 27344 9716 27396 9722
rect 27344 9658 27396 9664
rect 27356 9042 27384 9658
rect 27344 9036 27396 9042
rect 27344 8978 27396 8984
rect 27344 8628 27396 8634
rect 27344 8570 27396 8576
rect 27252 8560 27304 8566
rect 27252 8502 27304 8508
rect 27252 8424 27304 8430
rect 27252 8366 27304 8372
rect 27160 7880 27212 7886
rect 27160 7822 27212 7828
rect 27160 7540 27212 7546
rect 27160 7482 27212 7488
rect 27068 7268 27120 7274
rect 27068 7210 27120 7216
rect 27172 6458 27200 7482
rect 27160 6452 27212 6458
rect 27160 6394 27212 6400
rect 26976 5296 27028 5302
rect 26976 5238 27028 5244
rect 26884 5160 26936 5166
rect 26884 5102 26936 5108
rect 26976 5160 27028 5166
rect 26976 5102 27028 5108
rect 26896 5030 26924 5102
rect 26884 5024 26936 5030
rect 26884 4966 26936 4972
rect 26896 4826 26924 4966
rect 26884 4820 26936 4826
rect 26884 4762 26936 4768
rect 26988 4554 27016 5102
rect 27160 4616 27212 4622
rect 27160 4558 27212 4564
rect 26976 4548 27028 4554
rect 26976 4490 27028 4496
rect 26884 4276 26936 4282
rect 26884 4218 26936 4224
rect 26792 4208 26844 4214
rect 26792 4150 26844 4156
rect 26608 3664 26660 3670
rect 26608 3606 26660 3612
rect 26896 3398 26924 4218
rect 27172 3534 27200 4558
rect 27160 3528 27212 3534
rect 27160 3470 27212 3476
rect 26884 3392 26936 3398
rect 26884 3334 26936 3340
rect 26896 3194 26924 3334
rect 26884 3188 26936 3194
rect 26884 3130 26936 3136
rect 27264 2922 27292 8366
rect 27356 7585 27384 8570
rect 27342 7576 27398 7585
rect 27342 7511 27398 7520
rect 27344 7404 27396 7410
rect 27344 7346 27396 7352
rect 27356 7002 27384 7346
rect 27448 7206 27476 12038
rect 27540 7546 27568 12407
rect 27620 12378 27672 12384
rect 27620 12300 27672 12306
rect 27620 12242 27672 12248
rect 27632 11354 27660 12242
rect 27620 11348 27672 11354
rect 27620 11290 27672 11296
rect 27620 9376 27672 9382
rect 27620 9318 27672 9324
rect 27528 7540 27580 7546
rect 27528 7482 27580 7488
rect 27526 7304 27582 7313
rect 27526 7239 27582 7248
rect 27436 7200 27488 7206
rect 27436 7142 27488 7148
rect 27344 6996 27396 7002
rect 27344 6938 27396 6944
rect 27342 6488 27398 6497
rect 27342 6423 27344 6432
rect 27396 6423 27398 6432
rect 27344 6394 27396 6400
rect 27448 6118 27476 7142
rect 27436 6112 27488 6118
rect 27436 6054 27488 6060
rect 27344 5568 27396 5574
rect 27344 5510 27396 5516
rect 27356 3126 27384 5510
rect 27540 4010 27568 7239
rect 27528 4004 27580 4010
rect 27528 3946 27580 3952
rect 27344 3120 27396 3126
rect 27344 3062 27396 3068
rect 27252 2916 27304 2922
rect 27252 2858 27304 2864
rect 27252 2304 27304 2310
rect 27252 2246 27304 2252
rect 27264 2106 27292 2246
rect 27252 2100 27304 2106
rect 27252 2042 27304 2048
rect 27068 2032 27120 2038
rect 27068 1974 27120 1980
rect 27080 800 27108 1974
rect 27632 800 27660 9318
rect 27724 5710 27752 26522
rect 27816 10742 27844 27950
rect 27988 24812 28040 24818
rect 27988 24754 28040 24760
rect 27896 12436 27948 12442
rect 27896 12378 27948 12384
rect 27804 10736 27856 10742
rect 27804 10678 27856 10684
rect 27908 6186 27936 12378
rect 28000 7818 28028 24754
rect 28080 12640 28132 12646
rect 28080 12582 28132 12588
rect 28092 12102 28120 12582
rect 28080 12096 28132 12102
rect 28080 12038 28132 12044
rect 27988 7812 28040 7818
rect 27988 7754 28040 7760
rect 27896 6180 27948 6186
rect 27896 6122 27948 6128
rect 27712 5704 27764 5710
rect 27712 5646 27764 5652
rect 28172 5636 28224 5642
rect 28172 5578 28224 5584
rect 28184 800 28212 5578
rect 28724 3528 28776 3534
rect 28724 3470 28776 3476
rect 28736 800 28764 3470
rect 29000 2372 29052 2378
rect 29000 2314 29052 2320
rect 29012 800 29040 2314
rect 110 0 166 800
rect 294 0 350 800
rect 570 0 626 800
rect 846 0 902 800
rect 1122 0 1178 800
rect 1398 0 1454 800
rect 1674 0 1730 800
rect 1950 0 2006 800
rect 2226 0 2282 800
rect 2502 0 2558 800
rect 2778 0 2834 800
rect 3054 0 3110 800
rect 3330 0 3386 800
rect 3606 0 3662 800
rect 3882 0 3938 800
rect 4158 0 4214 800
rect 4342 0 4398 800
rect 4618 0 4674 800
rect 4894 0 4950 800
rect 5170 0 5226 800
rect 5446 0 5502 800
rect 5722 0 5778 800
rect 5998 0 6054 800
rect 6274 0 6330 800
rect 6550 0 6606 800
rect 6826 0 6882 800
rect 7102 0 7158 800
rect 7378 0 7434 800
rect 7654 0 7710 800
rect 7930 0 7986 800
rect 8206 0 8262 800
rect 8390 0 8446 800
rect 8666 0 8722 800
rect 8942 0 8998 800
rect 9218 0 9274 800
rect 9494 0 9550 800
rect 9770 0 9826 800
rect 10046 0 10102 800
rect 10322 0 10378 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11150 0 11206 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12530 0 12586 800
rect 12714 0 12770 800
rect 12990 0 13046 800
rect 13266 0 13322 800
rect 13542 0 13598 800
rect 13818 0 13874 800
rect 14094 0 14150 800
rect 14370 0 14426 800
rect 14646 0 14702 800
rect 14922 0 14978 800
rect 15198 0 15254 800
rect 15474 0 15530 800
rect 15750 0 15806 800
rect 16026 0 16082 800
rect 16302 0 16358 800
rect 16578 0 16634 800
rect 16762 0 16818 800
rect 17038 0 17094 800
rect 17314 0 17370 800
rect 17590 0 17646 800
rect 17866 0 17922 800
rect 18142 0 18198 800
rect 18418 0 18474 800
rect 18694 0 18750 800
rect 18970 0 19026 800
rect 19246 0 19302 800
rect 19522 0 19578 800
rect 19798 0 19854 800
rect 20074 0 20130 800
rect 20350 0 20406 800
rect 20626 0 20682 800
rect 20902 0 20958 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 21914 0 21970 800
rect 22190 0 22246 800
rect 22466 0 22522 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23294 0 23350 800
rect 23570 0 23626 800
rect 23846 0 23902 800
rect 24122 0 24178 800
rect 24398 0 24454 800
rect 24674 0 24730 800
rect 24950 0 25006 800
rect 25134 0 25190 800
rect 25410 0 25466 800
rect 25686 0 25742 800
rect 25962 0 26018 800
rect 26238 0 26294 800
rect 26514 0 26570 800
rect 26790 0 26846 800
rect 27066 0 27122 800
rect 27342 0 27398 800
rect 27618 0 27674 800
rect 27894 0 27950 800
rect 28170 0 28226 800
rect 28446 0 28502 800
rect 28722 0 28778 800
rect 28998 0 29054 800
<< via2 >>
rect 5448 28858 5504 28860
rect 5528 28858 5584 28860
rect 5608 28858 5664 28860
rect 5688 28858 5744 28860
rect 5448 28806 5494 28858
rect 5494 28806 5504 28858
rect 5528 28806 5558 28858
rect 5558 28806 5570 28858
rect 5570 28806 5584 28858
rect 5608 28806 5622 28858
rect 5622 28806 5634 28858
rect 5634 28806 5664 28858
rect 5688 28806 5698 28858
rect 5698 28806 5744 28858
rect 5448 28804 5504 28806
rect 5528 28804 5584 28806
rect 5608 28804 5664 28806
rect 5688 28804 5744 28806
rect 14434 28858 14490 28860
rect 14514 28858 14570 28860
rect 14594 28858 14650 28860
rect 14674 28858 14730 28860
rect 14434 28806 14480 28858
rect 14480 28806 14490 28858
rect 14514 28806 14544 28858
rect 14544 28806 14556 28858
rect 14556 28806 14570 28858
rect 14594 28806 14608 28858
rect 14608 28806 14620 28858
rect 14620 28806 14650 28858
rect 14674 28806 14684 28858
rect 14684 28806 14730 28858
rect 14434 28804 14490 28806
rect 14514 28804 14570 28806
rect 14594 28804 14650 28806
rect 14674 28804 14730 28806
rect 23419 28858 23475 28860
rect 23499 28858 23555 28860
rect 23579 28858 23635 28860
rect 23659 28858 23715 28860
rect 23419 28806 23465 28858
rect 23465 28806 23475 28858
rect 23499 28806 23529 28858
rect 23529 28806 23541 28858
rect 23541 28806 23555 28858
rect 23579 28806 23593 28858
rect 23593 28806 23605 28858
rect 23605 28806 23635 28858
rect 23659 28806 23669 28858
rect 23669 28806 23715 28858
rect 23419 28804 23475 28806
rect 23499 28804 23555 28806
rect 23579 28804 23635 28806
rect 23659 28804 23715 28806
rect 110 3440 166 3496
rect 1122 3576 1178 3632
rect 1398 6296 1454 6352
rect 1858 18808 1914 18864
rect 1858 15544 1914 15600
rect 1674 8880 1730 8936
rect 2686 23024 2742 23080
rect 2502 22344 2558 22400
rect 2226 20712 2282 20768
rect 2594 21800 2650 21856
rect 2686 20984 2742 21040
rect 2594 20168 2650 20224
rect 2502 19896 2558 19952
rect 2686 19352 2742 19408
rect 2594 19216 2650 19272
rect 2686 19080 2742 19136
rect 2686 18708 2688 18728
rect 2688 18708 2740 18728
rect 2740 18708 2742 18728
rect 2686 18672 2742 18708
rect 3054 26288 3110 26344
rect 2870 21936 2926 21992
rect 2870 20440 2926 20496
rect 2410 15680 2466 15736
rect 2226 8880 2282 8936
rect 2778 16224 2834 16280
rect 2686 15408 2742 15464
rect 2042 4256 2098 4312
rect 1306 2760 1362 2816
rect 3238 21528 3294 21584
rect 3146 20884 3148 20904
rect 3148 20884 3200 20904
rect 3200 20884 3202 20904
rect 3146 20848 3202 20884
rect 3238 20748 3240 20768
rect 3240 20748 3292 20768
rect 3292 20748 3294 20768
rect 3238 20712 3294 20748
rect 2686 12688 2742 12744
rect 2962 13640 3018 13696
rect 2962 12008 3018 12064
rect 3146 18944 3202 19000
rect 3146 18828 3202 18864
rect 3146 18808 3148 18828
rect 3148 18808 3200 18828
rect 3200 18808 3202 18828
rect 3146 14184 3202 14240
rect 3054 9968 3110 10024
rect 3054 6840 3110 6896
rect 2778 5344 2834 5400
rect 2962 5616 3018 5672
rect 2870 3168 2926 3224
rect 3238 13504 3294 13560
rect 3606 22752 3662 22808
rect 3422 18672 3478 18728
rect 3606 20304 3662 20360
rect 3606 19760 3662 19816
rect 3606 19660 3608 19680
rect 3608 19660 3660 19680
rect 3660 19660 3662 19680
rect 3606 19624 3662 19660
rect 3606 19508 3662 19544
rect 3606 19488 3608 19508
rect 3608 19488 3660 19508
rect 3660 19488 3662 19508
rect 3422 12824 3478 12880
rect 3606 12960 3662 13016
rect 3238 6840 3294 6896
rect 3330 6432 3386 6488
rect 3330 3168 3386 3224
rect 4434 25880 4490 25936
rect 4250 23704 4306 23760
rect 4526 25472 4582 25528
rect 4342 22888 4398 22944
rect 4250 22752 4306 22808
rect 4158 22616 4214 22672
rect 3974 21664 4030 21720
rect 3882 18264 3938 18320
rect 3882 15272 3938 15328
rect 3882 14320 3938 14376
rect 4158 20304 4214 20360
rect 4158 20168 4214 20224
rect 4066 18536 4122 18592
rect 4066 18400 4122 18456
rect 4250 18672 4306 18728
rect 4250 18128 4306 18184
rect 4526 22344 4582 22400
rect 5448 27770 5504 27772
rect 5528 27770 5584 27772
rect 5608 27770 5664 27772
rect 5688 27770 5744 27772
rect 5448 27718 5494 27770
rect 5494 27718 5504 27770
rect 5528 27718 5558 27770
rect 5558 27718 5570 27770
rect 5570 27718 5584 27770
rect 5608 27718 5622 27770
rect 5622 27718 5634 27770
rect 5634 27718 5664 27770
rect 5688 27718 5698 27770
rect 5698 27718 5744 27770
rect 5448 27716 5504 27718
rect 5528 27716 5584 27718
rect 5608 27716 5664 27718
rect 5688 27716 5744 27718
rect 5446 26832 5502 26888
rect 5448 26682 5504 26684
rect 5528 26682 5584 26684
rect 5608 26682 5664 26684
rect 5688 26682 5744 26684
rect 5448 26630 5494 26682
rect 5494 26630 5504 26682
rect 5528 26630 5558 26682
rect 5558 26630 5570 26682
rect 5570 26630 5584 26682
rect 5608 26630 5622 26682
rect 5622 26630 5634 26682
rect 5634 26630 5664 26682
rect 5688 26630 5698 26682
rect 5698 26630 5744 26682
rect 5448 26628 5504 26630
rect 5528 26628 5584 26630
rect 5608 26628 5664 26630
rect 5688 26628 5744 26630
rect 5262 26016 5318 26072
rect 5078 25472 5134 25528
rect 6182 27512 6238 27568
rect 5630 25880 5686 25936
rect 5448 25594 5504 25596
rect 5528 25594 5584 25596
rect 5608 25594 5664 25596
rect 5688 25594 5744 25596
rect 5448 25542 5494 25594
rect 5494 25542 5504 25594
rect 5528 25542 5558 25594
rect 5558 25542 5570 25594
rect 5570 25542 5584 25594
rect 5608 25542 5622 25594
rect 5622 25542 5634 25594
rect 5634 25542 5664 25594
rect 5688 25542 5698 25594
rect 5698 25542 5744 25594
rect 5448 25540 5504 25542
rect 5528 25540 5584 25542
rect 5608 25540 5664 25542
rect 5688 25540 5744 25542
rect 5906 25472 5962 25528
rect 5538 24656 5594 24712
rect 5448 24506 5504 24508
rect 5528 24506 5584 24508
rect 5608 24506 5664 24508
rect 5688 24506 5744 24508
rect 5448 24454 5494 24506
rect 5494 24454 5504 24506
rect 5528 24454 5558 24506
rect 5558 24454 5570 24506
rect 5570 24454 5584 24506
rect 5608 24454 5622 24506
rect 5622 24454 5634 24506
rect 5634 24454 5664 24506
rect 5688 24454 5698 24506
rect 5698 24454 5744 24506
rect 5448 24452 5504 24454
rect 5528 24452 5584 24454
rect 5608 24452 5664 24454
rect 5688 24452 5744 24454
rect 5170 23840 5226 23896
rect 4894 22480 4950 22536
rect 5078 21392 5134 21448
rect 4894 21292 4896 21312
rect 4896 21292 4948 21312
rect 4948 21292 4950 21312
rect 4894 21256 4950 21292
rect 4434 19216 4490 19272
rect 4618 18536 4674 18592
rect 4710 17584 4766 17640
rect 3882 13776 3938 13832
rect 4158 12416 4214 12472
rect 4066 12008 4122 12064
rect 3606 6860 3662 6896
rect 3606 6840 3608 6860
rect 3608 6840 3660 6860
rect 3660 6840 3662 6860
rect 3606 5072 3662 5128
rect 3974 8492 4030 8528
rect 3974 8472 3976 8492
rect 3976 8472 4028 8492
rect 4028 8472 4030 8492
rect 3790 5208 3846 5264
rect 4066 7112 4122 7168
rect 3698 3712 3754 3768
rect 4526 12280 4582 12336
rect 4250 8336 4306 8392
rect 4710 12416 4766 12472
rect 4710 12008 4766 12064
rect 5448 23418 5504 23420
rect 5528 23418 5584 23420
rect 5608 23418 5664 23420
rect 5688 23418 5744 23420
rect 5448 23366 5494 23418
rect 5494 23366 5504 23418
rect 5528 23366 5558 23418
rect 5558 23366 5570 23418
rect 5570 23366 5584 23418
rect 5608 23366 5622 23418
rect 5622 23366 5634 23418
rect 5634 23366 5664 23418
rect 5688 23366 5698 23418
rect 5698 23366 5744 23418
rect 5448 23364 5504 23366
rect 5528 23364 5584 23366
rect 5608 23364 5664 23366
rect 5688 23364 5744 23366
rect 5814 23024 5870 23080
rect 5446 22752 5502 22808
rect 5262 22480 5318 22536
rect 5448 22330 5504 22332
rect 5528 22330 5584 22332
rect 5608 22330 5664 22332
rect 5688 22330 5744 22332
rect 5448 22278 5494 22330
rect 5494 22278 5504 22330
rect 5528 22278 5558 22330
rect 5558 22278 5570 22330
rect 5570 22278 5584 22330
rect 5608 22278 5622 22330
rect 5622 22278 5634 22330
rect 5634 22278 5664 22330
rect 5688 22278 5698 22330
rect 5698 22278 5744 22330
rect 5448 22276 5504 22278
rect 5528 22276 5584 22278
rect 5608 22276 5664 22278
rect 5688 22276 5744 22278
rect 5448 21242 5504 21244
rect 5528 21242 5584 21244
rect 5608 21242 5664 21244
rect 5688 21242 5744 21244
rect 5448 21190 5494 21242
rect 5494 21190 5504 21242
rect 5528 21190 5558 21242
rect 5558 21190 5570 21242
rect 5570 21190 5584 21242
rect 5608 21190 5622 21242
rect 5622 21190 5634 21242
rect 5634 21190 5664 21242
rect 5688 21190 5698 21242
rect 5698 21190 5744 21242
rect 5448 21188 5504 21190
rect 5528 21188 5584 21190
rect 5608 21188 5664 21190
rect 5688 21188 5744 21190
rect 5354 20576 5410 20632
rect 5262 19080 5318 19136
rect 5448 20154 5504 20156
rect 5528 20154 5584 20156
rect 5608 20154 5664 20156
rect 5688 20154 5744 20156
rect 5448 20102 5494 20154
rect 5494 20102 5504 20154
rect 5528 20102 5558 20154
rect 5558 20102 5570 20154
rect 5570 20102 5584 20154
rect 5608 20102 5622 20154
rect 5622 20102 5634 20154
rect 5634 20102 5664 20154
rect 5688 20102 5698 20154
rect 5698 20102 5744 20154
rect 5448 20100 5504 20102
rect 5528 20100 5584 20102
rect 5608 20100 5664 20102
rect 5688 20100 5744 20102
rect 5448 19066 5504 19068
rect 5528 19066 5584 19068
rect 5608 19066 5664 19068
rect 5688 19066 5744 19068
rect 5448 19014 5494 19066
rect 5494 19014 5504 19066
rect 5528 19014 5558 19066
rect 5558 19014 5570 19066
rect 5570 19014 5584 19066
rect 5608 19014 5622 19066
rect 5622 19014 5634 19066
rect 5634 19014 5664 19066
rect 5688 19014 5698 19066
rect 5698 19014 5744 19066
rect 5448 19012 5504 19014
rect 5528 19012 5584 19014
rect 5608 19012 5664 19014
rect 5688 19012 5744 19014
rect 5538 18300 5540 18320
rect 5540 18300 5592 18320
rect 5592 18300 5594 18320
rect 5538 18264 5594 18300
rect 5446 18128 5502 18184
rect 5448 17978 5504 17980
rect 5528 17978 5584 17980
rect 5608 17978 5664 17980
rect 5688 17978 5744 17980
rect 5448 17926 5494 17978
rect 5494 17926 5504 17978
rect 5528 17926 5558 17978
rect 5558 17926 5570 17978
rect 5570 17926 5584 17978
rect 5608 17926 5622 17978
rect 5622 17926 5634 17978
rect 5634 17926 5664 17978
rect 5688 17926 5698 17978
rect 5698 17926 5744 17978
rect 5448 17924 5504 17926
rect 5528 17924 5584 17926
rect 5608 17924 5664 17926
rect 5688 17924 5744 17926
rect 5262 17312 5318 17368
rect 5906 20304 5962 20360
rect 4894 13232 4950 13288
rect 4802 9832 4858 9888
rect 5170 13232 5226 13288
rect 5078 11600 5134 11656
rect 5078 9696 5134 9752
rect 5078 6840 5134 6896
rect 5448 16890 5504 16892
rect 5528 16890 5584 16892
rect 5608 16890 5664 16892
rect 5688 16890 5744 16892
rect 5448 16838 5494 16890
rect 5494 16838 5504 16890
rect 5528 16838 5558 16890
rect 5558 16838 5570 16890
rect 5570 16838 5584 16890
rect 5608 16838 5622 16890
rect 5622 16838 5634 16890
rect 5634 16838 5664 16890
rect 5688 16838 5698 16890
rect 5698 16838 5744 16890
rect 5448 16836 5504 16838
rect 5528 16836 5584 16838
rect 5608 16836 5664 16838
rect 5688 16836 5744 16838
rect 5448 15802 5504 15804
rect 5528 15802 5584 15804
rect 5608 15802 5664 15804
rect 5688 15802 5744 15804
rect 5448 15750 5494 15802
rect 5494 15750 5504 15802
rect 5528 15750 5558 15802
rect 5558 15750 5570 15802
rect 5570 15750 5584 15802
rect 5608 15750 5622 15802
rect 5622 15750 5634 15802
rect 5634 15750 5664 15802
rect 5688 15750 5698 15802
rect 5698 15750 5744 15802
rect 5448 15748 5504 15750
rect 5528 15748 5584 15750
rect 5608 15748 5664 15750
rect 5688 15748 5744 15750
rect 5448 14714 5504 14716
rect 5528 14714 5584 14716
rect 5608 14714 5664 14716
rect 5688 14714 5744 14716
rect 5448 14662 5494 14714
rect 5494 14662 5504 14714
rect 5528 14662 5558 14714
rect 5558 14662 5570 14714
rect 5570 14662 5584 14714
rect 5608 14662 5622 14714
rect 5622 14662 5634 14714
rect 5634 14662 5664 14714
rect 5688 14662 5698 14714
rect 5698 14662 5744 14714
rect 5448 14660 5504 14662
rect 5528 14660 5584 14662
rect 5608 14660 5664 14662
rect 5688 14660 5744 14662
rect 5448 13626 5504 13628
rect 5528 13626 5584 13628
rect 5608 13626 5664 13628
rect 5688 13626 5744 13628
rect 5448 13574 5494 13626
rect 5494 13574 5504 13626
rect 5528 13574 5558 13626
rect 5558 13574 5570 13626
rect 5570 13574 5584 13626
rect 5608 13574 5622 13626
rect 5622 13574 5634 13626
rect 5634 13574 5664 13626
rect 5688 13574 5698 13626
rect 5698 13574 5744 13626
rect 5448 13572 5504 13574
rect 5528 13572 5584 13574
rect 5608 13572 5664 13574
rect 5688 13572 5744 13574
rect 5262 12552 5318 12608
rect 5262 12416 5318 12472
rect 5538 12860 5540 12880
rect 5540 12860 5592 12880
rect 5592 12860 5594 12880
rect 5538 12824 5594 12860
rect 5448 12538 5504 12540
rect 5528 12538 5584 12540
rect 5608 12538 5664 12540
rect 5688 12538 5744 12540
rect 5448 12486 5494 12538
rect 5494 12486 5504 12538
rect 5528 12486 5558 12538
rect 5558 12486 5570 12538
rect 5570 12486 5584 12538
rect 5608 12486 5622 12538
rect 5622 12486 5634 12538
rect 5634 12486 5664 12538
rect 5688 12486 5698 12538
rect 5698 12486 5744 12538
rect 5448 12484 5504 12486
rect 5528 12484 5584 12486
rect 5608 12484 5664 12486
rect 5688 12484 5744 12486
rect 6090 26988 6146 27024
rect 6090 26968 6092 26988
rect 6092 26968 6144 26988
rect 6144 26968 6146 26988
rect 6366 26016 6422 26072
rect 6182 24556 6184 24576
rect 6184 24556 6236 24576
rect 6236 24556 6238 24576
rect 6182 24520 6238 24556
rect 6458 25472 6514 25528
rect 6182 20576 6238 20632
rect 5448 11450 5504 11452
rect 5528 11450 5584 11452
rect 5608 11450 5664 11452
rect 5688 11450 5744 11452
rect 5448 11398 5494 11450
rect 5494 11398 5504 11450
rect 5528 11398 5558 11450
rect 5558 11398 5570 11450
rect 5570 11398 5584 11450
rect 5608 11398 5622 11450
rect 5622 11398 5634 11450
rect 5634 11398 5664 11450
rect 5688 11398 5698 11450
rect 5698 11398 5744 11450
rect 5448 11396 5504 11398
rect 5528 11396 5584 11398
rect 5608 11396 5664 11398
rect 5688 11396 5744 11398
rect 5448 10362 5504 10364
rect 5528 10362 5584 10364
rect 5608 10362 5664 10364
rect 5688 10362 5744 10364
rect 5448 10310 5494 10362
rect 5494 10310 5504 10362
rect 5528 10310 5558 10362
rect 5558 10310 5570 10362
rect 5570 10310 5584 10362
rect 5608 10310 5622 10362
rect 5622 10310 5634 10362
rect 5634 10310 5664 10362
rect 5688 10310 5698 10362
rect 5698 10310 5744 10362
rect 5448 10308 5504 10310
rect 5528 10308 5584 10310
rect 5608 10308 5664 10310
rect 5688 10308 5744 10310
rect 5448 9274 5504 9276
rect 5528 9274 5584 9276
rect 5608 9274 5664 9276
rect 5688 9274 5744 9276
rect 5448 9222 5494 9274
rect 5494 9222 5504 9274
rect 5528 9222 5558 9274
rect 5558 9222 5570 9274
rect 5570 9222 5584 9274
rect 5608 9222 5622 9274
rect 5622 9222 5634 9274
rect 5634 9222 5664 9274
rect 5688 9222 5698 9274
rect 5698 9222 5744 9274
rect 5448 9220 5504 9222
rect 5528 9220 5584 9222
rect 5608 9220 5664 9222
rect 5688 9220 5744 9222
rect 5448 8186 5504 8188
rect 5528 8186 5584 8188
rect 5608 8186 5664 8188
rect 5688 8186 5744 8188
rect 5448 8134 5494 8186
rect 5494 8134 5504 8186
rect 5528 8134 5558 8186
rect 5558 8134 5570 8186
rect 5570 8134 5584 8186
rect 5608 8134 5622 8186
rect 5622 8134 5634 8186
rect 5634 8134 5664 8186
rect 5688 8134 5698 8186
rect 5698 8134 5744 8186
rect 5448 8132 5504 8134
rect 5528 8132 5584 8134
rect 5608 8132 5664 8134
rect 5688 8132 5744 8134
rect 5448 7098 5504 7100
rect 5528 7098 5584 7100
rect 5608 7098 5664 7100
rect 5688 7098 5744 7100
rect 5448 7046 5494 7098
rect 5494 7046 5504 7098
rect 5528 7046 5558 7098
rect 5558 7046 5570 7098
rect 5570 7046 5584 7098
rect 5608 7046 5622 7098
rect 5622 7046 5634 7098
rect 5634 7046 5664 7098
rect 5688 7046 5698 7098
rect 5698 7046 5744 7098
rect 5448 7044 5504 7046
rect 5528 7044 5584 7046
rect 5608 7044 5664 7046
rect 5688 7044 5744 7046
rect 5906 6704 5962 6760
rect 5448 6010 5504 6012
rect 5528 6010 5584 6012
rect 5608 6010 5664 6012
rect 5688 6010 5744 6012
rect 5448 5958 5494 6010
rect 5494 5958 5504 6010
rect 5528 5958 5558 6010
rect 5558 5958 5570 6010
rect 5570 5958 5584 6010
rect 5608 5958 5622 6010
rect 5622 5958 5634 6010
rect 5634 5958 5664 6010
rect 5688 5958 5698 6010
rect 5698 5958 5744 6010
rect 5448 5956 5504 5958
rect 5528 5956 5584 5958
rect 5608 5956 5664 5958
rect 5688 5956 5744 5958
rect 5448 4922 5504 4924
rect 5528 4922 5584 4924
rect 5608 4922 5664 4924
rect 5688 4922 5744 4924
rect 5448 4870 5494 4922
rect 5494 4870 5504 4922
rect 5528 4870 5558 4922
rect 5558 4870 5570 4922
rect 5570 4870 5584 4922
rect 5608 4870 5622 4922
rect 5622 4870 5634 4922
rect 5634 4870 5664 4922
rect 5688 4870 5698 4922
rect 5698 4870 5744 4922
rect 5448 4868 5504 4870
rect 5528 4868 5584 4870
rect 5608 4868 5664 4870
rect 5688 4868 5744 4870
rect 5262 3712 5318 3768
rect 5262 3168 5318 3224
rect 5448 3834 5504 3836
rect 5528 3834 5584 3836
rect 5608 3834 5664 3836
rect 5688 3834 5744 3836
rect 5448 3782 5494 3834
rect 5494 3782 5504 3834
rect 5528 3782 5558 3834
rect 5558 3782 5570 3834
rect 5570 3782 5584 3834
rect 5608 3782 5622 3834
rect 5622 3782 5634 3834
rect 5634 3782 5664 3834
rect 5688 3782 5698 3834
rect 5698 3782 5744 3834
rect 5448 3780 5504 3782
rect 5528 3780 5584 3782
rect 5608 3780 5664 3782
rect 5688 3780 5744 3782
rect 5446 3576 5502 3632
rect 5448 2746 5504 2748
rect 5528 2746 5584 2748
rect 5608 2746 5664 2748
rect 5688 2746 5744 2748
rect 5448 2694 5494 2746
rect 5494 2694 5504 2746
rect 5528 2694 5558 2746
rect 5558 2694 5570 2746
rect 5570 2694 5584 2746
rect 5608 2694 5622 2746
rect 5622 2694 5634 2746
rect 5634 2694 5664 2746
rect 5688 2694 5698 2746
rect 5698 2694 5744 2746
rect 5448 2692 5504 2694
rect 5528 2692 5584 2694
rect 5608 2692 5664 2694
rect 5688 2692 5744 2694
rect 5722 2488 5778 2544
rect 6642 21428 6644 21448
rect 6644 21428 6696 21448
rect 6696 21428 6698 21448
rect 6642 21392 6698 21428
rect 6918 24692 6920 24712
rect 6920 24692 6972 24712
rect 6972 24692 6974 24712
rect 6918 24656 6974 24692
rect 6918 24556 6920 24576
rect 6920 24556 6972 24576
rect 6972 24556 6974 24576
rect 6918 24520 6974 24556
rect 6366 11872 6422 11928
rect 6274 9968 6330 10024
rect 7010 19352 7066 19408
rect 6918 18844 6920 18864
rect 6920 18844 6972 18864
rect 6972 18844 6974 18864
rect 6918 18808 6974 18844
rect 6918 18692 6974 18728
rect 6918 18672 6920 18692
rect 6920 18672 6972 18692
rect 6972 18672 6974 18692
rect 6826 15544 6882 15600
rect 6550 12552 6606 12608
rect 6550 12280 6606 12336
rect 6826 13912 6882 13968
rect 7010 18400 7066 18456
rect 6734 12280 6790 12336
rect 6366 8472 6422 8528
rect 6550 8472 6606 8528
rect 6826 12008 6882 12064
rect 7010 12416 7066 12472
rect 6918 9968 6974 10024
rect 6918 8472 6974 8528
rect 6550 4392 6606 4448
rect 6182 3848 6238 3904
rect 6274 3168 6330 3224
rect 7010 6724 7066 6760
rect 7010 6704 7012 6724
rect 7012 6704 7064 6724
rect 7064 6704 7066 6724
rect 6826 3168 6882 3224
rect 7010 2896 7066 2952
rect 7470 27512 7526 27568
rect 7194 26988 7250 27024
rect 7194 26968 7196 26988
rect 7196 26968 7248 26988
rect 7248 26968 7250 26988
rect 8666 27376 8722 27432
rect 7562 21800 7618 21856
rect 7562 21664 7618 21720
rect 7470 21564 7472 21584
rect 7472 21564 7524 21584
rect 7524 21564 7526 21584
rect 7470 21528 7526 21564
rect 7194 20576 7250 20632
rect 7286 20304 7342 20360
rect 7930 21800 7986 21856
rect 7378 19624 7434 19680
rect 7286 19080 7342 19136
rect 7378 17040 7434 17096
rect 7194 12280 7250 12336
rect 7194 12008 7250 12064
rect 7378 12588 7380 12608
rect 7380 12588 7432 12608
rect 7432 12588 7434 12608
rect 7378 12552 7434 12588
rect 7378 12416 7434 12472
rect 7378 12280 7434 12336
rect 8298 21800 8354 21856
rect 9941 28314 9997 28316
rect 10021 28314 10077 28316
rect 10101 28314 10157 28316
rect 10181 28314 10237 28316
rect 9941 28262 9987 28314
rect 9987 28262 9997 28314
rect 10021 28262 10051 28314
rect 10051 28262 10063 28314
rect 10063 28262 10077 28314
rect 10101 28262 10115 28314
rect 10115 28262 10127 28314
rect 10127 28262 10157 28314
rect 10181 28262 10191 28314
rect 10191 28262 10237 28314
rect 9941 28260 9997 28262
rect 10021 28260 10077 28262
rect 10101 28260 10157 28262
rect 10181 28260 10237 28262
rect 9941 27226 9997 27228
rect 10021 27226 10077 27228
rect 10101 27226 10157 27228
rect 10181 27226 10237 27228
rect 9941 27174 9987 27226
rect 9987 27174 9997 27226
rect 10021 27174 10051 27226
rect 10051 27174 10063 27226
rect 10063 27174 10077 27226
rect 10101 27174 10115 27226
rect 10115 27174 10127 27226
rect 10127 27174 10157 27226
rect 10181 27174 10191 27226
rect 10191 27174 10237 27226
rect 9941 27172 9997 27174
rect 10021 27172 10077 27174
rect 10101 27172 10157 27174
rect 10181 27172 10237 27174
rect 8666 20576 8722 20632
rect 8942 21800 8998 21856
rect 7930 19896 7986 19952
rect 8114 19896 8170 19952
rect 8114 19372 8170 19408
rect 8114 19352 8116 19372
rect 8116 19352 8168 19372
rect 8168 19352 8170 19372
rect 7838 18944 7894 19000
rect 8206 18536 8262 18592
rect 7930 18420 7986 18456
rect 7930 18400 7932 18420
rect 7932 18400 7984 18420
rect 7984 18400 7986 18420
rect 8022 18264 8078 18320
rect 7930 15020 7986 15056
rect 7930 15000 7932 15020
rect 7932 15000 7984 15020
rect 7984 15000 7986 15020
rect 7654 12416 7710 12472
rect 7930 13232 7986 13288
rect 7838 12688 7894 12744
rect 8666 19488 8722 19544
rect 8482 19080 8538 19136
rect 8758 19216 8814 19272
rect 7746 12280 7802 12336
rect 7654 11092 7656 11112
rect 7656 11092 7708 11112
rect 7708 11092 7710 11112
rect 7654 11056 7710 11092
rect 7286 7384 7342 7440
rect 7286 5344 7342 5400
rect 7562 8472 7618 8528
rect 7378 2896 7434 2952
rect 7746 7248 7802 7304
rect 8574 15000 8630 15056
rect 8850 14728 8906 14784
rect 9941 26138 9997 26140
rect 10021 26138 10077 26140
rect 10101 26138 10157 26140
rect 10181 26138 10237 26140
rect 9941 26086 9987 26138
rect 9987 26086 9997 26138
rect 10021 26086 10051 26138
rect 10051 26086 10063 26138
rect 10063 26086 10077 26138
rect 10101 26086 10115 26138
rect 10115 26086 10127 26138
rect 10127 26086 10157 26138
rect 10181 26086 10191 26138
rect 10191 26086 10237 26138
rect 9941 26084 9997 26086
rect 10021 26084 10077 26086
rect 10101 26084 10157 26086
rect 10181 26084 10237 26086
rect 9941 25050 9997 25052
rect 10021 25050 10077 25052
rect 10101 25050 10157 25052
rect 10181 25050 10237 25052
rect 9941 24998 9987 25050
rect 9987 24998 9997 25050
rect 10021 24998 10051 25050
rect 10051 24998 10063 25050
rect 10063 24998 10077 25050
rect 10101 24998 10115 25050
rect 10115 24998 10127 25050
rect 10127 24998 10157 25050
rect 10181 24998 10191 25050
rect 10191 24998 10237 25050
rect 9941 24996 9997 24998
rect 10021 24996 10077 24998
rect 10101 24996 10157 24998
rect 10181 24996 10237 24998
rect 9402 22072 9458 22128
rect 9941 23962 9997 23964
rect 10021 23962 10077 23964
rect 10101 23962 10157 23964
rect 10181 23962 10237 23964
rect 9941 23910 9987 23962
rect 9987 23910 9997 23962
rect 10021 23910 10051 23962
rect 10051 23910 10063 23962
rect 10063 23910 10077 23962
rect 10101 23910 10115 23962
rect 10115 23910 10127 23962
rect 10127 23910 10157 23962
rect 10181 23910 10191 23962
rect 10191 23910 10237 23962
rect 9941 23908 9997 23910
rect 10021 23908 10077 23910
rect 10101 23908 10157 23910
rect 10181 23908 10237 23910
rect 9941 22874 9997 22876
rect 10021 22874 10077 22876
rect 10101 22874 10157 22876
rect 10181 22874 10237 22876
rect 9941 22822 9987 22874
rect 9987 22822 9997 22874
rect 10021 22822 10051 22874
rect 10051 22822 10063 22874
rect 10063 22822 10077 22874
rect 10101 22822 10115 22874
rect 10115 22822 10127 22874
rect 10127 22822 10157 22874
rect 10181 22822 10191 22874
rect 10191 22822 10237 22874
rect 9941 22820 9997 22822
rect 10021 22820 10077 22822
rect 10101 22820 10157 22822
rect 10181 22820 10237 22822
rect 10874 26424 10930 26480
rect 10414 22092 10470 22128
rect 10414 22072 10416 22092
rect 10416 22072 10468 22092
rect 10468 22072 10470 22092
rect 9941 21786 9997 21788
rect 10021 21786 10077 21788
rect 10101 21786 10157 21788
rect 10181 21786 10237 21788
rect 9941 21734 9987 21786
rect 9987 21734 9997 21786
rect 10021 21734 10051 21786
rect 10051 21734 10063 21786
rect 10063 21734 10077 21786
rect 10101 21734 10115 21786
rect 10115 21734 10127 21786
rect 10127 21734 10157 21786
rect 10181 21734 10191 21786
rect 10191 21734 10237 21786
rect 9941 21732 9997 21734
rect 10021 21732 10077 21734
rect 10101 21732 10157 21734
rect 10181 21732 10237 21734
rect 9770 21392 9826 21448
rect 10322 21392 10378 21448
rect 9954 20884 9956 20904
rect 9956 20884 10008 20904
rect 10008 20884 10010 20904
rect 8574 12824 8630 12880
rect 9586 17720 9642 17776
rect 9954 20848 10010 20884
rect 9941 20698 9997 20700
rect 10021 20698 10077 20700
rect 10101 20698 10157 20700
rect 10181 20698 10237 20700
rect 9941 20646 9987 20698
rect 9987 20646 9997 20698
rect 10021 20646 10051 20698
rect 10051 20646 10063 20698
rect 10063 20646 10077 20698
rect 10101 20646 10115 20698
rect 10115 20646 10127 20698
rect 10127 20646 10157 20698
rect 10181 20646 10191 20698
rect 10191 20646 10237 20698
rect 9941 20644 9997 20646
rect 10021 20644 10077 20646
rect 10101 20644 10157 20646
rect 10181 20644 10237 20646
rect 9770 20576 9826 20632
rect 9126 13096 9182 13152
rect 9218 12960 9274 13016
rect 8850 12552 8906 12608
rect 8666 12416 8722 12472
rect 8206 12008 8262 12064
rect 8114 9832 8170 9888
rect 8022 4664 8078 4720
rect 8666 12280 8722 12336
rect 9402 12552 9458 12608
rect 9402 12416 9458 12472
rect 9941 19610 9997 19612
rect 10021 19610 10077 19612
rect 10101 19610 10157 19612
rect 10181 19610 10237 19612
rect 9941 19558 9987 19610
rect 9987 19558 9997 19610
rect 10021 19558 10051 19610
rect 10051 19558 10063 19610
rect 10063 19558 10077 19610
rect 10101 19558 10115 19610
rect 10115 19558 10127 19610
rect 10127 19558 10157 19610
rect 10181 19558 10191 19610
rect 10191 19558 10237 19610
rect 9941 19556 9997 19558
rect 10021 19556 10077 19558
rect 10101 19556 10157 19558
rect 10181 19556 10237 19558
rect 9941 18522 9997 18524
rect 10021 18522 10077 18524
rect 10101 18522 10157 18524
rect 10181 18522 10237 18524
rect 9941 18470 9987 18522
rect 9987 18470 9997 18522
rect 10021 18470 10051 18522
rect 10051 18470 10063 18522
rect 10063 18470 10077 18522
rect 10101 18470 10115 18522
rect 10115 18470 10127 18522
rect 10127 18470 10157 18522
rect 10181 18470 10191 18522
rect 10191 18470 10237 18522
rect 9941 18468 9997 18470
rect 10021 18468 10077 18470
rect 10101 18468 10157 18470
rect 10181 18468 10237 18470
rect 10414 18400 10470 18456
rect 10598 21548 10654 21584
rect 10598 21528 10600 21548
rect 10600 21528 10652 21548
rect 10652 21528 10654 21548
rect 10690 20304 10746 20360
rect 11150 22344 11206 22400
rect 10874 20884 10876 20904
rect 10876 20884 10928 20904
rect 10928 20884 10930 20904
rect 10874 20848 10930 20884
rect 10782 19216 10838 19272
rect 10598 18808 10654 18864
rect 10138 18128 10194 18184
rect 10138 18028 10140 18048
rect 10140 18028 10192 18048
rect 10192 18028 10194 18048
rect 10138 17992 10194 18028
rect 10046 17856 10102 17912
rect 9941 17434 9997 17436
rect 10021 17434 10077 17436
rect 10101 17434 10157 17436
rect 10181 17434 10237 17436
rect 9941 17382 9987 17434
rect 9987 17382 9997 17434
rect 10021 17382 10051 17434
rect 10051 17382 10063 17434
rect 10063 17382 10077 17434
rect 10101 17382 10115 17434
rect 10115 17382 10127 17434
rect 10127 17382 10157 17434
rect 10181 17382 10191 17434
rect 10191 17382 10237 17434
rect 9941 17380 9997 17382
rect 10021 17380 10077 17382
rect 10101 17380 10157 17382
rect 10181 17380 10237 17382
rect 9941 16346 9997 16348
rect 10021 16346 10077 16348
rect 10101 16346 10157 16348
rect 10181 16346 10237 16348
rect 9941 16294 9987 16346
rect 9987 16294 9997 16346
rect 10021 16294 10051 16346
rect 10051 16294 10063 16346
rect 10063 16294 10077 16346
rect 10101 16294 10115 16346
rect 10115 16294 10127 16346
rect 10127 16294 10157 16346
rect 10181 16294 10191 16346
rect 10191 16294 10237 16346
rect 9941 16292 9997 16294
rect 10021 16292 10077 16294
rect 10101 16292 10157 16294
rect 10181 16292 10237 16294
rect 9941 15258 9997 15260
rect 10021 15258 10077 15260
rect 10101 15258 10157 15260
rect 10181 15258 10237 15260
rect 9941 15206 9987 15258
rect 9987 15206 9997 15258
rect 10021 15206 10051 15258
rect 10051 15206 10063 15258
rect 10063 15206 10077 15258
rect 10101 15206 10115 15258
rect 10115 15206 10127 15258
rect 10127 15206 10157 15258
rect 10181 15206 10191 15258
rect 10191 15206 10237 15258
rect 9941 15204 9997 15206
rect 10021 15204 10077 15206
rect 10101 15204 10157 15206
rect 10181 15204 10237 15206
rect 10690 18536 10746 18592
rect 10966 18808 11022 18864
rect 10874 18692 10930 18728
rect 10874 18672 10876 18692
rect 10876 18672 10928 18692
rect 10928 18672 10930 18692
rect 10966 18536 11022 18592
rect 10690 17176 10746 17232
rect 9862 14592 9918 14648
rect 9941 14170 9997 14172
rect 10021 14170 10077 14172
rect 10101 14170 10157 14172
rect 10181 14170 10237 14172
rect 9941 14118 9987 14170
rect 9987 14118 9997 14170
rect 10021 14118 10051 14170
rect 10051 14118 10063 14170
rect 10063 14118 10077 14170
rect 10101 14118 10115 14170
rect 10115 14118 10127 14170
rect 10127 14118 10157 14170
rect 10181 14118 10191 14170
rect 10191 14118 10237 14170
rect 9941 14116 9997 14118
rect 10021 14116 10077 14118
rect 10101 14116 10157 14118
rect 10181 14116 10237 14118
rect 9586 12280 9642 12336
rect 9941 13082 9997 13084
rect 10021 13082 10077 13084
rect 10101 13082 10157 13084
rect 10181 13082 10237 13084
rect 9941 13030 9987 13082
rect 9987 13030 9997 13082
rect 10021 13030 10051 13082
rect 10051 13030 10063 13082
rect 10063 13030 10077 13082
rect 10101 13030 10115 13082
rect 10115 13030 10127 13082
rect 10127 13030 10157 13082
rect 10181 13030 10191 13082
rect 10191 13030 10237 13082
rect 9941 13028 9997 13030
rect 10021 13028 10077 13030
rect 10101 13028 10157 13030
rect 10181 13028 10237 13030
rect 10690 14320 10746 14376
rect 10874 14048 10930 14104
rect 10414 12688 10470 12744
rect 9586 11736 9642 11792
rect 9310 11192 9366 11248
rect 8942 10920 8998 10976
rect 8850 10784 8906 10840
rect 8942 6316 8998 6352
rect 8942 6296 8944 6316
rect 8944 6296 8996 6316
rect 8996 6296 8998 6316
rect 9941 11994 9997 11996
rect 10021 11994 10077 11996
rect 10101 11994 10157 11996
rect 10181 11994 10237 11996
rect 9941 11942 9987 11994
rect 9987 11942 9997 11994
rect 10021 11942 10051 11994
rect 10051 11942 10063 11994
rect 10063 11942 10077 11994
rect 10101 11942 10115 11994
rect 10115 11942 10127 11994
rect 10127 11942 10157 11994
rect 10181 11942 10191 11994
rect 10191 11942 10237 11994
rect 9941 11940 9997 11942
rect 10021 11940 10077 11942
rect 10101 11940 10157 11942
rect 10181 11940 10237 11942
rect 9770 11736 9826 11792
rect 9941 10906 9997 10908
rect 10021 10906 10077 10908
rect 10101 10906 10157 10908
rect 10181 10906 10237 10908
rect 9941 10854 9987 10906
rect 9987 10854 9997 10906
rect 10021 10854 10051 10906
rect 10051 10854 10063 10906
rect 10063 10854 10077 10906
rect 10101 10854 10115 10906
rect 10115 10854 10127 10906
rect 10127 10854 10157 10906
rect 10181 10854 10191 10906
rect 10191 10854 10237 10906
rect 9941 10852 9997 10854
rect 10021 10852 10077 10854
rect 10101 10852 10157 10854
rect 10181 10852 10237 10854
rect 9954 10668 10010 10704
rect 9954 10648 9956 10668
rect 9956 10648 10008 10668
rect 10008 10648 10010 10668
rect 10138 10376 10194 10432
rect 10138 10124 10194 10160
rect 10138 10104 10140 10124
rect 10140 10104 10192 10124
rect 10192 10104 10194 10124
rect 10598 12144 10654 12200
rect 9586 8900 9642 8936
rect 9586 8880 9588 8900
rect 9588 8880 9640 8900
rect 9640 8880 9642 8900
rect 9494 8372 9496 8392
rect 9496 8372 9548 8392
rect 9548 8372 9550 8392
rect 9494 8336 9550 8372
rect 10322 9832 10378 9888
rect 9941 9818 9997 9820
rect 10021 9818 10077 9820
rect 10101 9818 10157 9820
rect 10181 9818 10237 9820
rect 9941 9766 9987 9818
rect 9987 9766 9997 9818
rect 10021 9766 10051 9818
rect 10051 9766 10063 9818
rect 10063 9766 10077 9818
rect 10101 9766 10115 9818
rect 10115 9766 10127 9818
rect 10127 9766 10157 9818
rect 10181 9766 10191 9818
rect 10191 9766 10237 9818
rect 9941 9764 9997 9766
rect 10021 9764 10077 9766
rect 10101 9764 10157 9766
rect 10181 9764 10237 9766
rect 10322 9696 10378 9752
rect 9678 5636 9734 5672
rect 9678 5616 9680 5636
rect 9680 5616 9732 5636
rect 9732 5616 9734 5636
rect 10230 9444 10286 9480
rect 10230 9424 10232 9444
rect 10232 9424 10284 9444
rect 10284 9424 10286 9444
rect 9862 9288 9918 9344
rect 9941 8730 9997 8732
rect 10021 8730 10077 8732
rect 10101 8730 10157 8732
rect 10181 8730 10237 8732
rect 9941 8678 9987 8730
rect 9987 8678 9997 8730
rect 10021 8678 10051 8730
rect 10051 8678 10063 8730
rect 10063 8678 10077 8730
rect 10101 8678 10115 8730
rect 10115 8678 10127 8730
rect 10127 8678 10157 8730
rect 10181 8678 10191 8730
rect 10191 8678 10237 8730
rect 9941 8676 9997 8678
rect 10021 8676 10077 8678
rect 10101 8676 10157 8678
rect 10181 8676 10237 8678
rect 10138 8472 10194 8528
rect 10046 8336 10102 8392
rect 9941 7642 9997 7644
rect 10021 7642 10077 7644
rect 10101 7642 10157 7644
rect 10181 7642 10237 7644
rect 9941 7590 9987 7642
rect 9987 7590 9997 7642
rect 10021 7590 10051 7642
rect 10051 7590 10063 7642
rect 10063 7590 10077 7642
rect 10101 7590 10115 7642
rect 10115 7590 10127 7642
rect 10127 7590 10157 7642
rect 10181 7590 10191 7642
rect 10191 7590 10237 7642
rect 9941 7588 9997 7590
rect 10021 7588 10077 7590
rect 10101 7588 10157 7590
rect 10181 7588 10237 7590
rect 9941 6554 9997 6556
rect 10021 6554 10077 6556
rect 10101 6554 10157 6556
rect 10181 6554 10237 6556
rect 9941 6502 9987 6554
rect 9987 6502 9997 6554
rect 10021 6502 10051 6554
rect 10051 6502 10063 6554
rect 10063 6502 10077 6554
rect 10101 6502 10115 6554
rect 10115 6502 10127 6554
rect 10127 6502 10157 6554
rect 10181 6502 10191 6554
rect 10191 6502 10237 6554
rect 9941 6500 9997 6502
rect 10021 6500 10077 6502
rect 10101 6500 10157 6502
rect 10181 6500 10237 6502
rect 10230 6160 10286 6216
rect 9954 5616 10010 5672
rect 9941 5466 9997 5468
rect 10021 5466 10077 5468
rect 10101 5466 10157 5468
rect 10181 5466 10237 5468
rect 9941 5414 9987 5466
rect 9987 5414 9997 5466
rect 10021 5414 10051 5466
rect 10051 5414 10063 5466
rect 10063 5414 10077 5466
rect 10101 5414 10115 5466
rect 10115 5414 10127 5466
rect 10127 5414 10157 5466
rect 10181 5414 10191 5466
rect 10191 5414 10237 5466
rect 9941 5412 9997 5414
rect 10021 5412 10077 5414
rect 10101 5412 10157 5414
rect 10181 5412 10237 5414
rect 10230 5208 10286 5264
rect 9941 4378 9997 4380
rect 10021 4378 10077 4380
rect 10101 4378 10157 4380
rect 10181 4378 10237 4380
rect 9941 4326 9987 4378
rect 9987 4326 9997 4378
rect 10021 4326 10051 4378
rect 10051 4326 10063 4378
rect 10063 4326 10077 4378
rect 10101 4326 10115 4378
rect 10115 4326 10127 4378
rect 10127 4326 10157 4378
rect 10181 4326 10191 4378
rect 10191 4326 10237 4378
rect 9941 4324 9997 4326
rect 10021 4324 10077 4326
rect 10101 4324 10157 4326
rect 10181 4324 10237 4326
rect 11242 21936 11298 21992
rect 11242 18672 11298 18728
rect 11242 17992 11298 18048
rect 11334 17448 11390 17504
rect 11334 16224 11390 16280
rect 11610 18828 11666 18864
rect 11610 18808 11612 18828
rect 11612 18808 11664 18828
rect 11664 18808 11666 18828
rect 10874 12280 10930 12336
rect 10782 12144 10838 12200
rect 10690 10512 10746 10568
rect 9941 3290 9997 3292
rect 10021 3290 10077 3292
rect 10101 3290 10157 3292
rect 10181 3290 10237 3292
rect 9941 3238 9987 3290
rect 9987 3238 9997 3290
rect 10021 3238 10051 3290
rect 10051 3238 10063 3290
rect 10063 3238 10077 3290
rect 10101 3238 10115 3290
rect 10115 3238 10127 3290
rect 10127 3238 10157 3290
rect 10181 3238 10191 3290
rect 10191 3238 10237 3290
rect 9941 3236 9997 3238
rect 10021 3236 10077 3238
rect 10101 3236 10157 3238
rect 10181 3236 10237 3238
rect 9941 2202 9997 2204
rect 10021 2202 10077 2204
rect 10101 2202 10157 2204
rect 10181 2202 10237 2204
rect 9941 2150 9987 2202
rect 9987 2150 9997 2202
rect 10021 2150 10051 2202
rect 10051 2150 10063 2202
rect 10063 2150 10077 2202
rect 10101 2150 10115 2202
rect 10115 2150 10127 2202
rect 10127 2150 10157 2202
rect 10181 2150 10191 2202
rect 10191 2150 10237 2202
rect 9941 2148 9997 2150
rect 10021 2148 10077 2150
rect 10101 2148 10157 2150
rect 10181 2148 10237 2150
rect 10966 10784 11022 10840
rect 11058 8608 11114 8664
rect 11150 6840 11206 6896
rect 10782 5208 10838 5264
rect 11058 5072 11114 5128
rect 11058 2760 11114 2816
rect 10966 2488 11022 2544
rect 11334 14864 11390 14920
rect 11518 14184 11574 14240
rect 11518 13932 11574 13968
rect 11518 13912 11520 13932
rect 11520 13912 11572 13932
rect 11572 13912 11574 13932
rect 12162 27648 12218 27704
rect 13634 27376 13690 27432
rect 13266 26424 13322 26480
rect 12346 20304 12402 20360
rect 11978 17040 12034 17096
rect 11886 14592 11942 14648
rect 11426 10920 11482 10976
rect 11334 10648 11390 10704
rect 11702 10104 11758 10160
rect 11518 9424 11574 9480
rect 11794 9288 11850 9344
rect 11794 8880 11850 8936
rect 11610 8336 11666 8392
rect 12162 17196 12218 17232
rect 12162 17176 12164 17196
rect 12164 17176 12216 17196
rect 12216 17176 12218 17196
rect 12530 18944 12586 19000
rect 12622 17448 12678 17504
rect 12254 15816 12310 15872
rect 12162 14728 12218 14784
rect 12346 9968 12402 10024
rect 12346 9016 12402 9072
rect 12346 8372 12348 8392
rect 12348 8372 12400 8392
rect 12400 8372 12402 8392
rect 12346 8336 12402 8372
rect 11702 6724 11758 6760
rect 11702 6704 11704 6724
rect 11704 6704 11756 6724
rect 11756 6704 11758 6724
rect 12530 16088 12586 16144
rect 12622 15680 12678 15736
rect 13082 20984 13138 21040
rect 12806 20440 12862 20496
rect 12806 18400 12862 18456
rect 12990 19624 13046 19680
rect 12990 18536 13046 18592
rect 12714 15272 12770 15328
rect 12714 14456 12770 14512
rect 13082 18264 13138 18320
rect 14830 27920 14886 27976
rect 14434 27770 14490 27772
rect 14514 27770 14570 27772
rect 14594 27770 14650 27772
rect 14674 27770 14730 27772
rect 14434 27718 14480 27770
rect 14480 27718 14490 27770
rect 14514 27718 14544 27770
rect 14544 27718 14556 27770
rect 14556 27718 14570 27770
rect 14594 27718 14608 27770
rect 14608 27718 14620 27770
rect 14620 27718 14650 27770
rect 14674 27718 14684 27770
rect 14684 27718 14730 27770
rect 14434 27716 14490 27718
rect 14514 27716 14570 27718
rect 14594 27716 14650 27718
rect 14674 27716 14730 27718
rect 13910 27412 13912 27432
rect 13912 27412 13964 27432
rect 13964 27412 13966 27432
rect 13910 27376 13966 27412
rect 14434 26682 14490 26684
rect 14514 26682 14570 26684
rect 14594 26682 14650 26684
rect 14674 26682 14730 26684
rect 14434 26630 14480 26682
rect 14480 26630 14490 26682
rect 14514 26630 14544 26682
rect 14544 26630 14556 26682
rect 14556 26630 14570 26682
rect 14594 26630 14608 26682
rect 14608 26630 14620 26682
rect 14620 26630 14650 26682
rect 14674 26630 14684 26682
rect 14684 26630 14730 26682
rect 14434 26628 14490 26630
rect 14514 26628 14570 26630
rect 14594 26628 14650 26630
rect 14674 26628 14730 26630
rect 14554 26424 14610 26480
rect 13634 22344 13690 22400
rect 13450 19508 13506 19544
rect 13450 19488 13452 19508
rect 13452 19488 13504 19508
rect 13504 19488 13506 19508
rect 13266 18808 13322 18864
rect 13082 16360 13138 16416
rect 13082 15544 13138 15600
rect 13358 16088 13414 16144
rect 13174 13912 13230 13968
rect 13082 12416 13138 12472
rect 12530 10920 12586 10976
rect 12530 9036 12586 9072
rect 12530 9016 12532 9036
rect 12532 9016 12584 9036
rect 12584 9016 12586 9036
rect 13082 11192 13138 11248
rect 13082 10376 13138 10432
rect 13266 13368 13322 13424
rect 12990 6296 13046 6352
rect 12162 2760 12218 2816
rect 12622 3068 12624 3088
rect 12624 3068 12676 3088
rect 12676 3068 12678 3088
rect 12622 3032 12678 3068
rect 13174 8336 13230 8392
rect 13174 8200 13230 8256
rect 13542 14864 13598 14920
rect 13450 10920 13506 10976
rect 13542 9968 13598 10024
rect 14434 25594 14490 25596
rect 14514 25594 14570 25596
rect 14594 25594 14650 25596
rect 14674 25594 14730 25596
rect 14434 25542 14480 25594
rect 14480 25542 14490 25594
rect 14514 25542 14544 25594
rect 14544 25542 14556 25594
rect 14556 25542 14570 25594
rect 14594 25542 14608 25594
rect 14608 25542 14620 25594
rect 14620 25542 14650 25594
rect 14674 25542 14684 25594
rect 14684 25542 14730 25594
rect 14434 25540 14490 25542
rect 14514 25540 14570 25542
rect 14594 25540 14650 25542
rect 14674 25540 14730 25542
rect 14434 24506 14490 24508
rect 14514 24506 14570 24508
rect 14594 24506 14650 24508
rect 14674 24506 14730 24508
rect 14434 24454 14480 24506
rect 14480 24454 14490 24506
rect 14514 24454 14544 24506
rect 14544 24454 14556 24506
rect 14556 24454 14570 24506
rect 14594 24454 14608 24506
rect 14608 24454 14620 24506
rect 14620 24454 14650 24506
rect 14674 24454 14684 24506
rect 14684 24454 14730 24506
rect 14434 24452 14490 24454
rect 14514 24452 14570 24454
rect 14594 24452 14650 24454
rect 14674 24452 14730 24454
rect 14434 23418 14490 23420
rect 14514 23418 14570 23420
rect 14594 23418 14650 23420
rect 14674 23418 14730 23420
rect 14434 23366 14480 23418
rect 14480 23366 14490 23418
rect 14514 23366 14544 23418
rect 14544 23366 14556 23418
rect 14556 23366 14570 23418
rect 14594 23366 14608 23418
rect 14608 23366 14620 23418
rect 14620 23366 14650 23418
rect 14674 23366 14684 23418
rect 14684 23366 14730 23418
rect 14434 23364 14490 23366
rect 14514 23364 14570 23366
rect 14594 23364 14650 23366
rect 14674 23364 14730 23366
rect 14002 20984 14058 21040
rect 14434 22330 14490 22332
rect 14514 22330 14570 22332
rect 14594 22330 14650 22332
rect 14674 22330 14730 22332
rect 14434 22278 14480 22330
rect 14480 22278 14490 22330
rect 14514 22278 14544 22330
rect 14544 22278 14556 22330
rect 14556 22278 14570 22330
rect 14594 22278 14608 22330
rect 14608 22278 14620 22330
rect 14620 22278 14650 22330
rect 14674 22278 14684 22330
rect 14684 22278 14730 22330
rect 14434 22276 14490 22278
rect 14514 22276 14570 22278
rect 14594 22276 14650 22278
rect 14674 22276 14730 22278
rect 14434 21242 14490 21244
rect 14514 21242 14570 21244
rect 14594 21242 14650 21244
rect 14674 21242 14730 21244
rect 14434 21190 14480 21242
rect 14480 21190 14490 21242
rect 14514 21190 14544 21242
rect 14544 21190 14556 21242
rect 14556 21190 14570 21242
rect 14594 21190 14608 21242
rect 14608 21190 14620 21242
rect 14620 21190 14650 21242
rect 14674 21190 14684 21242
rect 14684 21190 14730 21242
rect 14434 21188 14490 21190
rect 14514 21188 14570 21190
rect 14594 21188 14650 21190
rect 14674 21188 14730 21190
rect 14186 20032 14242 20088
rect 14434 20154 14490 20156
rect 14514 20154 14570 20156
rect 14594 20154 14650 20156
rect 14674 20154 14730 20156
rect 14434 20102 14480 20154
rect 14480 20102 14490 20154
rect 14514 20102 14544 20154
rect 14544 20102 14556 20154
rect 14556 20102 14570 20154
rect 14594 20102 14608 20154
rect 14608 20102 14620 20154
rect 14620 20102 14650 20154
rect 14674 20102 14684 20154
rect 14684 20102 14730 20154
rect 14434 20100 14490 20102
rect 14514 20100 14570 20102
rect 14594 20100 14650 20102
rect 14674 20100 14730 20102
rect 14370 19916 14426 19952
rect 14370 19896 14372 19916
rect 14372 19896 14424 19916
rect 14424 19896 14426 19916
rect 14094 19760 14150 19816
rect 14186 19624 14242 19680
rect 13910 19488 13966 19544
rect 13910 19216 13966 19272
rect 13818 16108 13874 16144
rect 13818 16088 13820 16108
rect 13820 16088 13872 16108
rect 13872 16088 13874 16108
rect 14646 19660 14648 19680
rect 14648 19660 14700 19680
rect 14700 19660 14702 19680
rect 14646 19624 14702 19660
rect 14094 19116 14096 19136
rect 14096 19116 14148 19136
rect 14148 19116 14150 19136
rect 14094 19080 14150 19116
rect 14186 18944 14242 19000
rect 14830 19216 14886 19272
rect 14434 19066 14490 19068
rect 14514 19066 14570 19068
rect 14594 19066 14650 19068
rect 14674 19066 14730 19068
rect 14434 19014 14480 19066
rect 14480 19014 14490 19066
rect 14514 19014 14544 19066
rect 14544 19014 14556 19066
rect 14556 19014 14570 19066
rect 14594 19014 14608 19066
rect 14608 19014 14620 19066
rect 14620 19014 14650 19066
rect 14674 19014 14684 19066
rect 14684 19014 14730 19066
rect 14434 19012 14490 19014
rect 14514 19012 14570 19014
rect 14594 19012 14650 19014
rect 14674 19012 14730 19014
rect 14830 18672 14886 18728
rect 14094 17992 14150 18048
rect 13726 14320 13782 14376
rect 13726 12416 13782 12472
rect 14434 17978 14490 17980
rect 14514 17978 14570 17980
rect 14594 17978 14650 17980
rect 14674 17978 14730 17980
rect 14434 17926 14480 17978
rect 14480 17926 14490 17978
rect 14514 17926 14544 17978
rect 14544 17926 14556 17978
rect 14556 17926 14570 17978
rect 14594 17926 14608 17978
rect 14608 17926 14620 17978
rect 14620 17926 14650 17978
rect 14674 17926 14684 17978
rect 14684 17926 14730 17978
rect 14434 17924 14490 17926
rect 14514 17924 14570 17926
rect 14594 17924 14650 17926
rect 14674 17924 14730 17926
rect 14370 17196 14426 17232
rect 14370 17176 14372 17196
rect 14372 17176 14424 17196
rect 14424 17176 14426 17196
rect 14434 16890 14490 16892
rect 14514 16890 14570 16892
rect 14594 16890 14650 16892
rect 14674 16890 14730 16892
rect 14434 16838 14480 16890
rect 14480 16838 14490 16890
rect 14514 16838 14544 16890
rect 14544 16838 14556 16890
rect 14556 16838 14570 16890
rect 14594 16838 14608 16890
rect 14608 16838 14620 16890
rect 14620 16838 14650 16890
rect 14674 16838 14684 16890
rect 14684 16838 14730 16890
rect 14434 16836 14490 16838
rect 14514 16836 14570 16838
rect 14594 16836 14650 16838
rect 14674 16836 14730 16838
rect 14830 16360 14886 16416
rect 14370 15952 14426 16008
rect 14434 15802 14490 15804
rect 14514 15802 14570 15804
rect 14594 15802 14650 15804
rect 14674 15802 14730 15804
rect 14434 15750 14480 15802
rect 14480 15750 14490 15802
rect 14514 15750 14544 15802
rect 14544 15750 14556 15802
rect 14556 15750 14570 15802
rect 14594 15750 14608 15802
rect 14608 15750 14620 15802
rect 14620 15750 14650 15802
rect 14674 15750 14684 15802
rect 14684 15750 14730 15802
rect 14434 15748 14490 15750
rect 14514 15748 14570 15750
rect 14594 15748 14650 15750
rect 14674 15748 14730 15750
rect 14646 15544 14702 15600
rect 14002 12824 14058 12880
rect 13910 8608 13966 8664
rect 14554 15428 14610 15464
rect 14554 15408 14556 15428
rect 14556 15408 14608 15428
rect 14608 15408 14610 15428
rect 14434 14714 14490 14716
rect 14514 14714 14570 14716
rect 14594 14714 14650 14716
rect 14674 14714 14730 14716
rect 14434 14662 14480 14714
rect 14480 14662 14490 14714
rect 14514 14662 14544 14714
rect 14544 14662 14556 14714
rect 14556 14662 14570 14714
rect 14594 14662 14608 14714
rect 14608 14662 14620 14714
rect 14620 14662 14650 14714
rect 14674 14662 14684 14714
rect 14684 14662 14730 14714
rect 14434 14660 14490 14662
rect 14514 14660 14570 14662
rect 14594 14660 14650 14662
rect 14674 14660 14730 14662
rect 14646 14048 14702 14104
rect 14434 13626 14490 13628
rect 14514 13626 14570 13628
rect 14594 13626 14650 13628
rect 14674 13626 14730 13628
rect 14434 13574 14480 13626
rect 14480 13574 14490 13626
rect 14514 13574 14544 13626
rect 14544 13574 14556 13626
rect 14556 13574 14570 13626
rect 14594 13574 14608 13626
rect 14608 13574 14620 13626
rect 14620 13574 14650 13626
rect 14674 13574 14684 13626
rect 14684 13574 14730 13626
rect 14434 13572 14490 13574
rect 14514 13572 14570 13574
rect 14594 13572 14650 13574
rect 14674 13572 14730 13574
rect 15198 26288 15254 26344
rect 15014 21392 15070 21448
rect 15106 18128 15162 18184
rect 15106 15680 15162 15736
rect 15014 14184 15070 14240
rect 15014 13912 15070 13968
rect 14434 12538 14490 12540
rect 14514 12538 14570 12540
rect 14594 12538 14650 12540
rect 14674 12538 14730 12540
rect 14434 12486 14480 12538
rect 14480 12486 14490 12538
rect 14514 12486 14544 12538
rect 14544 12486 14556 12538
rect 14556 12486 14570 12538
rect 14594 12486 14608 12538
rect 14608 12486 14620 12538
rect 14620 12486 14650 12538
rect 14674 12486 14684 12538
rect 14684 12486 14730 12538
rect 14434 12484 14490 12486
rect 14514 12484 14570 12486
rect 14594 12484 14650 12486
rect 14674 12484 14730 12486
rect 14186 12008 14242 12064
rect 14646 11892 14702 11928
rect 14646 11872 14648 11892
rect 14648 11872 14700 11892
rect 14700 11872 14702 11892
rect 14434 11450 14490 11452
rect 14514 11450 14570 11452
rect 14594 11450 14650 11452
rect 14674 11450 14730 11452
rect 14434 11398 14480 11450
rect 14480 11398 14490 11450
rect 14514 11398 14544 11450
rect 14544 11398 14556 11450
rect 14556 11398 14570 11450
rect 14594 11398 14608 11450
rect 14608 11398 14620 11450
rect 14620 11398 14650 11450
rect 14674 11398 14684 11450
rect 14684 11398 14730 11450
rect 14434 11396 14490 11398
rect 14514 11396 14570 11398
rect 14594 11396 14650 11398
rect 14674 11396 14730 11398
rect 14094 10104 14150 10160
rect 14434 10362 14490 10364
rect 14514 10362 14570 10364
rect 14594 10362 14650 10364
rect 14674 10362 14730 10364
rect 14434 10310 14480 10362
rect 14480 10310 14490 10362
rect 14514 10310 14544 10362
rect 14544 10310 14556 10362
rect 14556 10310 14570 10362
rect 14594 10310 14608 10362
rect 14608 10310 14620 10362
rect 14620 10310 14650 10362
rect 14674 10310 14684 10362
rect 14684 10310 14730 10362
rect 14434 10308 14490 10310
rect 14514 10308 14570 10310
rect 14594 10308 14650 10310
rect 14674 10308 14730 10310
rect 14830 10104 14886 10160
rect 14186 9968 14242 10024
rect 14554 9832 14610 9888
rect 14094 8200 14150 8256
rect 14186 8064 14242 8120
rect 14434 9274 14490 9276
rect 14514 9274 14570 9276
rect 14594 9274 14650 9276
rect 14674 9274 14730 9276
rect 14434 9222 14480 9274
rect 14480 9222 14490 9274
rect 14514 9222 14544 9274
rect 14544 9222 14556 9274
rect 14556 9222 14570 9274
rect 14594 9222 14608 9274
rect 14608 9222 14620 9274
rect 14620 9222 14650 9274
rect 14674 9222 14684 9274
rect 14684 9222 14730 9274
rect 14434 9220 14490 9222
rect 14514 9220 14570 9222
rect 14594 9220 14650 9222
rect 14674 9220 14730 9222
rect 14434 8186 14490 8188
rect 14514 8186 14570 8188
rect 14594 8186 14650 8188
rect 14674 8186 14730 8188
rect 14434 8134 14480 8186
rect 14480 8134 14490 8186
rect 14514 8134 14544 8186
rect 14544 8134 14556 8186
rect 14556 8134 14570 8186
rect 14594 8134 14608 8186
rect 14608 8134 14620 8186
rect 14620 8134 14650 8186
rect 14674 8134 14684 8186
rect 14684 8134 14730 8186
rect 14434 8132 14490 8134
rect 14514 8132 14570 8134
rect 14594 8132 14650 8134
rect 14674 8132 14730 8134
rect 14370 7928 14426 7984
rect 14434 7098 14490 7100
rect 14514 7098 14570 7100
rect 14594 7098 14650 7100
rect 14674 7098 14730 7100
rect 14434 7046 14480 7098
rect 14480 7046 14490 7098
rect 14514 7046 14544 7098
rect 14544 7046 14556 7098
rect 14556 7046 14570 7098
rect 14594 7046 14608 7098
rect 14608 7046 14620 7098
rect 14620 7046 14650 7098
rect 14674 7046 14684 7098
rect 14684 7046 14730 7098
rect 14434 7044 14490 7046
rect 14514 7044 14570 7046
rect 14594 7044 14650 7046
rect 14674 7044 14730 7046
rect 15474 19292 15530 19348
rect 15658 21528 15714 21584
rect 15934 19896 15990 19952
rect 15474 16768 15530 16824
rect 15382 15272 15438 15328
rect 15474 14864 15530 14920
rect 15474 13912 15530 13968
rect 15198 11464 15254 11520
rect 14738 6196 14740 6216
rect 14740 6196 14792 6216
rect 14792 6196 14794 6216
rect 14738 6160 14794 6196
rect 14434 6010 14490 6012
rect 14514 6010 14570 6012
rect 14594 6010 14650 6012
rect 14674 6010 14730 6012
rect 14434 5958 14480 6010
rect 14480 5958 14490 6010
rect 14514 5958 14544 6010
rect 14544 5958 14556 6010
rect 14556 5958 14570 6010
rect 14594 5958 14608 6010
rect 14608 5958 14620 6010
rect 14620 5958 14650 6010
rect 14674 5958 14684 6010
rect 14684 5958 14730 6010
rect 14434 5956 14490 5958
rect 14514 5956 14570 5958
rect 14594 5956 14650 5958
rect 14674 5956 14730 5958
rect 14370 5752 14426 5808
rect 14434 4922 14490 4924
rect 14514 4922 14570 4924
rect 14594 4922 14650 4924
rect 14674 4922 14730 4924
rect 14434 4870 14480 4922
rect 14480 4870 14490 4922
rect 14514 4870 14544 4922
rect 14544 4870 14556 4922
rect 14556 4870 14570 4922
rect 14594 4870 14608 4922
rect 14608 4870 14620 4922
rect 14620 4870 14650 4922
rect 14674 4870 14684 4922
rect 14684 4870 14730 4922
rect 14434 4868 14490 4870
rect 14514 4868 14570 4870
rect 14594 4868 14650 4870
rect 14674 4868 14730 4870
rect 14434 3834 14490 3836
rect 14514 3834 14570 3836
rect 14594 3834 14650 3836
rect 14674 3834 14730 3836
rect 14434 3782 14480 3834
rect 14480 3782 14490 3834
rect 14514 3782 14544 3834
rect 14544 3782 14556 3834
rect 14556 3782 14570 3834
rect 14594 3782 14608 3834
rect 14608 3782 14620 3834
rect 14620 3782 14650 3834
rect 14674 3782 14684 3834
rect 14684 3782 14730 3834
rect 14434 3780 14490 3782
rect 14514 3780 14570 3782
rect 14594 3780 14650 3782
rect 14674 3780 14730 3782
rect 14434 2746 14490 2748
rect 14514 2746 14570 2748
rect 14594 2746 14650 2748
rect 14674 2746 14730 2748
rect 14434 2694 14480 2746
rect 14480 2694 14490 2746
rect 14514 2694 14544 2746
rect 14544 2694 14556 2746
rect 14556 2694 14570 2746
rect 14594 2694 14608 2746
rect 14608 2694 14620 2746
rect 14620 2694 14650 2746
rect 14674 2694 14684 2746
rect 14684 2694 14730 2746
rect 14434 2692 14490 2694
rect 14514 2692 14570 2694
rect 14594 2692 14650 2694
rect 14674 2692 14730 2694
rect 15106 5752 15162 5808
rect 15474 12960 15530 13016
rect 15858 19080 15914 19136
rect 15750 17992 15806 18048
rect 15658 16632 15714 16688
rect 15934 16516 15990 16552
rect 15934 16496 15936 16516
rect 15936 16496 15988 16516
rect 15988 16496 15990 16516
rect 15750 16360 15806 16416
rect 15658 15136 15714 15192
rect 16670 24792 16726 24848
rect 16210 18400 16266 18456
rect 15842 13776 15898 13832
rect 15842 12824 15898 12880
rect 15934 12280 15990 12336
rect 15934 11464 15990 11520
rect 16210 15136 16266 15192
rect 16026 10648 16082 10704
rect 15842 9016 15898 9072
rect 15842 8372 15844 8392
rect 15844 8372 15896 8392
rect 15896 8372 15898 8392
rect 15842 8336 15898 8372
rect 15566 6296 15622 6352
rect 15658 5616 15714 5672
rect 15934 6160 15990 6216
rect 16486 19252 16488 19272
rect 16488 19252 16540 19272
rect 16540 19252 16542 19272
rect 16486 19216 16542 19252
rect 16486 17720 16542 17776
rect 16486 17448 16542 17504
rect 16394 16768 16450 16824
rect 16762 17176 16818 17232
rect 16578 14612 16634 14648
rect 16578 14592 16580 14612
rect 16580 14592 16632 14612
rect 16632 14592 16634 14612
rect 16670 14456 16726 14512
rect 16670 10104 16726 10160
rect 16854 17040 16910 17096
rect 17038 18672 17094 18728
rect 16946 16904 17002 16960
rect 17222 18672 17278 18728
rect 17222 18128 17278 18184
rect 17130 17176 17186 17232
rect 18926 28314 18982 28316
rect 19006 28314 19062 28316
rect 19086 28314 19142 28316
rect 19166 28314 19222 28316
rect 18926 28262 18972 28314
rect 18972 28262 18982 28314
rect 19006 28262 19036 28314
rect 19036 28262 19048 28314
rect 19048 28262 19062 28314
rect 19086 28262 19100 28314
rect 19100 28262 19112 28314
rect 19112 28262 19142 28314
rect 19166 28262 19176 28314
rect 19176 28262 19222 28314
rect 18926 28260 18982 28262
rect 19006 28260 19062 28262
rect 19086 28260 19142 28262
rect 19166 28260 19222 28262
rect 18926 27226 18982 27228
rect 19006 27226 19062 27228
rect 19086 27226 19142 27228
rect 19166 27226 19222 27228
rect 18926 27174 18972 27226
rect 18972 27174 18982 27226
rect 19006 27174 19036 27226
rect 19036 27174 19048 27226
rect 19048 27174 19062 27226
rect 19086 27174 19100 27226
rect 19100 27174 19112 27226
rect 19112 27174 19142 27226
rect 19166 27174 19176 27226
rect 19176 27174 19222 27226
rect 18926 27172 18982 27174
rect 19006 27172 19062 27174
rect 19086 27172 19142 27174
rect 19166 27172 19222 27174
rect 19246 26288 19302 26344
rect 18926 26138 18982 26140
rect 19006 26138 19062 26140
rect 19086 26138 19142 26140
rect 19166 26138 19222 26140
rect 18926 26086 18972 26138
rect 18972 26086 18982 26138
rect 19006 26086 19036 26138
rect 19036 26086 19048 26138
rect 19048 26086 19062 26138
rect 19086 26086 19100 26138
rect 19100 26086 19112 26138
rect 19112 26086 19142 26138
rect 19166 26086 19176 26138
rect 19176 26086 19222 26138
rect 18926 26084 18982 26086
rect 19006 26084 19062 26086
rect 19086 26084 19142 26086
rect 19166 26084 19222 26086
rect 17406 17992 17462 18048
rect 17222 16088 17278 16144
rect 17130 15272 17186 15328
rect 17130 13368 17186 13424
rect 16946 12144 17002 12200
rect 16854 7656 16910 7712
rect 16762 7404 16818 7440
rect 16762 7384 16764 7404
rect 16764 7384 16816 7404
rect 16816 7384 16818 7404
rect 16670 6568 16726 6624
rect 16762 6160 16818 6216
rect 16946 7248 17002 7304
rect 17038 5480 17094 5536
rect 17314 11600 17370 11656
rect 17314 11056 17370 11112
rect 17774 20440 17830 20496
rect 17590 18128 17646 18184
rect 17866 17856 17922 17912
rect 17590 15000 17646 15056
rect 17590 13640 17646 13696
rect 17590 12280 17646 12336
rect 18234 21800 18290 21856
rect 18326 19896 18382 19952
rect 18234 18400 18290 18456
rect 19338 26152 19394 26208
rect 19522 26152 19578 26208
rect 19338 25880 19394 25936
rect 19522 25880 19578 25936
rect 18926 25050 18982 25052
rect 19006 25050 19062 25052
rect 19086 25050 19142 25052
rect 19166 25050 19222 25052
rect 18926 24998 18972 25050
rect 18972 24998 18982 25050
rect 19006 24998 19036 25050
rect 19036 24998 19048 25050
rect 19048 24998 19062 25050
rect 19086 24998 19100 25050
rect 19100 24998 19112 25050
rect 19112 24998 19142 25050
rect 19166 24998 19176 25050
rect 19176 24998 19222 25050
rect 18926 24996 18982 24998
rect 19006 24996 19062 24998
rect 19086 24996 19142 24998
rect 19166 24996 19222 24998
rect 18926 23962 18982 23964
rect 19006 23962 19062 23964
rect 19086 23962 19142 23964
rect 19166 23962 19222 23964
rect 18926 23910 18972 23962
rect 18972 23910 18982 23962
rect 19006 23910 19036 23962
rect 19036 23910 19048 23962
rect 19048 23910 19062 23962
rect 19086 23910 19100 23962
rect 19100 23910 19112 23962
rect 19112 23910 19142 23962
rect 19166 23910 19176 23962
rect 19176 23910 19222 23962
rect 18926 23908 18982 23910
rect 19006 23908 19062 23910
rect 19086 23908 19142 23910
rect 19166 23908 19222 23910
rect 19430 24792 19486 24848
rect 18926 22874 18982 22876
rect 19006 22874 19062 22876
rect 19086 22874 19142 22876
rect 19166 22874 19222 22876
rect 18926 22822 18972 22874
rect 18972 22822 18982 22874
rect 19006 22822 19036 22874
rect 19036 22822 19048 22874
rect 19048 22822 19062 22874
rect 19086 22822 19100 22874
rect 19100 22822 19112 22874
rect 19112 22822 19142 22874
rect 19166 22822 19176 22874
rect 19176 22822 19222 22874
rect 18926 22820 18982 22822
rect 19006 22820 19062 22822
rect 19086 22820 19142 22822
rect 19166 22820 19222 22822
rect 18926 21786 18982 21788
rect 19006 21786 19062 21788
rect 19086 21786 19142 21788
rect 19166 21786 19222 21788
rect 18926 21734 18972 21786
rect 18972 21734 18982 21786
rect 19006 21734 19036 21786
rect 19036 21734 19048 21786
rect 19048 21734 19062 21786
rect 19086 21734 19100 21786
rect 19100 21734 19112 21786
rect 19112 21734 19142 21786
rect 19166 21734 19176 21786
rect 19176 21734 19222 21786
rect 18926 21732 18982 21734
rect 19006 21732 19062 21734
rect 19086 21732 19142 21734
rect 19166 21732 19222 21734
rect 18142 17856 18198 17912
rect 18234 17040 18290 17096
rect 18050 13232 18106 13288
rect 17774 13096 17830 13152
rect 17958 12960 18014 13016
rect 17866 12824 17922 12880
rect 17590 12008 17646 12064
rect 17590 11872 17646 11928
rect 17682 11736 17738 11792
rect 17866 10784 17922 10840
rect 17774 9968 17830 10024
rect 17866 6704 17922 6760
rect 17866 6604 17868 6624
rect 17868 6604 17920 6624
rect 17920 6604 17922 6624
rect 17866 6568 17922 6604
rect 18510 18400 18566 18456
rect 18926 20698 18982 20700
rect 19006 20698 19062 20700
rect 19086 20698 19142 20700
rect 19166 20698 19222 20700
rect 18926 20646 18972 20698
rect 18972 20646 18982 20698
rect 19006 20646 19036 20698
rect 19036 20646 19048 20698
rect 19048 20646 19062 20698
rect 19086 20646 19100 20698
rect 19100 20646 19112 20698
rect 19112 20646 19142 20698
rect 19166 20646 19176 20698
rect 19176 20646 19222 20698
rect 18926 20644 18982 20646
rect 19006 20644 19062 20646
rect 19086 20644 19142 20646
rect 19166 20644 19222 20646
rect 19154 19796 19156 19816
rect 19156 19796 19208 19816
rect 19208 19796 19210 19816
rect 19154 19760 19210 19796
rect 18926 19610 18982 19612
rect 19006 19610 19062 19612
rect 19086 19610 19142 19612
rect 19166 19610 19222 19612
rect 18926 19558 18972 19610
rect 18972 19558 18982 19610
rect 19006 19558 19036 19610
rect 19036 19558 19048 19610
rect 19048 19558 19062 19610
rect 19086 19558 19100 19610
rect 19100 19558 19112 19610
rect 19112 19558 19142 19610
rect 19166 19558 19176 19610
rect 19176 19558 19222 19610
rect 18926 19556 18982 19558
rect 19006 19556 19062 19558
rect 19086 19556 19142 19558
rect 19166 19556 19222 19558
rect 18970 19352 19026 19408
rect 18602 18128 18658 18184
rect 18418 16904 18474 16960
rect 18786 19216 18842 19272
rect 18878 19080 18934 19136
rect 19522 24248 19578 24304
rect 19522 23724 19578 23760
rect 19522 23704 19524 23724
rect 19524 23704 19576 23724
rect 19576 23704 19578 23724
rect 19522 22888 19578 22944
rect 19522 22208 19578 22264
rect 20718 26288 20774 26344
rect 20626 26016 20682 26072
rect 19982 22208 20038 22264
rect 19798 21664 19854 21720
rect 19706 21528 19762 21584
rect 19890 21528 19946 21584
rect 18970 18944 19026 19000
rect 19062 18808 19118 18864
rect 18878 18672 18934 18728
rect 18926 18522 18982 18524
rect 19006 18522 19062 18524
rect 19086 18522 19142 18524
rect 19166 18522 19222 18524
rect 18926 18470 18972 18522
rect 18972 18470 18982 18522
rect 19006 18470 19036 18522
rect 19036 18470 19048 18522
rect 19048 18470 19062 18522
rect 19086 18470 19100 18522
rect 19100 18470 19112 18522
rect 19112 18470 19142 18522
rect 19166 18470 19176 18522
rect 19176 18470 19222 18522
rect 18926 18468 18982 18470
rect 19006 18468 19062 18470
rect 19086 18468 19142 18470
rect 19166 18468 19222 18470
rect 18878 18300 18880 18320
rect 18880 18300 18932 18320
rect 18932 18300 18934 18320
rect 18878 18264 18934 18300
rect 18970 17992 19026 18048
rect 19062 17756 19064 17776
rect 19064 17756 19116 17776
rect 19116 17756 19118 17776
rect 19062 17720 19118 17756
rect 18926 17434 18982 17436
rect 19006 17434 19062 17436
rect 19086 17434 19142 17436
rect 19166 17434 19222 17436
rect 18926 17382 18972 17434
rect 18972 17382 18982 17434
rect 19006 17382 19036 17434
rect 19036 17382 19048 17434
rect 19048 17382 19062 17434
rect 19086 17382 19100 17434
rect 19100 17382 19112 17434
rect 19112 17382 19142 17434
rect 19166 17382 19176 17434
rect 19176 17382 19222 17434
rect 18926 17380 18982 17382
rect 19006 17380 19062 17382
rect 19086 17380 19142 17382
rect 19166 17380 19222 17382
rect 18510 16768 18566 16824
rect 18510 16532 18512 16552
rect 18512 16532 18564 16552
rect 18564 16532 18566 16552
rect 18510 16496 18566 16532
rect 18510 14320 18566 14376
rect 18418 13932 18474 13968
rect 18418 13912 18420 13932
rect 18420 13912 18472 13932
rect 18472 13912 18474 13932
rect 18510 13132 18512 13152
rect 18512 13132 18564 13152
rect 18564 13132 18566 13152
rect 18326 12960 18382 13016
rect 18510 13096 18566 13132
rect 18510 12960 18566 13016
rect 18050 11056 18106 11112
rect 17866 6296 17922 6352
rect 17958 6024 18014 6080
rect 18234 6704 18290 6760
rect 18142 6296 18198 6352
rect 18970 16632 19026 16688
rect 18926 16346 18982 16348
rect 19006 16346 19062 16348
rect 19086 16346 19142 16348
rect 19166 16346 19222 16348
rect 18926 16294 18972 16346
rect 18972 16294 18982 16346
rect 19006 16294 19036 16346
rect 19036 16294 19048 16346
rect 19048 16294 19062 16346
rect 19086 16294 19100 16346
rect 19100 16294 19112 16346
rect 19112 16294 19142 16346
rect 19166 16294 19176 16346
rect 19176 16294 19222 16346
rect 18926 16292 18982 16294
rect 19006 16292 19062 16294
rect 19086 16292 19142 16294
rect 19166 16292 19222 16294
rect 18926 15258 18982 15260
rect 19006 15258 19062 15260
rect 19086 15258 19142 15260
rect 19166 15258 19222 15260
rect 18926 15206 18972 15258
rect 18972 15206 18982 15258
rect 19006 15206 19036 15258
rect 19036 15206 19048 15258
rect 19048 15206 19062 15258
rect 19086 15206 19100 15258
rect 19100 15206 19112 15258
rect 19112 15206 19142 15258
rect 19166 15206 19176 15258
rect 19176 15206 19222 15258
rect 18926 15204 18982 15206
rect 19006 15204 19062 15206
rect 19086 15204 19142 15206
rect 19166 15204 19222 15206
rect 19522 18264 19578 18320
rect 18926 14170 18982 14172
rect 19006 14170 19062 14172
rect 19086 14170 19142 14172
rect 19166 14170 19222 14172
rect 18926 14118 18972 14170
rect 18972 14118 18982 14170
rect 19006 14118 19036 14170
rect 19036 14118 19048 14170
rect 19048 14118 19062 14170
rect 19086 14118 19100 14170
rect 19100 14118 19112 14170
rect 19112 14118 19142 14170
rect 19166 14118 19176 14170
rect 19176 14118 19222 14170
rect 18926 14116 18982 14118
rect 19006 14116 19062 14118
rect 19086 14116 19142 14118
rect 19166 14116 19222 14118
rect 19154 13912 19210 13968
rect 19154 13504 19210 13560
rect 18694 12960 18750 13016
rect 18926 13082 18982 13084
rect 19006 13082 19062 13084
rect 19086 13082 19142 13084
rect 19166 13082 19222 13084
rect 18926 13030 18972 13082
rect 18972 13030 18982 13082
rect 19006 13030 19036 13082
rect 19036 13030 19048 13082
rect 19048 13030 19062 13082
rect 19086 13030 19100 13082
rect 19100 13030 19112 13082
rect 19112 13030 19142 13082
rect 19166 13030 19176 13082
rect 19176 13030 19222 13082
rect 18926 13028 18982 13030
rect 19006 13028 19062 13030
rect 19086 13028 19142 13030
rect 19166 13028 19222 13030
rect 18970 12144 19026 12200
rect 19522 13948 19524 13968
rect 19524 13948 19576 13968
rect 19576 13948 19578 13968
rect 19522 13912 19578 13948
rect 19522 13096 19578 13152
rect 18926 11994 18982 11996
rect 19006 11994 19062 11996
rect 19086 11994 19142 11996
rect 19166 11994 19222 11996
rect 18926 11942 18972 11994
rect 18972 11942 18982 11994
rect 19006 11942 19036 11994
rect 19036 11942 19048 11994
rect 19048 11942 19062 11994
rect 19086 11942 19100 11994
rect 19100 11942 19112 11994
rect 19112 11942 19142 11994
rect 19166 11942 19176 11994
rect 19176 11942 19222 11994
rect 18926 11940 18982 11942
rect 19006 11940 19062 11942
rect 19086 11940 19142 11942
rect 19166 11940 19222 11942
rect 18878 11756 18934 11792
rect 18878 11736 18880 11756
rect 18880 11736 18932 11756
rect 18932 11736 18934 11756
rect 18926 10906 18982 10908
rect 19006 10906 19062 10908
rect 19086 10906 19142 10908
rect 19166 10906 19222 10908
rect 18926 10854 18972 10906
rect 18972 10854 18982 10906
rect 19006 10854 19036 10906
rect 19036 10854 19048 10906
rect 19048 10854 19062 10906
rect 19086 10854 19100 10906
rect 19100 10854 19112 10906
rect 19112 10854 19142 10906
rect 19166 10854 19176 10906
rect 19176 10854 19222 10906
rect 18926 10852 18982 10854
rect 19006 10852 19062 10854
rect 19086 10852 19142 10854
rect 19166 10852 19222 10854
rect 19246 10648 19302 10704
rect 18926 9818 18982 9820
rect 19006 9818 19062 9820
rect 19086 9818 19142 9820
rect 19166 9818 19222 9820
rect 18926 9766 18972 9818
rect 18972 9766 18982 9818
rect 19006 9766 19036 9818
rect 19036 9766 19048 9818
rect 19048 9766 19062 9818
rect 19086 9766 19100 9818
rect 19100 9766 19112 9818
rect 19112 9766 19142 9818
rect 19166 9766 19176 9818
rect 19176 9766 19222 9818
rect 18926 9764 18982 9766
rect 19006 9764 19062 9766
rect 19086 9764 19142 9766
rect 19166 9764 19222 9766
rect 19430 10512 19486 10568
rect 19338 10104 19394 10160
rect 19430 9988 19486 10024
rect 19430 9968 19432 9988
rect 19432 9968 19484 9988
rect 19484 9968 19486 9988
rect 18694 8880 18750 8936
rect 19246 9016 19302 9072
rect 18926 8730 18982 8732
rect 19006 8730 19062 8732
rect 19086 8730 19142 8732
rect 19166 8730 19222 8732
rect 18926 8678 18972 8730
rect 18972 8678 18982 8730
rect 19006 8678 19036 8730
rect 19036 8678 19048 8730
rect 19048 8678 19062 8730
rect 19086 8678 19100 8730
rect 19100 8678 19112 8730
rect 19112 8678 19142 8730
rect 19166 8678 19176 8730
rect 19176 8678 19222 8730
rect 18926 8676 18982 8678
rect 19006 8676 19062 8678
rect 19086 8676 19142 8678
rect 19166 8676 19222 8678
rect 19430 8200 19486 8256
rect 18926 7642 18982 7644
rect 19006 7642 19062 7644
rect 19086 7642 19142 7644
rect 19166 7642 19222 7644
rect 18926 7590 18972 7642
rect 18972 7590 18982 7642
rect 19006 7590 19036 7642
rect 19036 7590 19048 7642
rect 19048 7590 19062 7642
rect 19086 7590 19100 7642
rect 19100 7590 19112 7642
rect 19112 7590 19142 7642
rect 19166 7590 19176 7642
rect 19176 7590 19222 7642
rect 18926 7588 18982 7590
rect 19006 7588 19062 7590
rect 19086 7588 19142 7590
rect 19166 7588 19222 7590
rect 18926 6554 18982 6556
rect 19006 6554 19062 6556
rect 19086 6554 19142 6556
rect 19166 6554 19222 6556
rect 18926 6502 18972 6554
rect 18972 6502 18982 6554
rect 19006 6502 19036 6554
rect 19036 6502 19048 6554
rect 19048 6502 19062 6554
rect 19086 6502 19100 6554
rect 19100 6502 19112 6554
rect 19112 6502 19142 6554
rect 19166 6502 19176 6554
rect 19176 6502 19222 6554
rect 18926 6500 18982 6502
rect 19006 6500 19062 6502
rect 19086 6500 19142 6502
rect 19166 6500 19222 6502
rect 18926 5466 18982 5468
rect 19006 5466 19062 5468
rect 19086 5466 19142 5468
rect 19166 5466 19222 5468
rect 18926 5414 18972 5466
rect 18972 5414 18982 5466
rect 19006 5414 19036 5466
rect 19036 5414 19048 5466
rect 19048 5414 19062 5466
rect 19086 5414 19100 5466
rect 19100 5414 19112 5466
rect 19112 5414 19142 5466
rect 19166 5414 19176 5466
rect 19176 5414 19222 5466
rect 18926 5412 18982 5414
rect 19006 5412 19062 5414
rect 19086 5412 19142 5414
rect 19166 5412 19222 5414
rect 18926 4378 18982 4380
rect 19006 4378 19062 4380
rect 19086 4378 19142 4380
rect 19166 4378 19222 4380
rect 18926 4326 18972 4378
rect 18972 4326 18982 4378
rect 19006 4326 19036 4378
rect 19036 4326 19048 4378
rect 19048 4326 19062 4378
rect 19086 4326 19100 4378
rect 19100 4326 19112 4378
rect 19112 4326 19142 4378
rect 19166 4326 19176 4378
rect 19176 4326 19222 4378
rect 18926 4324 18982 4326
rect 19006 4324 19062 4326
rect 19086 4324 19142 4326
rect 19166 4324 19222 4326
rect 19706 12300 19762 12336
rect 19706 12280 19708 12300
rect 19708 12280 19760 12300
rect 19760 12280 19762 12300
rect 20074 19216 20130 19272
rect 19890 15000 19946 15056
rect 19890 14612 19946 14648
rect 19890 14592 19892 14612
rect 19892 14592 19944 14612
rect 19944 14592 19946 14612
rect 19890 13776 19946 13832
rect 19890 11192 19946 11248
rect 20626 24792 20682 24848
rect 20350 19216 20406 19272
rect 19338 3984 19394 4040
rect 19430 3848 19486 3904
rect 18926 3290 18982 3292
rect 19006 3290 19062 3292
rect 19086 3290 19142 3292
rect 19166 3290 19222 3292
rect 18926 3238 18972 3290
rect 18972 3238 18982 3290
rect 19006 3238 19036 3290
rect 19036 3238 19048 3290
rect 19048 3238 19062 3290
rect 19086 3238 19100 3290
rect 19100 3238 19112 3290
rect 19112 3238 19142 3290
rect 19166 3238 19176 3290
rect 19176 3238 19222 3290
rect 18926 3236 18982 3238
rect 19006 3236 19062 3238
rect 19086 3236 19142 3238
rect 19166 3236 19222 3238
rect 18786 3168 18842 3224
rect 18926 2202 18982 2204
rect 19006 2202 19062 2204
rect 19086 2202 19142 2204
rect 19166 2202 19222 2204
rect 18926 2150 18972 2202
rect 18972 2150 18982 2202
rect 19006 2150 19036 2202
rect 19036 2150 19048 2202
rect 19048 2150 19062 2202
rect 19086 2150 19100 2202
rect 19100 2150 19112 2202
rect 19112 2150 19142 2202
rect 19166 2150 19176 2202
rect 19176 2150 19222 2202
rect 18926 2148 18982 2150
rect 19006 2148 19062 2150
rect 19086 2148 19142 2150
rect 19166 2148 19222 2150
rect 20718 23024 20774 23080
rect 20626 21528 20682 21584
rect 21270 24792 21326 24848
rect 21270 24248 21326 24304
rect 21178 23704 21234 23760
rect 21086 23432 21142 23488
rect 21178 23196 21180 23216
rect 21180 23196 21232 23216
rect 21232 23196 21234 23216
rect 21178 23160 21234 23196
rect 21086 22888 21142 22944
rect 21270 22888 21326 22944
rect 21454 23976 21510 24032
rect 21822 25900 21878 25936
rect 21822 25880 21824 25900
rect 21824 25880 21876 25900
rect 21876 25880 21878 25900
rect 21638 23568 21694 23624
rect 21546 23296 21602 23352
rect 20718 17176 20774 17232
rect 21178 19080 21234 19136
rect 21086 17176 21142 17232
rect 21178 16904 21234 16960
rect 20534 14456 20590 14512
rect 20718 15136 20774 15192
rect 20534 13368 20590 13424
rect 20626 13096 20682 13152
rect 20442 9696 20498 9752
rect 20442 8744 20498 8800
rect 20350 7384 20406 7440
rect 20718 10804 20774 10840
rect 20718 10784 20720 10804
rect 20720 10784 20772 10804
rect 20772 10784 20774 10804
rect 19982 5208 20038 5264
rect 20074 2916 20130 2952
rect 20074 2896 20076 2916
rect 20076 2896 20128 2916
rect 20128 2896 20130 2916
rect 20258 5480 20314 5536
rect 20350 5072 20406 5128
rect 21086 15544 21142 15600
rect 20994 12960 21050 13016
rect 20902 10956 20904 10976
rect 20904 10956 20956 10976
rect 20956 10956 20958 10976
rect 20902 10920 20958 10956
rect 21546 17584 21602 17640
rect 21546 17176 21602 17232
rect 21546 14476 21602 14512
rect 21546 14456 21548 14476
rect 21548 14456 21600 14476
rect 21600 14456 21602 14476
rect 21454 14184 21510 14240
rect 21454 13912 21510 13968
rect 21270 12552 21326 12608
rect 21270 12416 21326 12472
rect 21178 11872 21234 11928
rect 21546 13640 21602 13696
rect 22098 23976 22154 24032
rect 22006 23316 22062 23352
rect 22006 23296 22008 23316
rect 22008 23296 22060 23316
rect 22060 23296 22062 23316
rect 22374 23568 22430 23624
rect 22282 23432 22338 23488
rect 22190 22208 22246 22264
rect 21822 20712 21878 20768
rect 22282 20712 22338 20768
rect 22006 19352 22062 19408
rect 22190 19488 22246 19544
rect 22374 19508 22430 19544
rect 22374 19488 22376 19508
rect 22376 19488 22428 19508
rect 22428 19488 22430 19508
rect 21822 17040 21878 17096
rect 22098 18264 22154 18320
rect 22006 16632 22062 16688
rect 22190 15308 22192 15328
rect 22192 15308 22244 15328
rect 22244 15308 22246 15328
rect 22190 15272 22246 15308
rect 22190 15020 22246 15056
rect 22190 15000 22192 15020
rect 22192 15000 22244 15020
rect 22244 15000 22246 15020
rect 22098 14320 22154 14376
rect 21730 13912 21786 13968
rect 22006 13912 22062 13968
rect 21178 10512 21234 10568
rect 20810 7384 20866 7440
rect 20626 5364 20682 5400
rect 20626 5344 20628 5364
rect 20628 5344 20680 5364
rect 20680 5344 20682 5364
rect 20626 5072 20682 5128
rect 20994 6296 21050 6352
rect 20994 5908 21050 5944
rect 20994 5888 20996 5908
rect 20996 5888 21048 5908
rect 21048 5888 21050 5908
rect 20994 2896 21050 2952
rect 21362 6432 21418 6488
rect 21362 5752 21418 5808
rect 21730 12008 21786 12064
rect 21638 9052 21640 9072
rect 21640 9052 21692 9072
rect 21692 9052 21694 9072
rect 21638 9016 21694 9052
rect 21546 7248 21602 7304
rect 21730 7656 21786 7712
rect 21730 7248 21786 7304
rect 22190 14184 22246 14240
rect 22282 13776 22338 13832
rect 22098 13232 22154 13288
rect 22006 11600 22062 11656
rect 21914 10104 21970 10160
rect 22006 7928 22062 7984
rect 21822 5636 21878 5672
rect 21822 5616 21824 5636
rect 21824 5616 21876 5636
rect 21876 5616 21878 5636
rect 21914 5364 21970 5400
rect 21914 5344 21916 5364
rect 21916 5344 21968 5364
rect 21968 5344 21970 5364
rect 22834 23316 22890 23352
rect 22834 23296 22836 23316
rect 22836 23296 22888 23316
rect 22888 23296 22890 23316
rect 22650 19488 22706 19544
rect 22650 19372 22706 19408
rect 22650 19352 22652 19372
rect 22652 19352 22704 19372
rect 22704 19352 22706 19372
rect 22374 9560 22430 9616
rect 22282 6024 22338 6080
rect 22282 5208 22338 5264
rect 22650 14592 22706 14648
rect 22650 14320 22706 14376
rect 22650 13776 22706 13832
rect 22834 19352 22890 19408
rect 23419 27770 23475 27772
rect 23499 27770 23555 27772
rect 23579 27770 23635 27772
rect 23659 27770 23715 27772
rect 23419 27718 23465 27770
rect 23465 27718 23475 27770
rect 23499 27718 23529 27770
rect 23529 27718 23541 27770
rect 23541 27718 23555 27770
rect 23579 27718 23593 27770
rect 23593 27718 23605 27770
rect 23605 27718 23635 27770
rect 23659 27718 23669 27770
rect 23669 27718 23715 27770
rect 23419 27716 23475 27718
rect 23499 27716 23555 27718
rect 23579 27716 23635 27718
rect 23659 27716 23715 27718
rect 23846 27648 23902 27704
rect 23419 26682 23475 26684
rect 23499 26682 23555 26684
rect 23579 26682 23635 26684
rect 23659 26682 23715 26684
rect 23419 26630 23465 26682
rect 23465 26630 23475 26682
rect 23499 26630 23529 26682
rect 23529 26630 23541 26682
rect 23541 26630 23555 26682
rect 23579 26630 23593 26682
rect 23593 26630 23605 26682
rect 23605 26630 23635 26682
rect 23659 26630 23669 26682
rect 23669 26630 23715 26682
rect 23419 26628 23475 26630
rect 23499 26628 23555 26630
rect 23579 26628 23635 26630
rect 23659 26628 23715 26630
rect 23202 26288 23258 26344
rect 23202 25900 23258 25936
rect 23202 25880 23204 25900
rect 23204 25880 23256 25900
rect 23256 25880 23258 25900
rect 23419 25594 23475 25596
rect 23499 25594 23555 25596
rect 23579 25594 23635 25596
rect 23659 25594 23715 25596
rect 23419 25542 23465 25594
rect 23465 25542 23475 25594
rect 23499 25542 23529 25594
rect 23529 25542 23541 25594
rect 23541 25542 23555 25594
rect 23579 25542 23593 25594
rect 23593 25542 23605 25594
rect 23605 25542 23635 25594
rect 23659 25542 23669 25594
rect 23669 25542 23715 25594
rect 23419 25540 23475 25542
rect 23499 25540 23555 25542
rect 23579 25540 23635 25542
rect 23659 25540 23715 25542
rect 23419 24506 23475 24508
rect 23499 24506 23555 24508
rect 23579 24506 23635 24508
rect 23659 24506 23715 24508
rect 23419 24454 23465 24506
rect 23465 24454 23475 24506
rect 23499 24454 23529 24506
rect 23529 24454 23541 24506
rect 23541 24454 23555 24506
rect 23579 24454 23593 24506
rect 23593 24454 23605 24506
rect 23605 24454 23635 24506
rect 23659 24454 23669 24506
rect 23669 24454 23715 24506
rect 23419 24452 23475 24454
rect 23499 24452 23555 24454
rect 23579 24452 23635 24454
rect 23659 24452 23715 24454
rect 23419 23418 23475 23420
rect 23499 23418 23555 23420
rect 23579 23418 23635 23420
rect 23659 23418 23715 23420
rect 23419 23366 23465 23418
rect 23465 23366 23475 23418
rect 23499 23366 23529 23418
rect 23529 23366 23541 23418
rect 23541 23366 23555 23418
rect 23579 23366 23593 23418
rect 23593 23366 23605 23418
rect 23605 23366 23635 23418
rect 23659 23366 23669 23418
rect 23669 23366 23715 23418
rect 23419 23364 23475 23366
rect 23499 23364 23555 23366
rect 23579 23364 23635 23366
rect 23659 23364 23715 23366
rect 23386 23160 23442 23216
rect 23419 22330 23475 22332
rect 23499 22330 23555 22332
rect 23579 22330 23635 22332
rect 23659 22330 23715 22332
rect 23419 22278 23465 22330
rect 23465 22278 23475 22330
rect 23499 22278 23529 22330
rect 23529 22278 23541 22330
rect 23541 22278 23555 22330
rect 23579 22278 23593 22330
rect 23593 22278 23605 22330
rect 23605 22278 23635 22330
rect 23659 22278 23669 22330
rect 23669 22278 23715 22330
rect 23419 22276 23475 22278
rect 23499 22276 23555 22278
rect 23579 22276 23635 22278
rect 23659 22276 23715 22278
rect 23419 21242 23475 21244
rect 23499 21242 23555 21244
rect 23579 21242 23635 21244
rect 23659 21242 23715 21244
rect 23419 21190 23465 21242
rect 23465 21190 23475 21242
rect 23499 21190 23529 21242
rect 23529 21190 23541 21242
rect 23541 21190 23555 21242
rect 23579 21190 23593 21242
rect 23593 21190 23605 21242
rect 23605 21190 23635 21242
rect 23659 21190 23669 21242
rect 23669 21190 23715 21242
rect 23419 21188 23475 21190
rect 23499 21188 23555 21190
rect 23579 21188 23635 21190
rect 23659 21188 23715 21190
rect 23846 26016 23902 26072
rect 23419 20154 23475 20156
rect 23499 20154 23555 20156
rect 23579 20154 23635 20156
rect 23659 20154 23715 20156
rect 23419 20102 23465 20154
rect 23465 20102 23475 20154
rect 23499 20102 23529 20154
rect 23529 20102 23541 20154
rect 23541 20102 23555 20154
rect 23579 20102 23593 20154
rect 23593 20102 23605 20154
rect 23605 20102 23635 20154
rect 23659 20102 23669 20154
rect 23669 20102 23715 20154
rect 23419 20100 23475 20102
rect 23499 20100 23555 20102
rect 23579 20100 23635 20102
rect 23659 20100 23715 20102
rect 23662 19252 23664 19272
rect 23664 19252 23716 19272
rect 23716 19252 23718 19272
rect 23662 19216 23718 19252
rect 23202 19080 23258 19136
rect 23419 19066 23475 19068
rect 23499 19066 23555 19068
rect 23579 19066 23635 19068
rect 23659 19066 23715 19068
rect 23419 19014 23465 19066
rect 23465 19014 23475 19066
rect 23499 19014 23529 19066
rect 23529 19014 23541 19066
rect 23541 19014 23555 19066
rect 23579 19014 23593 19066
rect 23593 19014 23605 19066
rect 23605 19014 23635 19066
rect 23659 19014 23669 19066
rect 23669 19014 23715 19066
rect 23419 19012 23475 19014
rect 23499 19012 23555 19014
rect 23579 19012 23635 19014
rect 23659 19012 23715 19014
rect 23419 17978 23475 17980
rect 23499 17978 23555 17980
rect 23579 17978 23635 17980
rect 23659 17978 23715 17980
rect 23419 17926 23465 17978
rect 23465 17926 23475 17978
rect 23499 17926 23529 17978
rect 23529 17926 23541 17978
rect 23541 17926 23555 17978
rect 23579 17926 23593 17978
rect 23593 17926 23605 17978
rect 23605 17926 23635 17978
rect 23659 17926 23669 17978
rect 23669 17926 23715 17978
rect 23419 17924 23475 17926
rect 23499 17924 23555 17926
rect 23579 17924 23635 17926
rect 23659 17924 23715 17926
rect 23018 17448 23074 17504
rect 23018 16904 23074 16960
rect 24398 22888 24454 22944
rect 23294 17040 23350 17096
rect 23018 16360 23074 16416
rect 23419 16890 23475 16892
rect 23499 16890 23555 16892
rect 23579 16890 23635 16892
rect 23659 16890 23715 16892
rect 23419 16838 23465 16890
rect 23465 16838 23475 16890
rect 23499 16838 23529 16890
rect 23529 16838 23541 16890
rect 23541 16838 23555 16890
rect 23579 16838 23593 16890
rect 23593 16838 23605 16890
rect 23605 16838 23635 16890
rect 23659 16838 23669 16890
rect 23669 16838 23715 16890
rect 23419 16836 23475 16838
rect 23499 16836 23555 16838
rect 23579 16836 23635 16838
rect 23659 16836 23715 16838
rect 23419 15802 23475 15804
rect 23499 15802 23555 15804
rect 23579 15802 23635 15804
rect 23659 15802 23715 15804
rect 23419 15750 23465 15802
rect 23465 15750 23475 15802
rect 23499 15750 23529 15802
rect 23529 15750 23541 15802
rect 23541 15750 23555 15802
rect 23579 15750 23593 15802
rect 23593 15750 23605 15802
rect 23605 15750 23635 15802
rect 23659 15750 23669 15802
rect 23669 15750 23715 15802
rect 23419 15748 23475 15750
rect 23499 15748 23555 15750
rect 23579 15748 23635 15750
rect 23659 15748 23715 15750
rect 23202 15408 23258 15464
rect 23110 15136 23166 15192
rect 23662 15136 23718 15192
rect 23202 14592 23258 14648
rect 23478 14884 23534 14920
rect 23478 14864 23480 14884
rect 23480 14864 23532 14884
rect 23532 14864 23534 14884
rect 23419 14714 23475 14716
rect 23499 14714 23555 14716
rect 23579 14714 23635 14716
rect 23659 14714 23715 14716
rect 23419 14662 23465 14714
rect 23465 14662 23475 14714
rect 23499 14662 23529 14714
rect 23529 14662 23541 14714
rect 23541 14662 23555 14714
rect 23579 14662 23593 14714
rect 23593 14662 23605 14714
rect 23605 14662 23635 14714
rect 23659 14662 23669 14714
rect 23669 14662 23715 14714
rect 23419 14660 23475 14662
rect 23499 14660 23555 14662
rect 23579 14660 23635 14662
rect 23659 14660 23715 14662
rect 23662 14456 23718 14512
rect 24490 19488 24546 19544
rect 24214 17720 24270 17776
rect 23110 14320 23166 14376
rect 23478 13912 23534 13968
rect 22650 6316 22706 6352
rect 22650 6296 22652 6316
rect 22652 6296 22704 6316
rect 22704 6296 22706 6316
rect 22466 5908 22522 5944
rect 22466 5888 22468 5908
rect 22468 5888 22520 5908
rect 22520 5888 22522 5908
rect 22558 4664 22614 4720
rect 23419 13626 23475 13628
rect 23499 13626 23555 13628
rect 23579 13626 23635 13628
rect 23659 13626 23715 13628
rect 23419 13574 23465 13626
rect 23465 13574 23475 13626
rect 23499 13574 23529 13626
rect 23529 13574 23541 13626
rect 23541 13574 23555 13626
rect 23579 13574 23593 13626
rect 23593 13574 23605 13626
rect 23605 13574 23635 13626
rect 23659 13574 23669 13626
rect 23669 13574 23715 13626
rect 23419 13572 23475 13574
rect 23499 13572 23555 13574
rect 23579 13572 23635 13574
rect 23659 13572 23715 13574
rect 23386 13096 23442 13152
rect 23419 12538 23475 12540
rect 23499 12538 23555 12540
rect 23579 12538 23635 12540
rect 23659 12538 23715 12540
rect 23419 12486 23465 12538
rect 23465 12486 23475 12538
rect 23499 12486 23529 12538
rect 23529 12486 23541 12538
rect 23541 12486 23555 12538
rect 23579 12486 23593 12538
rect 23593 12486 23605 12538
rect 23605 12486 23635 12538
rect 23659 12486 23669 12538
rect 23669 12486 23715 12538
rect 23419 12484 23475 12486
rect 23499 12484 23555 12486
rect 23579 12484 23635 12486
rect 23659 12484 23715 12486
rect 24030 13232 24086 13288
rect 24214 13948 24216 13968
rect 24216 13948 24268 13968
rect 24268 13948 24270 13968
rect 24214 13912 24270 13948
rect 24122 12688 24178 12744
rect 24122 12416 24178 12472
rect 23754 11600 23810 11656
rect 23419 11450 23475 11452
rect 23499 11450 23555 11452
rect 23579 11450 23635 11452
rect 23659 11450 23715 11452
rect 23419 11398 23465 11450
rect 23465 11398 23475 11450
rect 23499 11398 23529 11450
rect 23529 11398 23541 11450
rect 23541 11398 23555 11450
rect 23579 11398 23593 11450
rect 23593 11398 23605 11450
rect 23605 11398 23635 11450
rect 23659 11398 23669 11450
rect 23669 11398 23715 11450
rect 23419 11396 23475 11398
rect 23499 11396 23555 11398
rect 23579 11396 23635 11398
rect 23659 11396 23715 11398
rect 23419 10362 23475 10364
rect 23499 10362 23555 10364
rect 23579 10362 23635 10364
rect 23659 10362 23715 10364
rect 23419 10310 23465 10362
rect 23465 10310 23475 10362
rect 23499 10310 23529 10362
rect 23529 10310 23541 10362
rect 23541 10310 23555 10362
rect 23579 10310 23593 10362
rect 23593 10310 23605 10362
rect 23605 10310 23635 10362
rect 23659 10310 23669 10362
rect 23669 10310 23715 10362
rect 23419 10308 23475 10310
rect 23499 10308 23555 10310
rect 23579 10308 23635 10310
rect 23659 10308 23715 10310
rect 23294 9560 23350 9616
rect 23754 9424 23810 9480
rect 23419 9274 23475 9276
rect 23499 9274 23555 9276
rect 23579 9274 23635 9276
rect 23659 9274 23715 9276
rect 23419 9222 23465 9274
rect 23465 9222 23475 9274
rect 23499 9222 23529 9274
rect 23529 9222 23541 9274
rect 23541 9222 23555 9274
rect 23579 9222 23593 9274
rect 23593 9222 23605 9274
rect 23605 9222 23635 9274
rect 23659 9222 23669 9274
rect 23669 9222 23715 9274
rect 23419 9220 23475 9222
rect 23499 9220 23555 9222
rect 23579 9220 23635 9222
rect 23659 9220 23715 9222
rect 23662 8628 23718 8664
rect 23662 8608 23664 8628
rect 23664 8608 23716 8628
rect 23716 8608 23718 8628
rect 23386 8336 23442 8392
rect 23419 8186 23475 8188
rect 23499 8186 23555 8188
rect 23579 8186 23635 8188
rect 23659 8186 23715 8188
rect 23419 8134 23465 8186
rect 23465 8134 23475 8186
rect 23499 8134 23529 8186
rect 23529 8134 23541 8186
rect 23541 8134 23555 8186
rect 23579 8134 23593 8186
rect 23593 8134 23605 8186
rect 23605 8134 23635 8186
rect 23659 8134 23669 8186
rect 23669 8134 23715 8186
rect 23419 8132 23475 8134
rect 23499 8132 23555 8134
rect 23579 8132 23635 8134
rect 23659 8132 23715 8134
rect 23662 7928 23718 7984
rect 23110 5752 23166 5808
rect 23419 7098 23475 7100
rect 23499 7098 23555 7100
rect 23579 7098 23635 7100
rect 23659 7098 23715 7100
rect 23419 7046 23465 7098
rect 23465 7046 23475 7098
rect 23499 7046 23529 7098
rect 23529 7046 23541 7098
rect 23541 7046 23555 7098
rect 23579 7046 23593 7098
rect 23593 7046 23605 7098
rect 23605 7046 23635 7098
rect 23659 7046 23669 7098
rect 23669 7046 23715 7098
rect 23419 7044 23475 7046
rect 23499 7044 23555 7046
rect 23579 7044 23635 7046
rect 23659 7044 23715 7046
rect 23294 6432 23350 6488
rect 23419 6010 23475 6012
rect 23499 6010 23555 6012
rect 23579 6010 23635 6012
rect 23659 6010 23715 6012
rect 23419 5958 23465 6010
rect 23465 5958 23475 6010
rect 23499 5958 23529 6010
rect 23529 5958 23541 6010
rect 23541 5958 23555 6010
rect 23579 5958 23593 6010
rect 23593 5958 23605 6010
rect 23605 5958 23635 6010
rect 23659 5958 23669 6010
rect 23669 5958 23715 6010
rect 23419 5956 23475 5958
rect 23499 5956 23555 5958
rect 23579 5956 23635 5958
rect 23659 5956 23715 5958
rect 23478 5480 23534 5536
rect 23419 4922 23475 4924
rect 23499 4922 23555 4924
rect 23579 4922 23635 4924
rect 23659 4922 23715 4924
rect 23419 4870 23465 4922
rect 23465 4870 23475 4922
rect 23499 4870 23529 4922
rect 23529 4870 23541 4922
rect 23541 4870 23555 4922
rect 23579 4870 23593 4922
rect 23593 4870 23605 4922
rect 23605 4870 23635 4922
rect 23659 4870 23669 4922
rect 23669 4870 23715 4922
rect 23419 4868 23475 4870
rect 23499 4868 23555 4870
rect 23579 4868 23635 4870
rect 23659 4868 23715 4870
rect 23386 4664 23442 4720
rect 23419 3834 23475 3836
rect 23499 3834 23555 3836
rect 23579 3834 23635 3836
rect 23659 3834 23715 3836
rect 23419 3782 23465 3834
rect 23465 3782 23475 3834
rect 23499 3782 23529 3834
rect 23529 3782 23541 3834
rect 23541 3782 23555 3834
rect 23579 3782 23593 3834
rect 23593 3782 23605 3834
rect 23605 3782 23635 3834
rect 23659 3782 23669 3834
rect 23669 3782 23715 3834
rect 23419 3780 23475 3782
rect 23499 3780 23555 3782
rect 23579 3780 23635 3782
rect 23659 3780 23715 3782
rect 23419 2746 23475 2748
rect 23499 2746 23555 2748
rect 23579 2746 23635 2748
rect 23659 2746 23715 2748
rect 23419 2694 23465 2746
rect 23465 2694 23475 2746
rect 23499 2694 23529 2746
rect 23529 2694 23541 2746
rect 23541 2694 23555 2746
rect 23579 2694 23593 2746
rect 23593 2694 23605 2746
rect 23605 2694 23635 2746
rect 23659 2694 23669 2746
rect 23669 2694 23715 2746
rect 23419 2692 23475 2694
rect 23499 2692 23555 2694
rect 23579 2692 23635 2694
rect 23659 2692 23715 2694
rect 24122 8744 24178 8800
rect 24490 10104 24546 10160
rect 24306 7112 24362 7168
rect 24398 6840 24454 6896
rect 24398 6568 24454 6624
rect 24674 19488 24730 19544
rect 25594 23704 25650 23760
rect 25134 15000 25190 15056
rect 25318 14320 25374 14376
rect 25226 13776 25282 13832
rect 25870 21664 25926 21720
rect 26422 24928 26478 24984
rect 26146 21664 26202 21720
rect 25962 19624 26018 19680
rect 25778 19488 25834 19544
rect 24950 7404 25006 7440
rect 24950 7384 24952 7404
rect 24952 7384 25004 7404
rect 25004 7384 25006 7404
rect 24674 7112 24730 7168
rect 24582 6976 24638 7032
rect 24766 6704 24822 6760
rect 24214 5072 24270 5128
rect 25042 6704 25098 6760
rect 24674 5072 24730 5128
rect 25042 6432 25098 6488
rect 25318 8628 25374 8664
rect 25318 8608 25320 8628
rect 25320 8608 25372 8628
rect 25372 8608 25374 8628
rect 25318 8336 25374 8392
rect 25502 7248 25558 7304
rect 25410 5480 25466 5536
rect 26238 19216 26294 19272
rect 25870 12280 25926 12336
rect 25870 9696 25926 9752
rect 26790 25064 26846 25120
rect 27250 27276 27252 27296
rect 27252 27276 27304 27296
rect 27304 27276 27306 27296
rect 27250 27240 27306 27276
rect 27158 25336 27214 25392
rect 26790 17584 26846 17640
rect 26606 16768 26662 16824
rect 26514 14456 26570 14512
rect 26422 13368 26478 13424
rect 26146 12688 26202 12744
rect 25686 5344 25742 5400
rect 25962 7656 26018 7712
rect 26238 7928 26294 7984
rect 26054 6296 26110 6352
rect 26238 3848 26294 3904
rect 26606 12824 26662 12880
rect 26790 15544 26846 15600
rect 27250 19488 27306 19544
rect 27066 12688 27122 12744
rect 27526 12416 27582 12472
rect 27250 11620 27306 11656
rect 27250 11600 27252 11620
rect 27252 11600 27304 11620
rect 27304 11600 27306 11620
rect 27342 7520 27398 7576
rect 27526 7248 27582 7304
rect 27342 6452 27398 6488
rect 27342 6432 27344 6452
rect 27344 6432 27396 6452
rect 27396 6432 27398 6452
<< metal3 >>
rect 5436 28864 5756 28865
rect 5436 28800 5444 28864
rect 5508 28800 5524 28864
rect 5588 28800 5604 28864
rect 5668 28800 5684 28864
rect 5748 28800 5756 28864
rect 5436 28799 5756 28800
rect 14422 28864 14742 28865
rect 14422 28800 14430 28864
rect 14494 28800 14510 28864
rect 14574 28800 14590 28864
rect 14654 28800 14670 28864
rect 14734 28800 14742 28864
rect 14422 28799 14742 28800
rect 23407 28864 23727 28865
rect 23407 28800 23415 28864
rect 23479 28800 23495 28864
rect 23559 28800 23575 28864
rect 23639 28800 23655 28864
rect 23719 28800 23727 28864
rect 23407 28799 23727 28800
rect 9929 28320 10249 28321
rect 9929 28256 9937 28320
rect 10001 28256 10017 28320
rect 10081 28256 10097 28320
rect 10161 28256 10177 28320
rect 10241 28256 10249 28320
rect 9929 28255 10249 28256
rect 18914 28320 19234 28321
rect 18914 28256 18922 28320
rect 18986 28256 19002 28320
rect 19066 28256 19082 28320
rect 19146 28256 19162 28320
rect 19226 28256 19234 28320
rect 18914 28255 19234 28256
rect 14222 27916 14228 27980
rect 14292 27978 14298 27980
rect 14825 27978 14891 27981
rect 14292 27976 14891 27978
rect 14292 27920 14830 27976
rect 14886 27920 14891 27976
rect 14292 27918 14891 27920
rect 14292 27916 14298 27918
rect 14825 27915 14891 27918
rect 5436 27776 5756 27777
rect 5436 27712 5444 27776
rect 5508 27712 5524 27776
rect 5588 27712 5604 27776
rect 5668 27712 5684 27776
rect 5748 27712 5756 27776
rect 5436 27711 5756 27712
rect 14422 27776 14742 27777
rect 14422 27712 14430 27776
rect 14494 27712 14510 27776
rect 14574 27712 14590 27776
rect 14654 27712 14670 27776
rect 14734 27712 14742 27776
rect 14422 27711 14742 27712
rect 23407 27776 23727 27777
rect 23407 27712 23415 27776
rect 23479 27712 23495 27776
rect 23559 27712 23575 27776
rect 23639 27712 23655 27776
rect 23719 27712 23727 27776
rect 23407 27711 23727 27712
rect 12157 27708 12223 27709
rect 23841 27708 23907 27709
rect 12157 27704 12204 27708
rect 12268 27706 12274 27708
rect 12157 27648 12162 27704
rect 12157 27644 12204 27648
rect 12268 27646 12314 27706
rect 12268 27644 12274 27646
rect 23790 27644 23796 27708
rect 23860 27706 23907 27708
rect 23860 27704 23952 27706
rect 23902 27648 23952 27704
rect 23860 27646 23952 27648
rect 23860 27644 23907 27646
rect 12157 27643 12223 27644
rect 23841 27643 23907 27644
rect 6177 27570 6243 27573
rect 7465 27570 7531 27573
rect 6177 27568 7531 27570
rect 6177 27512 6182 27568
rect 6238 27512 7470 27568
rect 7526 27512 7531 27568
rect 6177 27510 7531 27512
rect 6177 27507 6243 27510
rect 7465 27507 7531 27510
rect 8661 27434 8727 27437
rect 13629 27434 13695 27437
rect 13905 27434 13971 27437
rect 8661 27432 13971 27434
rect 8661 27376 8666 27432
rect 8722 27376 13634 27432
rect 13690 27376 13910 27432
rect 13966 27376 13971 27432
rect 8661 27374 13971 27376
rect 8661 27371 8727 27374
rect 13629 27371 13695 27374
rect 13905 27371 13971 27374
rect 27245 27298 27311 27301
rect 28373 27298 29173 27328
rect 27245 27296 29173 27298
rect 27245 27240 27250 27296
rect 27306 27240 29173 27296
rect 27245 27238 29173 27240
rect 27245 27235 27311 27238
rect 9929 27232 10249 27233
rect 9929 27168 9937 27232
rect 10001 27168 10017 27232
rect 10081 27168 10097 27232
rect 10161 27168 10177 27232
rect 10241 27168 10249 27232
rect 9929 27167 10249 27168
rect 18914 27232 19234 27233
rect 18914 27168 18922 27232
rect 18986 27168 19002 27232
rect 19066 27168 19082 27232
rect 19146 27168 19162 27232
rect 19226 27168 19234 27232
rect 28373 27208 29173 27238
rect 18914 27167 19234 27168
rect 6085 27026 6151 27029
rect 7189 27026 7255 27029
rect 6085 27024 7255 27026
rect 6085 26968 6090 27024
rect 6146 26968 7194 27024
rect 7250 26968 7255 27024
rect 6085 26966 7255 26968
rect 6085 26963 6151 26966
rect 7189 26963 7255 26966
rect 5441 26890 5507 26893
rect 6494 26890 6500 26892
rect 5441 26888 6500 26890
rect 5441 26832 5446 26888
rect 5502 26832 6500 26888
rect 5441 26830 6500 26832
rect 5441 26827 5507 26830
rect 6494 26828 6500 26830
rect 6564 26828 6570 26892
rect 5436 26688 5756 26689
rect 5436 26624 5444 26688
rect 5508 26624 5524 26688
rect 5588 26624 5604 26688
rect 5668 26624 5684 26688
rect 5748 26624 5756 26688
rect 5436 26623 5756 26624
rect 14422 26688 14742 26689
rect 14422 26624 14430 26688
rect 14494 26624 14510 26688
rect 14574 26624 14590 26688
rect 14654 26624 14670 26688
rect 14734 26624 14742 26688
rect 14422 26623 14742 26624
rect 23407 26688 23727 26689
rect 23407 26624 23415 26688
rect 23479 26624 23495 26688
rect 23559 26624 23575 26688
rect 23639 26624 23655 26688
rect 23719 26624 23727 26688
rect 23407 26623 23727 26624
rect 10869 26482 10935 26485
rect 11462 26482 11468 26484
rect 10869 26480 11468 26482
rect 10869 26424 10874 26480
rect 10930 26424 11468 26480
rect 10869 26422 11468 26424
rect 10869 26419 10935 26422
rect 11462 26420 11468 26422
rect 11532 26420 11538 26484
rect 13261 26482 13327 26485
rect 14549 26482 14615 26485
rect 13261 26480 14615 26482
rect 13261 26424 13266 26480
rect 13322 26424 14554 26480
rect 14610 26424 14615 26480
rect 13261 26422 14615 26424
rect 13261 26419 13327 26422
rect 14549 26419 14615 26422
rect 3049 26346 3115 26349
rect 3366 26346 3372 26348
rect 3049 26344 3372 26346
rect 3049 26288 3054 26344
rect 3110 26288 3372 26344
rect 3049 26286 3372 26288
rect 3049 26283 3115 26286
rect 3366 26284 3372 26286
rect 3436 26284 3442 26348
rect 15193 26346 15259 26349
rect 15326 26346 15332 26348
rect 15193 26344 15332 26346
rect 15193 26288 15198 26344
rect 15254 26288 15332 26344
rect 15193 26286 15332 26288
rect 15193 26283 15259 26286
rect 15326 26284 15332 26286
rect 15396 26284 15402 26348
rect 18270 26284 18276 26348
rect 18340 26346 18346 26348
rect 19241 26346 19307 26349
rect 18340 26344 19307 26346
rect 18340 26288 19246 26344
rect 19302 26288 19307 26344
rect 18340 26286 19307 26288
rect 18340 26284 18346 26286
rect 19241 26283 19307 26286
rect 19558 26284 19564 26348
rect 19628 26346 19634 26348
rect 20713 26346 20779 26349
rect 19628 26344 20779 26346
rect 19628 26288 20718 26344
rect 20774 26288 20779 26344
rect 19628 26286 20779 26288
rect 19628 26284 19634 26286
rect 20713 26283 20779 26286
rect 23197 26348 23263 26349
rect 23197 26344 23244 26348
rect 23308 26346 23314 26348
rect 23197 26288 23202 26344
rect 23197 26284 23244 26288
rect 23308 26286 23354 26346
rect 23308 26284 23314 26286
rect 23197 26283 23263 26284
rect 19333 26208 19399 26213
rect 19333 26152 19338 26208
rect 19394 26152 19399 26208
rect 19333 26147 19399 26152
rect 19517 26210 19583 26213
rect 19517 26208 19626 26210
rect 19517 26152 19522 26208
rect 19578 26152 19626 26208
rect 19517 26147 19626 26152
rect 9929 26144 10249 26145
rect 9929 26080 9937 26144
rect 10001 26080 10017 26144
rect 10081 26080 10097 26144
rect 10161 26080 10177 26144
rect 10241 26080 10249 26144
rect 9929 26079 10249 26080
rect 18914 26144 19234 26145
rect 18914 26080 18922 26144
rect 18986 26080 19002 26144
rect 19066 26080 19082 26144
rect 19146 26080 19162 26144
rect 19226 26080 19234 26144
rect 18914 26079 19234 26080
rect 5257 26074 5323 26077
rect 6361 26074 6427 26077
rect 5257 26072 6427 26074
rect 5257 26016 5262 26072
rect 5318 26016 6366 26072
rect 6422 26016 6427 26072
rect 5257 26014 6427 26016
rect 5257 26011 5323 26014
rect 6361 26011 6427 26014
rect 19336 25941 19396 26147
rect 19566 25941 19626 26147
rect 20621 26074 20687 26077
rect 23841 26074 23907 26077
rect 20621 26072 23907 26074
rect 20621 26016 20626 26072
rect 20682 26016 23846 26072
rect 23902 26016 23907 26072
rect 20621 26014 23907 26016
rect 20621 26011 20687 26014
rect 23841 26011 23907 26014
rect 4429 25938 4495 25941
rect 5625 25938 5691 25941
rect 4429 25936 5691 25938
rect 4429 25880 4434 25936
rect 4490 25880 5630 25936
rect 5686 25880 5691 25936
rect 4429 25878 5691 25880
rect 4429 25875 4495 25878
rect 5625 25875 5691 25878
rect 19333 25936 19399 25941
rect 19333 25880 19338 25936
rect 19394 25880 19399 25936
rect 19333 25875 19399 25880
rect 19517 25936 19626 25941
rect 19517 25880 19522 25936
rect 19578 25880 19626 25936
rect 19517 25878 19626 25880
rect 21817 25938 21883 25941
rect 23197 25938 23263 25941
rect 21817 25936 23263 25938
rect 21817 25880 21822 25936
rect 21878 25880 23202 25936
rect 23258 25880 23263 25936
rect 21817 25878 23263 25880
rect 19517 25875 19583 25878
rect 21817 25875 21883 25878
rect 23197 25875 23263 25878
rect 5436 25600 5756 25601
rect 5436 25536 5444 25600
rect 5508 25536 5524 25600
rect 5588 25536 5604 25600
rect 5668 25536 5684 25600
rect 5748 25536 5756 25600
rect 5436 25535 5756 25536
rect 14422 25600 14742 25601
rect 14422 25536 14430 25600
rect 14494 25536 14510 25600
rect 14574 25536 14590 25600
rect 14654 25536 14670 25600
rect 14734 25536 14742 25600
rect 14422 25535 14742 25536
rect 23407 25600 23727 25601
rect 23407 25536 23415 25600
rect 23479 25536 23495 25600
rect 23559 25536 23575 25600
rect 23639 25536 23655 25600
rect 23719 25536 23727 25600
rect 23407 25535 23727 25536
rect 4521 25530 4587 25533
rect 5073 25530 5139 25533
rect 4521 25528 5139 25530
rect 4521 25472 4526 25528
rect 4582 25472 5078 25528
rect 5134 25472 5139 25528
rect 4521 25470 5139 25472
rect 4521 25467 4587 25470
rect 5073 25467 5139 25470
rect 5901 25530 5967 25533
rect 6453 25530 6519 25533
rect 5901 25528 6519 25530
rect 5901 25472 5906 25528
rect 5962 25472 6458 25528
rect 6514 25472 6519 25528
rect 5901 25470 6519 25472
rect 5901 25467 5967 25470
rect 6453 25467 6519 25470
rect 27153 25394 27219 25397
rect 27470 25394 27476 25396
rect 27153 25392 27476 25394
rect 27153 25336 27158 25392
rect 27214 25336 27476 25392
rect 27153 25334 27476 25336
rect 27153 25331 27219 25334
rect 27470 25332 27476 25334
rect 27540 25332 27546 25396
rect 25078 25060 25084 25124
rect 25148 25122 25154 25124
rect 26785 25122 26851 25125
rect 25148 25120 26851 25122
rect 25148 25064 26790 25120
rect 26846 25064 26851 25120
rect 25148 25062 26851 25064
rect 25148 25060 25154 25062
rect 26785 25059 26851 25062
rect 9929 25056 10249 25057
rect 9929 24992 9937 25056
rect 10001 24992 10017 25056
rect 10081 24992 10097 25056
rect 10161 24992 10177 25056
rect 10241 24992 10249 25056
rect 9929 24991 10249 24992
rect 18914 25056 19234 25057
rect 18914 24992 18922 25056
rect 18986 24992 19002 25056
rect 19066 24992 19082 25056
rect 19146 24992 19162 25056
rect 19226 24992 19234 25056
rect 18914 24991 19234 24992
rect 25262 24924 25268 24988
rect 25332 24986 25338 24988
rect 26417 24986 26483 24989
rect 25332 24984 26483 24986
rect 25332 24928 26422 24984
rect 26478 24928 26483 24984
rect 25332 24926 26483 24928
rect 25332 24924 25338 24926
rect 26417 24923 26483 24926
rect 15694 24788 15700 24852
rect 15764 24850 15770 24852
rect 16665 24850 16731 24853
rect 15764 24848 16731 24850
rect 15764 24792 16670 24848
rect 16726 24792 16731 24848
rect 15764 24790 16731 24792
rect 15764 24788 15770 24790
rect 16665 24787 16731 24790
rect 19425 24850 19491 24853
rect 20621 24850 20687 24853
rect 21265 24850 21331 24853
rect 19425 24848 21331 24850
rect 19425 24792 19430 24848
rect 19486 24792 20626 24848
rect 20682 24792 21270 24848
rect 21326 24792 21331 24848
rect 19425 24790 21331 24792
rect 19425 24787 19491 24790
rect 20621 24787 20687 24790
rect 21265 24787 21331 24790
rect 5533 24714 5599 24717
rect 6913 24714 6979 24717
rect 5533 24712 6979 24714
rect 5533 24656 5538 24712
rect 5594 24656 6918 24712
rect 6974 24656 6979 24712
rect 5533 24654 6979 24656
rect 5533 24651 5599 24654
rect 6913 24651 6979 24654
rect 6177 24578 6243 24581
rect 6913 24578 6979 24581
rect 6177 24576 6979 24578
rect 6177 24520 6182 24576
rect 6238 24520 6918 24576
rect 6974 24520 6979 24576
rect 6177 24518 6979 24520
rect 6177 24515 6243 24518
rect 6913 24515 6979 24518
rect 5436 24512 5756 24513
rect 5436 24448 5444 24512
rect 5508 24448 5524 24512
rect 5588 24448 5604 24512
rect 5668 24448 5684 24512
rect 5748 24448 5756 24512
rect 5436 24447 5756 24448
rect 14422 24512 14742 24513
rect 14422 24448 14430 24512
rect 14494 24448 14510 24512
rect 14574 24448 14590 24512
rect 14654 24448 14670 24512
rect 14734 24448 14742 24512
rect 14422 24447 14742 24448
rect 23407 24512 23727 24513
rect 23407 24448 23415 24512
rect 23479 24448 23495 24512
rect 23559 24448 23575 24512
rect 23639 24448 23655 24512
rect 23719 24448 23727 24512
rect 23407 24447 23727 24448
rect 19517 24306 19583 24309
rect 21265 24306 21331 24309
rect 19517 24304 21331 24306
rect 19517 24248 19522 24304
rect 19578 24248 21270 24304
rect 21326 24248 21331 24304
rect 19517 24246 21331 24248
rect 19517 24243 19583 24246
rect 21265 24243 21331 24246
rect 21449 24034 21515 24037
rect 22093 24034 22159 24037
rect 22686 24034 22692 24036
rect 21449 24032 22692 24034
rect 21449 23976 21454 24032
rect 21510 23976 22098 24032
rect 22154 23976 22692 24032
rect 21449 23974 22692 23976
rect 21449 23971 21515 23974
rect 22093 23971 22159 23974
rect 22686 23972 22692 23974
rect 22756 23972 22762 24036
rect 9929 23968 10249 23969
rect 9929 23904 9937 23968
rect 10001 23904 10017 23968
rect 10081 23904 10097 23968
rect 10161 23904 10177 23968
rect 10241 23904 10249 23968
rect 9929 23903 10249 23904
rect 18914 23968 19234 23969
rect 18914 23904 18922 23968
rect 18986 23904 19002 23968
rect 19066 23904 19082 23968
rect 19146 23904 19162 23968
rect 19226 23904 19234 23968
rect 18914 23903 19234 23904
rect 5165 23896 5231 23901
rect 5165 23840 5170 23896
rect 5226 23840 5231 23896
rect 5165 23835 5231 23840
rect 4245 23762 4311 23765
rect 5168 23762 5228 23835
rect 4245 23760 5228 23762
rect 4245 23704 4250 23760
rect 4306 23704 5228 23760
rect 4245 23702 5228 23704
rect 19517 23762 19583 23765
rect 21173 23762 21239 23765
rect 19517 23760 21239 23762
rect 19517 23704 19522 23760
rect 19578 23704 21178 23760
rect 21234 23704 21239 23760
rect 19517 23702 21239 23704
rect 4245 23699 4311 23702
rect 19517 23699 19583 23702
rect 21173 23699 21239 23702
rect 23974 23700 23980 23764
rect 24044 23762 24050 23764
rect 25589 23762 25655 23765
rect 24044 23760 25655 23762
rect 24044 23704 25594 23760
rect 25650 23704 25655 23760
rect 24044 23702 25655 23704
rect 24044 23700 24050 23702
rect 25589 23699 25655 23702
rect 21633 23626 21699 23629
rect 22369 23626 22435 23629
rect 21633 23624 22435 23626
rect 21633 23568 21638 23624
rect 21694 23568 22374 23624
rect 22430 23568 22435 23624
rect 21633 23566 22435 23568
rect 21633 23563 21699 23566
rect 22369 23563 22435 23566
rect 21081 23490 21147 23493
rect 22277 23492 22343 23493
rect 21214 23490 21220 23492
rect 21081 23488 21220 23490
rect 21081 23432 21086 23488
rect 21142 23432 21220 23488
rect 21081 23430 21220 23432
rect 21081 23427 21147 23430
rect 21214 23428 21220 23430
rect 21284 23428 21290 23492
rect 22277 23488 22324 23492
rect 22388 23490 22394 23492
rect 22277 23432 22282 23488
rect 22277 23428 22324 23432
rect 22388 23430 22434 23490
rect 22388 23428 22394 23430
rect 22277 23427 22343 23428
rect 5436 23424 5756 23425
rect 5436 23360 5444 23424
rect 5508 23360 5524 23424
rect 5588 23360 5604 23424
rect 5668 23360 5684 23424
rect 5748 23360 5756 23424
rect 5436 23359 5756 23360
rect 14422 23424 14742 23425
rect 14422 23360 14430 23424
rect 14494 23360 14510 23424
rect 14574 23360 14590 23424
rect 14654 23360 14670 23424
rect 14734 23360 14742 23424
rect 14422 23359 14742 23360
rect 23407 23424 23727 23425
rect 23407 23360 23415 23424
rect 23479 23360 23495 23424
rect 23559 23360 23575 23424
rect 23639 23360 23655 23424
rect 23719 23360 23727 23424
rect 23407 23359 23727 23360
rect 21541 23354 21607 23357
rect 20348 23352 21607 23354
rect 20348 23296 21546 23352
rect 21602 23296 21607 23352
rect 20348 23294 21607 23296
rect 2681 23082 2747 23085
rect 5809 23082 5875 23085
rect 2681 23080 5875 23082
rect 2681 23024 2686 23080
rect 2742 23024 5814 23080
rect 5870 23024 5875 23080
rect 2681 23022 5875 23024
rect 2681 23019 2747 23022
rect 5809 23019 5875 23022
rect 4337 22946 4403 22949
rect 4470 22946 4476 22948
rect 4337 22944 4476 22946
rect 4337 22888 4342 22944
rect 4398 22888 4476 22944
rect 4337 22886 4476 22888
rect 4337 22883 4403 22886
rect 4470 22884 4476 22886
rect 4540 22884 4546 22948
rect 19517 22946 19583 22949
rect 20348 22946 20408 23294
rect 21541 23291 21607 23294
rect 22001 23354 22067 23357
rect 22829 23354 22895 23357
rect 22001 23352 22895 23354
rect 22001 23296 22006 23352
rect 22062 23296 22834 23352
rect 22890 23296 22895 23352
rect 22001 23294 22895 23296
rect 22001 23291 22067 23294
rect 22829 23291 22895 23294
rect 21173 23218 21239 23221
rect 23238 23218 23244 23220
rect 21038 23216 21239 23218
rect 21038 23160 21178 23216
rect 21234 23160 21239 23216
rect 21038 23158 21239 23160
rect 20478 23020 20484 23084
rect 20548 23082 20554 23084
rect 20713 23082 20779 23085
rect 20548 23080 20779 23082
rect 20548 23024 20718 23080
rect 20774 23024 20779 23080
rect 20548 23022 20779 23024
rect 20548 23020 20554 23022
rect 20713 23019 20779 23022
rect 19517 22944 20408 22946
rect 19517 22888 19522 22944
rect 19578 22888 20408 22944
rect 19517 22886 20408 22888
rect 21038 22949 21098 23158
rect 21173 23155 21239 23158
rect 22050 23158 23244 23218
rect 21038 22944 21147 22949
rect 21038 22888 21086 22944
rect 21142 22888 21147 22944
rect 21038 22886 21147 22888
rect 19517 22883 19583 22886
rect 21081 22883 21147 22886
rect 21265 22946 21331 22949
rect 22050 22946 22110 23158
rect 23238 23156 23244 23158
rect 23308 23218 23314 23220
rect 23381 23218 23447 23221
rect 23308 23216 23447 23218
rect 23308 23160 23386 23216
rect 23442 23160 23447 23216
rect 23308 23158 23447 23160
rect 23308 23156 23314 23158
rect 23381 23155 23447 23158
rect 21265 22944 22110 22946
rect 21265 22888 21270 22944
rect 21326 22888 22110 22944
rect 21265 22886 22110 22888
rect 21265 22883 21331 22886
rect 9929 22880 10249 22881
rect 9929 22816 9937 22880
rect 10001 22816 10017 22880
rect 10081 22816 10097 22880
rect 10161 22816 10177 22880
rect 10241 22816 10249 22880
rect 9929 22815 10249 22816
rect 18914 22880 19234 22881
rect 18914 22816 18922 22880
rect 18986 22816 19002 22880
rect 19066 22816 19082 22880
rect 19146 22816 19162 22880
rect 19226 22816 19234 22880
rect 18914 22815 19234 22816
rect 3601 22810 3667 22813
rect 4245 22810 4311 22813
rect 5441 22810 5507 22813
rect 3601 22808 5507 22810
rect 3601 22752 3606 22808
rect 3662 22752 4250 22808
rect 4306 22752 5446 22808
rect 5502 22752 5507 22808
rect 3601 22750 5507 22752
rect 3601 22747 3667 22750
rect 4245 22747 4311 22750
rect 5441 22747 5507 22750
rect 4153 22676 4219 22677
rect 4102 22612 4108 22676
rect 4172 22674 4219 22676
rect 4172 22672 4264 22674
rect 4214 22616 4264 22672
rect 4172 22614 4264 22616
rect 4172 22612 4219 22614
rect 4153 22611 4219 22612
rect 4889 22540 4955 22541
rect 5257 22540 5323 22541
rect 4838 22476 4844 22540
rect 4908 22538 4955 22540
rect 4908 22536 5000 22538
rect 4950 22480 5000 22536
rect 4908 22478 5000 22480
rect 4908 22476 4955 22478
rect 5206 22476 5212 22540
rect 5276 22538 5323 22540
rect 5276 22536 5368 22538
rect 5318 22480 5368 22536
rect 5276 22478 5368 22480
rect 5276 22476 5323 22478
rect 4889 22475 4955 22476
rect 5257 22475 5323 22476
rect 2497 22402 2563 22405
rect 4521 22402 4587 22405
rect 2497 22400 4587 22402
rect 2497 22344 2502 22400
rect 2558 22344 4526 22400
rect 4582 22344 4587 22400
rect 2497 22342 4587 22344
rect 2497 22339 2563 22342
rect 4521 22339 4587 22342
rect 11145 22402 11211 22405
rect 13629 22402 13695 22405
rect 11145 22400 13695 22402
rect 11145 22344 11150 22400
rect 11206 22344 13634 22400
rect 13690 22344 13695 22400
rect 11145 22342 13695 22344
rect 11145 22339 11211 22342
rect 13629 22339 13695 22342
rect 5436 22336 5756 22337
rect 5436 22272 5444 22336
rect 5508 22272 5524 22336
rect 5588 22272 5604 22336
rect 5668 22272 5684 22336
rect 5748 22272 5756 22336
rect 5436 22271 5756 22272
rect 14422 22336 14742 22337
rect 14422 22272 14430 22336
rect 14494 22272 14510 22336
rect 14574 22272 14590 22336
rect 14654 22272 14670 22336
rect 14734 22272 14742 22336
rect 14422 22271 14742 22272
rect 19517 22266 19583 22269
rect 19977 22266 20043 22269
rect 19517 22264 20043 22266
rect 19517 22208 19522 22264
rect 19578 22208 19982 22264
rect 20038 22208 20043 22264
rect 19517 22206 20043 22208
rect 22050 22266 22110 22886
rect 22502 22884 22508 22948
rect 22572 22946 22578 22948
rect 24393 22946 24459 22949
rect 22572 22944 24459 22946
rect 22572 22888 24398 22944
rect 24454 22888 24459 22944
rect 22572 22886 24459 22888
rect 22572 22884 22578 22886
rect 24393 22883 24459 22886
rect 23407 22336 23727 22337
rect 23407 22272 23415 22336
rect 23479 22272 23495 22336
rect 23559 22272 23575 22336
rect 23639 22272 23655 22336
rect 23719 22272 23727 22336
rect 23407 22271 23727 22272
rect 22185 22266 22251 22269
rect 22050 22264 22251 22266
rect 22050 22208 22190 22264
rect 22246 22208 22251 22264
rect 22050 22206 22251 22208
rect 19517 22203 19583 22206
rect 19977 22203 20043 22206
rect 22185 22203 22251 22206
rect 9397 22130 9463 22133
rect 10409 22130 10475 22133
rect 9397 22128 10475 22130
rect 9397 22072 9402 22128
rect 9458 22072 10414 22128
rect 10470 22072 10475 22128
rect 9397 22070 10475 22072
rect 9397 22067 9463 22070
rect 10409 22067 10475 22070
rect 2865 21994 2931 21997
rect 11237 21994 11303 21997
rect 2865 21992 11303 21994
rect 2865 21936 2870 21992
rect 2926 21936 11242 21992
rect 11298 21936 11303 21992
rect 2865 21934 11303 21936
rect 2865 21931 2931 21934
rect 11237 21931 11303 21934
rect 2589 21858 2655 21861
rect 6310 21858 6316 21860
rect 2589 21856 6316 21858
rect 2589 21800 2594 21856
rect 2650 21800 6316 21856
rect 2589 21798 6316 21800
rect 2589 21795 2655 21798
rect 6310 21796 6316 21798
rect 6380 21796 6386 21860
rect 7557 21858 7623 21861
rect 7925 21858 7991 21861
rect 7557 21856 7991 21858
rect 7557 21800 7562 21856
rect 7618 21800 7930 21856
rect 7986 21800 7991 21856
rect 7557 21798 7991 21800
rect 7557 21795 7623 21798
rect 7925 21795 7991 21798
rect 8293 21858 8359 21861
rect 8937 21858 9003 21861
rect 18229 21860 18295 21861
rect 18229 21858 18276 21860
rect 8293 21856 9003 21858
rect 8293 21800 8298 21856
rect 8354 21800 8942 21856
rect 8998 21800 9003 21856
rect 8293 21798 9003 21800
rect 18184 21856 18276 21858
rect 18184 21800 18234 21856
rect 18184 21798 18276 21800
rect 8293 21795 8359 21798
rect 8937 21795 9003 21798
rect 18229 21796 18276 21798
rect 18340 21796 18346 21860
rect 18229 21795 18295 21796
rect 9929 21792 10249 21793
rect 9929 21728 9937 21792
rect 10001 21728 10017 21792
rect 10081 21728 10097 21792
rect 10161 21728 10177 21792
rect 10241 21728 10249 21792
rect 9929 21727 10249 21728
rect 18914 21792 19234 21793
rect 18914 21728 18922 21792
rect 18986 21728 19002 21792
rect 19066 21728 19082 21792
rect 19146 21728 19162 21792
rect 19226 21728 19234 21792
rect 18914 21727 19234 21728
rect 3969 21722 4035 21725
rect 7557 21722 7623 21725
rect 3969 21720 7623 21722
rect 3969 21664 3974 21720
rect 4030 21664 7562 21720
rect 7618 21664 7623 21720
rect 3969 21662 7623 21664
rect 3969 21659 4035 21662
rect 7557 21659 7623 21662
rect 19793 21722 19859 21725
rect 25865 21722 25931 21725
rect 26141 21722 26207 21725
rect 19793 21720 20178 21722
rect 19793 21664 19798 21720
rect 19854 21664 20178 21720
rect 19793 21662 20178 21664
rect 19793 21659 19859 21662
rect 3233 21586 3299 21589
rect 7465 21586 7531 21589
rect 3233 21584 7531 21586
rect 3233 21528 3238 21584
rect 3294 21528 7470 21584
rect 7526 21528 7531 21584
rect 3233 21526 7531 21528
rect 3233 21523 3299 21526
rect 7465 21523 7531 21526
rect 10593 21586 10659 21589
rect 15653 21586 15719 21589
rect 10593 21584 15719 21586
rect 10593 21528 10598 21584
rect 10654 21528 15658 21584
rect 15714 21528 15719 21584
rect 10593 21526 15719 21528
rect 10593 21523 10659 21526
rect 15653 21523 15719 21526
rect 19701 21586 19767 21589
rect 19885 21586 19951 21589
rect 19701 21584 19951 21586
rect 19701 21528 19706 21584
rect 19762 21528 19890 21584
rect 19946 21528 19951 21584
rect 19701 21526 19951 21528
rect 20118 21586 20178 21662
rect 25865 21720 26207 21722
rect 25865 21664 25870 21720
rect 25926 21664 26146 21720
rect 26202 21664 26207 21720
rect 25865 21662 26207 21664
rect 25865 21659 25931 21662
rect 26141 21659 26207 21662
rect 20621 21586 20687 21589
rect 20118 21584 20687 21586
rect 20118 21528 20626 21584
rect 20682 21528 20687 21584
rect 20118 21526 20687 21528
rect 19701 21523 19767 21526
rect 19885 21523 19951 21526
rect 20621 21523 20687 21526
rect 5073 21450 5139 21453
rect 5206 21450 5212 21452
rect 5073 21448 5212 21450
rect 5073 21392 5078 21448
rect 5134 21392 5212 21448
rect 5073 21390 5212 21392
rect 5073 21387 5139 21390
rect 5206 21388 5212 21390
rect 5276 21388 5282 21452
rect 6637 21450 6703 21453
rect 7230 21450 7236 21452
rect 6637 21448 7236 21450
rect 6637 21392 6642 21448
rect 6698 21392 7236 21448
rect 6637 21390 7236 21392
rect 6637 21387 6703 21390
rect 7230 21388 7236 21390
rect 7300 21388 7306 21452
rect 9765 21450 9831 21453
rect 10317 21450 10383 21453
rect 15009 21452 15075 21453
rect 14958 21450 14964 21452
rect 9765 21448 10383 21450
rect 9765 21392 9770 21448
rect 9826 21392 10322 21448
rect 10378 21392 10383 21448
rect 9765 21390 10383 21392
rect 14918 21390 14964 21450
rect 15028 21448 15075 21452
rect 15070 21392 15075 21448
rect 9765 21387 9831 21390
rect 10317 21387 10383 21390
rect 14958 21388 14964 21390
rect 15028 21388 15075 21392
rect 15009 21387 15075 21388
rect 4889 21314 4955 21317
rect 5206 21314 5212 21316
rect 4889 21312 5212 21314
rect 4889 21256 4894 21312
rect 4950 21256 5212 21312
rect 4889 21254 5212 21256
rect 4889 21251 4955 21254
rect 5206 21252 5212 21254
rect 5276 21252 5282 21316
rect 5436 21248 5756 21249
rect 5436 21184 5444 21248
rect 5508 21184 5524 21248
rect 5588 21184 5604 21248
rect 5668 21184 5684 21248
rect 5748 21184 5756 21248
rect 5436 21183 5756 21184
rect 14422 21248 14742 21249
rect 14422 21184 14430 21248
rect 14494 21184 14510 21248
rect 14574 21184 14590 21248
rect 14654 21184 14670 21248
rect 14734 21184 14742 21248
rect 14422 21183 14742 21184
rect 23407 21248 23727 21249
rect 23407 21184 23415 21248
rect 23479 21184 23495 21248
rect 23559 21184 23575 21248
rect 23639 21184 23655 21248
rect 23719 21184 23727 21248
rect 23407 21183 23727 21184
rect 2681 21042 2747 21045
rect 6126 21042 6132 21044
rect 2681 21040 6132 21042
rect 2681 20984 2686 21040
rect 2742 20984 6132 21040
rect 2681 20982 6132 20984
rect 2681 20979 2747 20982
rect 6126 20980 6132 20982
rect 6196 20980 6202 21044
rect 13077 21042 13143 21045
rect 13997 21044 14063 21045
rect 13670 21042 13676 21044
rect 13077 21040 13676 21042
rect 13077 20984 13082 21040
rect 13138 20984 13676 21040
rect 13077 20982 13676 20984
rect 13077 20979 13143 20982
rect 13670 20980 13676 20982
rect 13740 20980 13746 21044
rect 13997 21040 14044 21044
rect 14108 21042 14114 21044
rect 13997 20984 14002 21040
rect 13997 20980 14044 20984
rect 14108 20982 14154 21042
rect 14108 20980 14114 20982
rect 13997 20979 14063 20980
rect 3141 20906 3207 20909
rect 9622 20906 9628 20908
rect 3141 20904 9628 20906
rect 3141 20848 3146 20904
rect 3202 20848 9628 20904
rect 3141 20846 9628 20848
rect 3141 20843 3207 20846
rect 9622 20844 9628 20846
rect 9692 20844 9698 20908
rect 9949 20906 10015 20909
rect 10869 20906 10935 20909
rect 11278 20906 11284 20908
rect 9949 20904 11284 20906
rect 9949 20848 9954 20904
rect 10010 20848 10874 20904
rect 10930 20848 11284 20904
rect 9949 20846 11284 20848
rect 9949 20843 10015 20846
rect 10869 20843 10935 20846
rect 11278 20844 11284 20846
rect 11348 20844 11354 20908
rect 2221 20770 2287 20773
rect 3233 20770 3299 20773
rect 9254 20770 9260 20772
rect 2221 20768 9260 20770
rect 2221 20712 2226 20768
rect 2282 20712 3238 20768
rect 3294 20712 9260 20768
rect 2221 20710 9260 20712
rect 2221 20707 2287 20710
rect 3233 20707 3299 20710
rect 9254 20708 9260 20710
rect 9324 20708 9330 20772
rect 21817 20770 21883 20773
rect 21950 20770 21956 20772
rect 21817 20768 21956 20770
rect 21817 20712 21822 20768
rect 21878 20712 21956 20768
rect 21817 20710 21956 20712
rect 21817 20707 21883 20710
rect 21950 20708 21956 20710
rect 22020 20708 22026 20772
rect 22134 20708 22140 20772
rect 22204 20770 22210 20772
rect 22277 20770 22343 20773
rect 22204 20768 22343 20770
rect 22204 20712 22282 20768
rect 22338 20712 22343 20768
rect 22204 20710 22343 20712
rect 22204 20708 22210 20710
rect 22277 20707 22343 20710
rect 9929 20704 10249 20705
rect 9929 20640 9937 20704
rect 10001 20640 10017 20704
rect 10081 20640 10097 20704
rect 10161 20640 10177 20704
rect 10241 20640 10249 20704
rect 9929 20639 10249 20640
rect 18914 20704 19234 20705
rect 18914 20640 18922 20704
rect 18986 20640 19002 20704
rect 19066 20640 19082 20704
rect 19146 20640 19162 20704
rect 19226 20640 19234 20704
rect 18914 20639 19234 20640
rect 4838 20572 4844 20636
rect 4908 20634 4914 20636
rect 5349 20634 5415 20637
rect 4908 20632 5415 20634
rect 4908 20576 5354 20632
rect 5410 20576 5415 20632
rect 4908 20574 5415 20576
rect 4908 20572 4914 20574
rect 5349 20571 5415 20574
rect 6177 20634 6243 20637
rect 7189 20634 7255 20637
rect 6177 20632 7255 20634
rect 6177 20576 6182 20632
rect 6238 20576 7194 20632
rect 7250 20576 7255 20632
rect 6177 20574 7255 20576
rect 6177 20571 6243 20574
rect 7189 20571 7255 20574
rect 8661 20634 8727 20637
rect 9765 20634 9831 20637
rect 8661 20632 9831 20634
rect 8661 20576 8666 20632
rect 8722 20576 9770 20632
rect 9826 20576 9831 20632
rect 8661 20574 9831 20576
rect 8661 20571 8727 20574
rect 9765 20571 9831 20574
rect 2865 20498 2931 20501
rect 7966 20498 7972 20500
rect 2865 20496 7972 20498
rect 2865 20440 2870 20496
rect 2926 20440 7972 20496
rect 2865 20438 7972 20440
rect 2865 20435 2931 20438
rect 7966 20436 7972 20438
rect 8036 20436 8042 20500
rect 12801 20498 12867 20501
rect 17769 20498 17835 20501
rect 12801 20496 17835 20498
rect 12801 20440 12806 20496
rect 12862 20440 17774 20496
rect 17830 20440 17835 20496
rect 12801 20438 17835 20440
rect 12801 20435 12867 20438
rect 17769 20435 17835 20438
rect 3601 20364 3667 20365
rect 3550 20300 3556 20364
rect 3620 20362 3667 20364
rect 4153 20362 4219 20365
rect 5901 20362 5967 20365
rect 3620 20360 3712 20362
rect 3662 20304 3712 20360
rect 3620 20302 3712 20304
rect 4153 20360 5967 20362
rect 4153 20304 4158 20360
rect 4214 20304 5906 20360
rect 5962 20304 5967 20360
rect 4153 20302 5967 20304
rect 3620 20300 3667 20302
rect 3601 20299 3667 20300
rect 4153 20299 4219 20302
rect 5901 20299 5967 20302
rect 7281 20362 7347 20365
rect 10685 20362 10751 20365
rect 12341 20362 12407 20365
rect 7281 20360 12407 20362
rect 7281 20304 7286 20360
rect 7342 20304 10690 20360
rect 10746 20304 12346 20360
rect 12402 20304 12407 20360
rect 7281 20302 12407 20304
rect 7281 20299 7347 20302
rect 10685 20299 10751 20302
rect 12341 20299 12407 20302
rect 2589 20226 2655 20229
rect 4153 20226 4219 20229
rect 2589 20224 4219 20226
rect 2589 20168 2594 20224
rect 2650 20168 4158 20224
rect 4214 20168 4219 20224
rect 2589 20166 4219 20168
rect 2589 20163 2655 20166
rect 4153 20163 4219 20166
rect 5436 20160 5756 20161
rect 5436 20096 5444 20160
rect 5508 20096 5524 20160
rect 5588 20096 5604 20160
rect 5668 20096 5684 20160
rect 5748 20096 5756 20160
rect 5436 20095 5756 20096
rect 14422 20160 14742 20161
rect 14422 20096 14430 20160
rect 14494 20096 14510 20160
rect 14574 20096 14590 20160
rect 14654 20096 14670 20160
rect 14734 20096 14742 20160
rect 14422 20095 14742 20096
rect 23407 20160 23727 20161
rect 23407 20096 23415 20160
rect 23479 20096 23495 20160
rect 23559 20096 23575 20160
rect 23639 20096 23655 20160
rect 23719 20096 23727 20160
rect 23407 20095 23727 20096
rect 13486 20028 13492 20092
rect 13556 20090 13562 20092
rect 14181 20090 14247 20093
rect 13556 20088 14247 20090
rect 13556 20032 14186 20088
rect 14242 20032 14247 20088
rect 13556 20030 14247 20032
rect 13556 20028 13562 20030
rect 14181 20027 14247 20030
rect 2497 19954 2563 19957
rect 7782 19954 7788 19956
rect 2497 19952 7788 19954
rect 2497 19896 2502 19952
rect 2558 19896 7788 19952
rect 2497 19894 7788 19896
rect 2497 19891 2563 19894
rect 7782 19892 7788 19894
rect 7852 19954 7858 19956
rect 7925 19954 7991 19957
rect 7852 19952 7991 19954
rect 7852 19896 7930 19952
rect 7986 19896 7991 19952
rect 7852 19894 7991 19896
rect 7852 19892 7858 19894
rect 7925 19891 7991 19894
rect 8109 19956 8175 19957
rect 8109 19952 8156 19956
rect 8220 19954 8226 19956
rect 14365 19954 14431 19957
rect 15929 19956 15995 19957
rect 15878 19954 15884 19956
rect 8109 19896 8114 19952
rect 8109 19892 8156 19896
rect 8220 19894 8266 19954
rect 14365 19952 15884 19954
rect 15948 19952 15995 19956
rect 14365 19896 14370 19952
rect 14426 19896 15884 19952
rect 15990 19896 15995 19952
rect 14365 19894 15884 19896
rect 8220 19892 8226 19894
rect 8109 19891 8175 19892
rect 14365 19891 14431 19894
rect 15878 19892 15884 19894
rect 15948 19892 15995 19896
rect 15929 19891 15995 19892
rect 18321 19954 18387 19957
rect 18454 19954 18460 19956
rect 18321 19952 18460 19954
rect 18321 19896 18326 19952
rect 18382 19896 18460 19952
rect 18321 19894 18460 19896
rect 18321 19891 18387 19894
rect 18454 19892 18460 19894
rect 18524 19892 18530 19956
rect 3601 19818 3667 19821
rect 14089 19818 14155 19821
rect 16430 19818 16436 19820
rect 3601 19816 6378 19818
rect 3601 19760 3606 19816
rect 3662 19760 6378 19816
rect 3601 19758 6378 19760
rect 3601 19755 3667 19758
rect 3601 19682 3667 19685
rect 5942 19682 5948 19684
rect 3601 19680 5948 19682
rect 3601 19624 3606 19680
rect 3662 19624 5948 19680
rect 3601 19622 5948 19624
rect 3601 19619 3667 19622
rect 5942 19620 5948 19622
rect 6012 19620 6018 19684
rect 6318 19682 6378 19758
rect 14089 19816 16436 19818
rect 14089 19760 14094 19816
rect 14150 19760 16436 19816
rect 14089 19758 16436 19760
rect 14089 19755 14155 19758
rect 16430 19756 16436 19758
rect 16500 19756 16506 19820
rect 19149 19818 19215 19821
rect 18784 19816 19215 19818
rect 18784 19760 19154 19816
rect 19210 19760 19215 19816
rect 18784 19758 19215 19760
rect 7373 19682 7439 19685
rect 6318 19680 7439 19682
rect 6318 19624 7378 19680
rect 7434 19624 7439 19680
rect 6318 19622 7439 19624
rect 7373 19619 7439 19622
rect 12985 19682 13051 19685
rect 14181 19682 14247 19685
rect 12985 19680 14247 19682
rect 12985 19624 12990 19680
rect 13046 19624 14186 19680
rect 14242 19624 14247 19680
rect 12985 19622 14247 19624
rect 12985 19619 13051 19622
rect 14181 19619 14247 19622
rect 14641 19682 14707 19685
rect 15142 19682 15148 19684
rect 14641 19680 15148 19682
rect 14641 19624 14646 19680
rect 14702 19624 15148 19680
rect 14641 19622 15148 19624
rect 14641 19619 14707 19622
rect 15142 19620 15148 19622
rect 15212 19620 15218 19684
rect 9929 19616 10249 19617
rect 9929 19552 9937 19616
rect 10001 19552 10017 19616
rect 10081 19552 10097 19616
rect 10161 19552 10177 19616
rect 10241 19552 10249 19616
rect 9929 19551 10249 19552
rect 3601 19546 3667 19549
rect 8661 19546 8727 19549
rect 13445 19548 13511 19549
rect 13445 19546 13492 19548
rect 3601 19544 8727 19546
rect 3601 19488 3606 19544
rect 3662 19488 8666 19544
rect 8722 19488 8727 19544
rect 3601 19486 8727 19488
rect 13400 19544 13492 19546
rect 13400 19488 13450 19544
rect 13400 19486 13492 19488
rect 3601 19483 3667 19486
rect 8661 19483 8727 19486
rect 13445 19484 13492 19486
rect 13556 19484 13562 19548
rect 13905 19544 13971 19549
rect 13905 19488 13910 19544
rect 13966 19488 13971 19544
rect 13445 19483 13511 19484
rect 13905 19483 13971 19488
rect 2681 19410 2747 19413
rect 7005 19410 7071 19413
rect 2681 19408 7071 19410
rect 2681 19352 2686 19408
rect 2742 19352 7010 19408
rect 7066 19352 7071 19408
rect 2681 19350 7071 19352
rect 2681 19347 2747 19350
rect 7005 19347 7071 19350
rect 8109 19412 8175 19413
rect 8109 19408 8156 19412
rect 8220 19410 8226 19412
rect 8109 19352 8114 19408
rect 8109 19348 8156 19352
rect 8220 19350 8266 19410
rect 8220 19348 8226 19350
rect 8109 19347 8175 19348
rect 13908 19277 13968 19483
rect 18784 19410 18844 19758
rect 19149 19755 19215 19758
rect 25957 19682 26023 19685
rect 22188 19680 26023 19682
rect 22188 19624 25962 19680
rect 26018 19624 26023 19680
rect 22188 19622 26023 19624
rect 18914 19616 19234 19617
rect 18914 19552 18922 19616
rect 18986 19552 19002 19616
rect 19066 19552 19082 19616
rect 19146 19552 19162 19616
rect 19226 19552 19234 19616
rect 18914 19551 19234 19552
rect 22188 19549 22248 19622
rect 25957 19619 26023 19622
rect 22185 19544 22251 19549
rect 22185 19488 22190 19544
rect 22246 19488 22251 19544
rect 22185 19483 22251 19488
rect 22369 19546 22435 19549
rect 22645 19546 22711 19549
rect 22369 19544 22711 19546
rect 22369 19488 22374 19544
rect 22430 19488 22650 19544
rect 22706 19488 22711 19544
rect 22369 19486 22711 19488
rect 22369 19483 22435 19486
rect 22645 19483 22711 19486
rect 24485 19546 24551 19549
rect 24669 19546 24735 19549
rect 25773 19546 25839 19549
rect 24485 19544 25839 19546
rect 24485 19488 24490 19544
rect 24546 19488 24674 19544
rect 24730 19488 25778 19544
rect 25834 19488 25839 19544
rect 24485 19486 25839 19488
rect 24485 19483 24551 19486
rect 24669 19483 24735 19486
rect 25773 19483 25839 19486
rect 27245 19546 27311 19549
rect 28373 19546 29173 19576
rect 27245 19544 29173 19546
rect 27245 19488 27250 19544
rect 27306 19488 29173 19544
rect 27245 19486 29173 19488
rect 27245 19483 27311 19486
rect 28373 19456 29173 19486
rect 18965 19410 19031 19413
rect 18784 19408 19031 19410
rect 15469 19348 15535 19353
rect 18784 19352 18970 19408
rect 19026 19352 19031 19408
rect 18784 19350 19031 19352
rect 15469 19292 15474 19348
rect 15530 19308 15535 19348
rect 18965 19347 19031 19350
rect 22001 19410 22067 19413
rect 22645 19410 22711 19413
rect 22001 19408 22711 19410
rect 22001 19352 22006 19408
rect 22062 19352 22650 19408
rect 22706 19352 22711 19408
rect 22001 19350 22711 19352
rect 22001 19347 22067 19350
rect 22645 19347 22711 19350
rect 22829 19412 22895 19413
rect 22829 19408 22876 19412
rect 22940 19410 22946 19412
rect 22829 19352 22834 19408
rect 22829 19348 22876 19352
rect 22940 19350 22986 19410
rect 22940 19348 22946 19350
rect 22829 19347 22895 19348
rect 15530 19292 15946 19308
rect 15469 19287 15946 19292
rect 2589 19274 2655 19277
rect 2998 19274 3004 19276
rect 2589 19272 3004 19274
rect 2589 19216 2594 19272
rect 2650 19216 3004 19272
rect 2589 19214 3004 19216
rect 2589 19211 2655 19214
rect 2998 19212 3004 19214
rect 3068 19212 3074 19276
rect 4429 19274 4495 19277
rect 8753 19274 8819 19277
rect 4429 19272 8819 19274
rect 4429 19216 4434 19272
rect 4490 19216 8758 19272
rect 8814 19216 8819 19272
rect 4429 19214 8819 19216
rect 4429 19211 4495 19214
rect 8753 19211 8819 19214
rect 10777 19274 10843 19277
rect 11094 19274 11100 19276
rect 10777 19272 11100 19274
rect 10777 19216 10782 19272
rect 10838 19216 11100 19272
rect 10777 19214 11100 19216
rect 10777 19211 10843 19214
rect 11094 19212 11100 19214
rect 11164 19212 11170 19276
rect 13905 19272 13971 19277
rect 14825 19274 14891 19277
rect 13905 19216 13910 19272
rect 13966 19216 13971 19272
rect 13905 19211 13971 19216
rect 14782 19272 14891 19274
rect 14782 19216 14830 19272
rect 14886 19240 14891 19272
rect 15472 19274 15946 19287
rect 16246 19274 16252 19276
rect 15472 19248 16252 19274
rect 14886 19216 15210 19240
rect 14782 19180 15210 19216
rect 15886 19214 16252 19248
rect 16246 19212 16252 19214
rect 16316 19212 16322 19276
rect 16481 19274 16547 19277
rect 16614 19274 16620 19276
rect 16481 19272 16620 19274
rect 16481 19216 16486 19272
rect 16542 19216 16620 19272
rect 16481 19214 16620 19216
rect 16481 19211 16547 19214
rect 16614 19212 16620 19214
rect 16684 19212 16690 19276
rect 18781 19274 18847 19277
rect 20069 19274 20135 19277
rect 18781 19272 20135 19274
rect 18781 19216 18786 19272
rect 18842 19216 20074 19272
rect 20130 19216 20135 19272
rect 18781 19214 20135 19216
rect 18781 19211 18847 19214
rect 20069 19211 20135 19214
rect 20345 19274 20411 19277
rect 23657 19274 23723 19277
rect 26233 19274 26299 19277
rect 20345 19272 22110 19274
rect 20345 19216 20350 19272
rect 20406 19216 22110 19272
rect 20345 19214 22110 19216
rect 20345 19211 20411 19214
rect 2681 19138 2747 19141
rect 5257 19138 5323 19141
rect 2681 19136 5323 19138
rect 2681 19080 2686 19136
rect 2742 19080 5262 19136
rect 5318 19080 5323 19136
rect 2681 19078 5323 19080
rect 2681 19075 2747 19078
rect 5257 19075 5323 19078
rect 7281 19138 7347 19141
rect 8150 19138 8156 19140
rect 7281 19136 8156 19138
rect 7281 19080 7286 19136
rect 7342 19080 8156 19136
rect 7281 19078 8156 19080
rect 7281 19075 7347 19078
rect 8150 19076 8156 19078
rect 8220 19076 8226 19140
rect 8477 19138 8543 19141
rect 14089 19138 14155 19141
rect 8477 19136 14155 19138
rect 8477 19080 8482 19136
rect 8538 19080 14094 19136
rect 14150 19080 14155 19136
rect 8477 19078 14155 19080
rect 15150 19138 15210 19180
rect 15510 19138 15516 19140
rect 15150 19078 15516 19138
rect 8477 19075 8543 19078
rect 14089 19075 14155 19078
rect 15510 19076 15516 19078
rect 15580 19076 15586 19140
rect 15853 19138 15919 19141
rect 16798 19138 16804 19140
rect 15853 19136 16804 19138
rect 15853 19080 15858 19136
rect 15914 19080 16804 19136
rect 15853 19078 16804 19080
rect 15853 19075 15919 19078
rect 16798 19076 16804 19078
rect 16868 19076 16874 19140
rect 18873 19138 18939 19141
rect 21173 19138 21239 19141
rect 18873 19136 21239 19138
rect 18873 19080 18878 19136
rect 18934 19080 21178 19136
rect 21234 19080 21239 19136
rect 18873 19078 21239 19080
rect 22050 19138 22110 19214
rect 23657 19272 26299 19274
rect 23657 19216 23662 19272
rect 23718 19216 26238 19272
rect 26294 19216 26299 19272
rect 23657 19214 26299 19216
rect 23657 19211 23723 19214
rect 26233 19211 26299 19214
rect 23197 19138 23263 19141
rect 22050 19136 23263 19138
rect 22050 19080 23202 19136
rect 23258 19080 23263 19136
rect 22050 19078 23263 19080
rect 18873 19075 18939 19078
rect 21173 19075 21239 19078
rect 23197 19075 23263 19078
rect 5436 19072 5756 19073
rect 5436 19008 5444 19072
rect 5508 19008 5524 19072
rect 5588 19008 5604 19072
rect 5668 19008 5684 19072
rect 5748 19008 5756 19072
rect 5436 19007 5756 19008
rect 14422 19072 14742 19073
rect 14422 19008 14430 19072
rect 14494 19008 14510 19072
rect 14574 19008 14590 19072
rect 14654 19008 14670 19072
rect 14734 19008 14742 19072
rect 14422 19007 14742 19008
rect 23407 19072 23727 19073
rect 23407 19008 23415 19072
rect 23479 19008 23495 19072
rect 23559 19008 23575 19072
rect 23639 19008 23655 19072
rect 23719 19008 23727 19072
rect 23407 19007 23727 19008
rect 3141 19002 3207 19005
rect 4654 19002 4660 19004
rect 3141 19000 4660 19002
rect 3141 18944 3146 19000
rect 3202 18944 4660 19000
rect 3141 18942 4660 18944
rect 3141 18939 3207 18942
rect 4654 18940 4660 18942
rect 4724 18940 4730 19004
rect 5942 18940 5948 19004
rect 6012 19002 6018 19004
rect 7833 19002 7899 19005
rect 6012 19000 7899 19002
rect 6012 18944 7838 19000
rect 7894 18944 7899 19000
rect 6012 18942 7899 18944
rect 6012 18940 6018 18942
rect 7833 18939 7899 18942
rect 9622 18940 9628 19004
rect 9692 19002 9698 19004
rect 12014 19002 12020 19004
rect 9692 18942 12020 19002
rect 9692 18940 9698 18942
rect 12014 18940 12020 18942
rect 12084 18940 12090 19004
rect 12525 19002 12591 19005
rect 14181 19002 14247 19005
rect 12525 19000 14247 19002
rect 12525 18944 12530 19000
rect 12586 18944 14186 19000
rect 14242 18944 14247 19000
rect 12525 18942 14247 18944
rect 12525 18939 12591 18942
rect 14181 18939 14247 18942
rect 17902 18940 17908 19004
rect 17972 19002 17978 19004
rect 18965 19002 19031 19005
rect 17972 19000 19031 19002
rect 17972 18944 18970 19000
rect 19026 18944 19031 19000
rect 17972 18942 19031 18944
rect 17972 18940 17978 18942
rect 18965 18939 19031 18942
rect 1853 18866 1919 18869
rect 2630 18866 2636 18868
rect 1853 18864 2636 18866
rect 1853 18808 1858 18864
rect 1914 18808 2636 18864
rect 1853 18806 2636 18808
rect 1853 18803 1919 18806
rect 2630 18804 2636 18806
rect 2700 18804 2706 18868
rect 3141 18866 3207 18869
rect 6913 18866 6979 18869
rect 3141 18864 6979 18866
rect 3141 18808 3146 18864
rect 3202 18808 6918 18864
rect 6974 18808 6979 18864
rect 3141 18806 6979 18808
rect 3141 18803 3207 18806
rect 6913 18803 6979 18806
rect 10593 18866 10659 18869
rect 10726 18866 10732 18868
rect 10593 18864 10732 18866
rect 10593 18808 10598 18864
rect 10654 18808 10732 18864
rect 10593 18806 10732 18808
rect 10593 18803 10659 18806
rect 10726 18804 10732 18806
rect 10796 18804 10802 18868
rect 10961 18866 11027 18869
rect 11605 18866 11671 18869
rect 10961 18864 11671 18866
rect 10961 18808 10966 18864
rect 11022 18808 11610 18864
rect 11666 18808 11671 18864
rect 10961 18806 11671 18808
rect 10961 18803 11027 18806
rect 11605 18803 11671 18806
rect 13261 18866 13327 18869
rect 18086 18866 18092 18868
rect 13261 18864 18092 18866
rect 13261 18808 13266 18864
rect 13322 18808 18092 18864
rect 13261 18806 18092 18808
rect 13261 18803 13327 18806
rect 18086 18804 18092 18806
rect 18156 18866 18162 18868
rect 19057 18866 19123 18869
rect 18156 18864 19123 18866
rect 18156 18808 19062 18864
rect 19118 18808 19123 18864
rect 18156 18806 19123 18808
rect 18156 18804 18162 18806
rect 19057 18803 19123 18806
rect 2681 18730 2747 18733
rect 2814 18730 2820 18732
rect 2681 18728 2820 18730
rect 2681 18672 2686 18728
rect 2742 18672 2820 18728
rect 2681 18670 2820 18672
rect 2681 18667 2747 18670
rect 2814 18668 2820 18670
rect 2884 18668 2890 18732
rect 3182 18668 3188 18732
rect 3252 18730 3258 18732
rect 3417 18730 3483 18733
rect 3252 18728 3483 18730
rect 3252 18672 3422 18728
rect 3478 18672 3483 18728
rect 3252 18670 3483 18672
rect 3252 18668 3258 18670
rect 3417 18667 3483 18670
rect 4245 18730 4311 18733
rect 6913 18730 6979 18733
rect 4245 18728 6979 18730
rect 4245 18672 4250 18728
rect 4306 18672 6918 18728
rect 6974 18672 6979 18728
rect 4245 18670 6979 18672
rect 4245 18667 4311 18670
rect 6913 18667 6979 18670
rect 10869 18730 10935 18733
rect 11237 18730 11303 18733
rect 10869 18728 11303 18730
rect 10869 18672 10874 18728
rect 10930 18672 11242 18728
rect 11298 18672 11303 18728
rect 10869 18670 11303 18672
rect 10869 18667 10935 18670
rect 11237 18667 11303 18670
rect 14825 18730 14891 18733
rect 15510 18730 15516 18732
rect 14825 18728 15516 18730
rect 14825 18672 14830 18728
rect 14886 18672 15516 18728
rect 14825 18670 15516 18672
rect 14825 18667 14891 18670
rect 15510 18668 15516 18670
rect 15580 18668 15586 18732
rect 16062 18668 16068 18732
rect 16132 18730 16138 18732
rect 17033 18730 17099 18733
rect 17217 18730 17283 18733
rect 18873 18730 18939 18733
rect 16132 18728 17099 18730
rect 16132 18672 17038 18728
rect 17094 18672 17099 18728
rect 16132 18670 17099 18672
rect 16132 18668 16138 18670
rect 17033 18667 17099 18670
rect 17174 18728 17283 18730
rect 17174 18672 17222 18728
rect 17278 18672 17283 18728
rect 17174 18667 17283 18672
rect 18646 18728 18939 18730
rect 18646 18672 18878 18728
rect 18934 18672 18939 18728
rect 18646 18670 18939 18672
rect 3918 18532 3924 18596
rect 3988 18594 3994 18596
rect 4061 18594 4127 18597
rect 3988 18592 4127 18594
rect 3988 18536 4066 18592
rect 4122 18536 4127 18592
rect 3988 18534 4127 18536
rect 3988 18532 3994 18534
rect 4061 18531 4127 18534
rect 4613 18594 4679 18597
rect 5942 18594 5948 18596
rect 4613 18592 5948 18594
rect 4613 18536 4618 18592
rect 4674 18536 5948 18592
rect 4613 18534 5948 18536
rect 4613 18531 4679 18534
rect 5942 18532 5948 18534
rect 6012 18532 6018 18596
rect 6310 18532 6316 18596
rect 6380 18594 6386 18596
rect 8201 18594 8267 18597
rect 6380 18592 8267 18594
rect 6380 18536 8206 18592
rect 8262 18536 8267 18592
rect 6380 18534 8267 18536
rect 6380 18532 6386 18534
rect 8201 18531 8267 18534
rect 10685 18594 10751 18597
rect 10961 18594 11027 18597
rect 10685 18592 11027 18594
rect 10685 18536 10690 18592
rect 10746 18536 10966 18592
rect 11022 18536 11027 18592
rect 10685 18534 11027 18536
rect 10685 18531 10751 18534
rect 10961 18531 11027 18534
rect 12985 18594 13051 18597
rect 17174 18594 17234 18667
rect 12985 18592 17234 18594
rect 12985 18536 12990 18592
rect 13046 18536 17234 18592
rect 12985 18534 17234 18536
rect 12985 18531 13051 18534
rect 9929 18528 10249 18529
rect 9929 18464 9937 18528
rect 10001 18464 10017 18528
rect 10081 18464 10097 18528
rect 10161 18464 10177 18528
rect 10241 18464 10249 18528
rect 9929 18463 10249 18464
rect 4061 18458 4127 18461
rect 4061 18456 4538 18458
rect 4061 18400 4066 18456
rect 4122 18400 4538 18456
rect 4061 18398 4538 18400
rect 4061 18395 4127 18398
rect 3877 18322 3943 18325
rect 4286 18322 4292 18324
rect 3877 18320 4292 18322
rect 3877 18264 3882 18320
rect 3938 18264 4292 18320
rect 3877 18262 4292 18264
rect 3877 18259 3943 18262
rect 4286 18260 4292 18262
rect 4356 18260 4362 18324
rect 4478 18322 4538 18398
rect 5206 18396 5212 18460
rect 5276 18458 5282 18460
rect 7005 18458 7071 18461
rect 5276 18456 7071 18458
rect 5276 18400 7010 18456
rect 7066 18400 7071 18456
rect 5276 18398 7071 18400
rect 5276 18396 5282 18398
rect 7005 18395 7071 18398
rect 7782 18396 7788 18460
rect 7852 18458 7858 18460
rect 7925 18458 7991 18461
rect 7852 18456 7991 18458
rect 7852 18400 7930 18456
rect 7986 18400 7991 18456
rect 7852 18398 7991 18400
rect 7852 18396 7858 18398
rect 7925 18395 7991 18398
rect 10409 18458 10475 18461
rect 10910 18458 10916 18460
rect 10409 18456 10916 18458
rect 10409 18400 10414 18456
rect 10470 18400 10916 18456
rect 10409 18398 10916 18400
rect 10409 18395 10475 18398
rect 10910 18396 10916 18398
rect 10980 18396 10986 18460
rect 12801 18458 12867 18461
rect 16205 18458 16271 18461
rect 12801 18456 16271 18458
rect 12801 18400 12806 18456
rect 12862 18400 16210 18456
rect 16266 18400 16271 18456
rect 12801 18398 16271 18400
rect 12801 18395 12867 18398
rect 16205 18395 16271 18398
rect 18229 18460 18295 18461
rect 18229 18456 18276 18460
rect 18340 18458 18346 18460
rect 18505 18458 18571 18461
rect 18646 18458 18706 18670
rect 18873 18667 18939 18670
rect 18914 18528 19234 18529
rect 18914 18464 18922 18528
rect 18986 18464 19002 18528
rect 19066 18464 19082 18528
rect 19146 18464 19162 18528
rect 19226 18464 19234 18528
rect 18914 18463 19234 18464
rect 18229 18400 18234 18456
rect 18229 18396 18276 18400
rect 18340 18398 18386 18458
rect 18505 18456 18706 18458
rect 18505 18400 18510 18456
rect 18566 18400 18706 18456
rect 18505 18398 18706 18400
rect 18340 18396 18346 18398
rect 18229 18395 18295 18396
rect 18505 18395 18571 18398
rect 5533 18322 5599 18325
rect 4478 18320 5599 18322
rect 4478 18264 5538 18320
rect 5594 18264 5599 18320
rect 4478 18262 5599 18264
rect 5533 18259 5599 18262
rect 6494 18260 6500 18324
rect 6564 18322 6570 18324
rect 8017 18322 8083 18325
rect 6564 18320 8083 18322
rect 6564 18264 8022 18320
rect 8078 18264 8083 18320
rect 6564 18262 8083 18264
rect 6564 18260 6570 18262
rect 8017 18259 8083 18262
rect 13077 18322 13143 18325
rect 18873 18322 18939 18325
rect 13077 18320 18939 18322
rect 13077 18264 13082 18320
rect 13138 18264 18878 18320
rect 18934 18264 18939 18320
rect 13077 18262 18939 18264
rect 13077 18259 13143 18262
rect 18873 18259 18939 18262
rect 19517 18322 19583 18325
rect 22093 18322 22159 18325
rect 19517 18320 22159 18322
rect 19517 18264 19522 18320
rect 19578 18264 22098 18320
rect 22154 18264 22159 18320
rect 19517 18262 22159 18264
rect 19517 18259 19583 18262
rect 22093 18259 22159 18262
rect 4245 18186 4311 18189
rect 5022 18186 5028 18188
rect 4245 18184 5028 18186
rect 4245 18128 4250 18184
rect 4306 18128 5028 18184
rect 4245 18126 5028 18128
rect 4245 18123 4311 18126
rect 5022 18124 5028 18126
rect 5092 18124 5098 18188
rect 5206 18124 5212 18188
rect 5276 18186 5282 18188
rect 5441 18186 5507 18189
rect 5276 18184 5507 18186
rect 5276 18128 5446 18184
rect 5502 18128 5507 18184
rect 5276 18126 5507 18128
rect 5276 18124 5282 18126
rect 5441 18123 5507 18126
rect 10133 18186 10199 18189
rect 10358 18186 10364 18188
rect 10133 18184 10364 18186
rect 10133 18128 10138 18184
rect 10194 18128 10364 18184
rect 10133 18126 10364 18128
rect 10133 18123 10199 18126
rect 10358 18124 10364 18126
rect 10428 18124 10434 18188
rect 13670 18124 13676 18188
rect 13740 18186 13746 18188
rect 15101 18186 15167 18189
rect 13740 18184 15167 18186
rect 13740 18128 15106 18184
rect 15162 18128 15167 18184
rect 13740 18126 15167 18128
rect 13740 18124 13746 18126
rect 15101 18123 15167 18126
rect 16982 18124 16988 18188
rect 17052 18186 17058 18188
rect 17217 18186 17283 18189
rect 17052 18184 17283 18186
rect 17052 18128 17222 18184
rect 17278 18128 17283 18184
rect 17052 18126 17283 18128
rect 17052 18124 17058 18126
rect 17217 18123 17283 18126
rect 17585 18186 17651 18189
rect 18597 18186 18663 18189
rect 17585 18184 18663 18186
rect 17585 18128 17590 18184
rect 17646 18128 18602 18184
rect 18658 18128 18663 18184
rect 17585 18126 18663 18128
rect 17585 18123 17651 18126
rect 18597 18123 18663 18126
rect 10133 18050 10199 18053
rect 11237 18050 11303 18053
rect 10133 18048 11303 18050
rect 10133 17992 10138 18048
rect 10194 17992 11242 18048
rect 11298 17992 11303 18048
rect 10133 17990 11303 17992
rect 10133 17987 10199 17990
rect 11237 17987 11303 17990
rect 11462 17988 11468 18052
rect 11532 18050 11538 18052
rect 14089 18050 14155 18053
rect 11532 18048 14155 18050
rect 11532 17992 14094 18048
rect 14150 17992 14155 18048
rect 11532 17990 14155 17992
rect 11532 17988 11538 17990
rect 14089 17987 14155 17990
rect 15745 18050 15811 18053
rect 16798 18050 16804 18052
rect 15745 18048 16804 18050
rect 15745 17992 15750 18048
rect 15806 17992 16804 18048
rect 15745 17990 16804 17992
rect 15745 17987 15811 17990
rect 16798 17988 16804 17990
rect 16868 17988 16874 18052
rect 17401 18050 17467 18053
rect 18965 18050 19031 18053
rect 17401 18048 19031 18050
rect 17401 17992 17406 18048
rect 17462 17992 18970 18048
rect 19026 17992 19031 18048
rect 17401 17990 19031 17992
rect 17401 17987 17467 17990
rect 18965 17987 19031 17990
rect 5436 17984 5756 17985
rect 5436 17920 5444 17984
rect 5508 17920 5524 17984
rect 5588 17920 5604 17984
rect 5668 17920 5684 17984
rect 5748 17920 5756 17984
rect 5436 17919 5756 17920
rect 14422 17984 14742 17985
rect 14422 17920 14430 17984
rect 14494 17920 14510 17984
rect 14574 17920 14590 17984
rect 14654 17920 14670 17984
rect 14734 17920 14742 17984
rect 14422 17919 14742 17920
rect 23407 17984 23727 17985
rect 23407 17920 23415 17984
rect 23479 17920 23495 17984
rect 23559 17920 23575 17984
rect 23639 17920 23655 17984
rect 23719 17920 23727 17984
rect 23407 17919 23727 17920
rect 10041 17914 10107 17917
rect 10542 17914 10548 17916
rect 10041 17912 10548 17914
rect 10041 17856 10046 17912
rect 10102 17856 10548 17912
rect 10041 17854 10548 17856
rect 10041 17851 10107 17854
rect 10542 17852 10548 17854
rect 10612 17852 10618 17916
rect 17861 17914 17927 17917
rect 18137 17914 18203 17917
rect 17861 17912 18203 17914
rect 17861 17856 17866 17912
rect 17922 17856 18142 17912
rect 18198 17856 18203 17912
rect 17861 17854 18203 17856
rect 17861 17851 17927 17854
rect 18137 17851 18203 17854
rect 2814 17716 2820 17780
rect 2884 17778 2890 17780
rect 9581 17778 9647 17781
rect 2884 17776 9647 17778
rect 2884 17720 9586 17776
rect 9642 17720 9647 17776
rect 2884 17718 9647 17720
rect 2884 17716 2890 17718
rect 9581 17715 9647 17718
rect 13486 17716 13492 17780
rect 13556 17778 13562 17780
rect 16481 17778 16547 17781
rect 19057 17778 19123 17781
rect 13556 17776 19123 17778
rect 13556 17720 16486 17776
rect 16542 17720 19062 17776
rect 19118 17720 19123 17776
rect 13556 17718 19123 17720
rect 13556 17716 13562 17718
rect 16481 17715 16547 17718
rect 19057 17715 19123 17718
rect 21030 17716 21036 17780
rect 21100 17778 21106 17780
rect 24209 17778 24275 17781
rect 21100 17776 24275 17778
rect 21100 17720 24214 17776
rect 24270 17720 24275 17776
rect 21100 17718 24275 17720
rect 21100 17716 21106 17718
rect 24209 17715 24275 17718
rect 4705 17642 4771 17645
rect 4838 17642 4844 17644
rect 4705 17640 4844 17642
rect 4705 17584 4710 17640
rect 4766 17584 4844 17640
rect 4705 17582 4844 17584
rect 4705 17579 4771 17582
rect 4838 17580 4844 17582
rect 4908 17580 4914 17644
rect 15142 17580 15148 17644
rect 15212 17642 15218 17644
rect 21541 17642 21607 17645
rect 26785 17642 26851 17645
rect 15212 17640 21607 17642
rect 15212 17584 21546 17640
rect 21602 17584 21607 17640
rect 15212 17582 21607 17584
rect 15212 17580 15218 17582
rect 21541 17579 21607 17582
rect 26742 17640 26851 17642
rect 26742 17584 26790 17640
rect 26846 17584 26851 17640
rect 26742 17579 26851 17584
rect 11329 17506 11395 17509
rect 11462 17506 11468 17508
rect 11329 17504 11468 17506
rect 11329 17448 11334 17504
rect 11390 17448 11468 17504
rect 11329 17446 11468 17448
rect 11329 17443 11395 17446
rect 11462 17444 11468 17446
rect 11532 17444 11538 17508
rect 12617 17506 12683 17509
rect 12390 17504 12683 17506
rect 12390 17448 12622 17504
rect 12678 17448 12683 17504
rect 12390 17446 12683 17448
rect 9929 17440 10249 17441
rect 9929 17376 9937 17440
rect 10001 17376 10017 17440
rect 10081 17376 10097 17440
rect 10161 17376 10177 17440
rect 10241 17376 10249 17440
rect 9929 17375 10249 17376
rect 5257 17370 5323 17373
rect 7046 17370 7052 17372
rect 5257 17368 7052 17370
rect 5257 17312 5262 17368
rect 5318 17312 7052 17368
rect 5257 17310 7052 17312
rect 5257 17307 5323 17310
rect 7046 17308 7052 17310
rect 7116 17308 7122 17372
rect 12390 17370 12450 17446
rect 12617 17443 12683 17446
rect 16481 17506 16547 17509
rect 17350 17506 17356 17508
rect 16481 17504 17356 17506
rect 16481 17448 16486 17504
rect 16542 17448 17356 17504
rect 16481 17446 17356 17448
rect 16481 17443 16547 17446
rect 17350 17444 17356 17446
rect 17420 17444 17426 17508
rect 23013 17506 23079 17509
rect 22050 17504 23079 17506
rect 22050 17448 23018 17504
rect 23074 17448 23079 17504
rect 22050 17446 23079 17448
rect 18914 17440 19234 17441
rect 18914 17376 18922 17440
rect 18986 17376 19002 17440
rect 19066 17376 19082 17440
rect 19146 17376 19162 17440
rect 19226 17376 19234 17440
rect 18914 17375 19234 17376
rect 22050 17370 22110 17446
rect 23013 17443 23079 17446
rect 10734 17310 12450 17370
rect 21774 17310 22110 17370
rect 10734 17237 10794 17310
rect 10685 17232 10794 17237
rect 10685 17176 10690 17232
rect 10746 17176 10794 17232
rect 10685 17174 10794 17176
rect 12157 17234 12223 17237
rect 14038 17234 14044 17236
rect 12157 17232 14044 17234
rect 12157 17176 12162 17232
rect 12218 17176 14044 17232
rect 12157 17174 14044 17176
rect 10685 17171 10751 17174
rect 12157 17171 12223 17174
rect 14038 17172 14044 17174
rect 14108 17234 14114 17236
rect 14365 17234 14431 17237
rect 14108 17232 14431 17234
rect 14108 17176 14370 17232
rect 14426 17176 14431 17232
rect 14108 17174 14431 17176
rect 14108 17172 14114 17174
rect 14365 17171 14431 17174
rect 16757 17234 16823 17237
rect 17125 17234 17191 17237
rect 16757 17232 17191 17234
rect 16757 17176 16762 17232
rect 16818 17176 17130 17232
rect 17186 17176 17191 17232
rect 16757 17174 17191 17176
rect 16757 17171 16823 17174
rect 17125 17171 17191 17174
rect 20713 17234 20779 17237
rect 21081 17234 21147 17237
rect 20713 17232 21147 17234
rect 20713 17176 20718 17232
rect 20774 17176 21086 17232
rect 21142 17176 21147 17232
rect 20713 17174 21147 17176
rect 20713 17171 20779 17174
rect 21081 17171 21147 17174
rect 21541 17234 21607 17237
rect 21774 17234 21834 17310
rect 21541 17232 21834 17234
rect 21541 17176 21546 17232
rect 21602 17176 21834 17232
rect 21541 17174 21834 17176
rect 21541 17171 21607 17174
rect 7373 17100 7439 17101
rect 7373 17096 7420 17100
rect 7484 17098 7490 17100
rect 7373 17040 7378 17096
rect 7373 17036 7420 17040
rect 7484 17038 7530 17098
rect 7484 17036 7490 17038
rect 11830 17036 11836 17100
rect 11900 17098 11906 17100
rect 11973 17098 12039 17101
rect 11900 17096 12039 17098
rect 11900 17040 11978 17096
rect 12034 17040 12039 17096
rect 11900 17038 12039 17040
rect 11900 17036 11906 17038
rect 7373 17035 7439 17036
rect 11973 17035 12039 17038
rect 16849 17098 16915 17101
rect 18229 17100 18295 17101
rect 17166 17098 17172 17100
rect 16849 17096 17172 17098
rect 16849 17040 16854 17096
rect 16910 17040 17172 17096
rect 16849 17038 17172 17040
rect 16849 17035 16915 17038
rect 17166 17036 17172 17038
rect 17236 17036 17242 17100
rect 18229 17098 18276 17100
rect 18184 17096 18276 17098
rect 18184 17040 18234 17096
rect 18184 17038 18276 17040
rect 18229 17036 18276 17038
rect 18340 17036 18346 17100
rect 21817 17098 21883 17101
rect 23289 17098 23355 17101
rect 21817 17096 23355 17098
rect 21817 17040 21822 17096
rect 21878 17040 23294 17096
rect 23350 17040 23355 17096
rect 21817 17038 23355 17040
rect 18229 17035 18295 17036
rect 21817 17035 21883 17038
rect 23289 17035 23355 17038
rect 16798 16900 16804 16964
rect 16868 16962 16874 16964
rect 16941 16962 17007 16965
rect 18413 16964 18479 16965
rect 18413 16962 18460 16964
rect 16868 16960 17007 16962
rect 16868 16904 16946 16960
rect 17002 16904 17007 16960
rect 16868 16902 17007 16904
rect 18368 16960 18460 16962
rect 18368 16904 18418 16960
rect 18368 16902 18460 16904
rect 16868 16900 16874 16902
rect 16941 16899 17007 16902
rect 18413 16900 18460 16902
rect 18524 16900 18530 16964
rect 21173 16962 21239 16965
rect 23013 16962 23079 16965
rect 21173 16960 23079 16962
rect 21173 16904 21178 16960
rect 21234 16904 23018 16960
rect 23074 16904 23079 16960
rect 21173 16902 23079 16904
rect 18413 16899 18479 16900
rect 21173 16899 21239 16902
rect 23013 16899 23079 16902
rect 5436 16896 5756 16897
rect 5436 16832 5444 16896
rect 5508 16832 5524 16896
rect 5588 16832 5604 16896
rect 5668 16832 5684 16896
rect 5748 16832 5756 16896
rect 5436 16831 5756 16832
rect 14422 16896 14742 16897
rect 14422 16832 14430 16896
rect 14494 16832 14510 16896
rect 14574 16832 14590 16896
rect 14654 16832 14670 16896
rect 14734 16832 14742 16896
rect 14422 16831 14742 16832
rect 23407 16896 23727 16897
rect 23407 16832 23415 16896
rect 23479 16832 23495 16896
rect 23559 16832 23575 16896
rect 23639 16832 23655 16896
rect 23719 16832 23727 16896
rect 23407 16831 23727 16832
rect 15469 16826 15535 16829
rect 16246 16826 16252 16828
rect 15469 16824 16252 16826
rect 15469 16768 15474 16824
rect 15530 16768 16252 16824
rect 15469 16766 16252 16768
rect 15469 16763 15535 16766
rect 16246 16764 16252 16766
rect 16316 16764 16322 16828
rect 16389 16826 16455 16829
rect 18270 16826 18276 16828
rect 16389 16824 18276 16826
rect 16389 16768 16394 16824
rect 16450 16768 18276 16824
rect 16389 16766 18276 16768
rect 16389 16763 16455 16766
rect 18270 16764 18276 16766
rect 18340 16826 18346 16828
rect 18505 16826 18571 16829
rect 18340 16824 18571 16826
rect 18340 16768 18510 16824
rect 18566 16768 18571 16824
rect 18340 16766 18571 16768
rect 18340 16764 18346 16766
rect 18505 16763 18571 16766
rect 26601 16826 26667 16829
rect 26742 16826 26802 17579
rect 26601 16824 26802 16826
rect 26601 16768 26606 16824
rect 26662 16768 26802 16824
rect 26601 16766 26802 16768
rect 26601 16763 26667 16766
rect 15510 16628 15516 16692
rect 15580 16690 15586 16692
rect 15653 16690 15719 16693
rect 18965 16690 19031 16693
rect 15580 16688 19031 16690
rect 15580 16632 15658 16688
rect 15714 16632 18970 16688
rect 19026 16632 19031 16688
rect 15580 16630 19031 16632
rect 15580 16628 15586 16630
rect 15653 16627 15719 16630
rect 18965 16627 19031 16630
rect 22001 16690 22067 16693
rect 22686 16690 22692 16692
rect 22001 16688 22692 16690
rect 22001 16632 22006 16688
rect 22062 16632 22692 16688
rect 22001 16630 22692 16632
rect 22001 16627 22067 16630
rect 22686 16628 22692 16630
rect 22756 16628 22762 16692
rect 15929 16554 15995 16557
rect 18505 16554 18571 16557
rect 15929 16552 18571 16554
rect 15929 16496 15934 16552
rect 15990 16496 18510 16552
rect 18566 16496 18571 16552
rect 15929 16494 18571 16496
rect 15929 16491 15995 16494
rect 18505 16491 18571 16494
rect 13077 16418 13143 16421
rect 14825 16418 14891 16421
rect 13077 16416 14891 16418
rect 13077 16360 13082 16416
rect 13138 16360 14830 16416
rect 14886 16360 14891 16416
rect 13077 16358 14891 16360
rect 13077 16355 13143 16358
rect 14825 16355 14891 16358
rect 15745 16418 15811 16421
rect 16614 16418 16620 16420
rect 15745 16416 16620 16418
rect 15745 16360 15750 16416
rect 15806 16360 16620 16416
rect 15745 16358 16620 16360
rect 15745 16355 15811 16358
rect 16614 16356 16620 16358
rect 16684 16356 16690 16420
rect 22870 16356 22876 16420
rect 22940 16418 22946 16420
rect 23013 16418 23079 16421
rect 22940 16416 23079 16418
rect 22940 16360 23018 16416
rect 23074 16360 23079 16416
rect 22940 16358 23079 16360
rect 22940 16356 22946 16358
rect 23013 16355 23079 16358
rect 9929 16352 10249 16353
rect 9929 16288 9937 16352
rect 10001 16288 10017 16352
rect 10081 16288 10097 16352
rect 10161 16288 10177 16352
rect 10241 16288 10249 16352
rect 9929 16287 10249 16288
rect 18914 16352 19234 16353
rect 18914 16288 18922 16352
rect 18986 16288 19002 16352
rect 19066 16288 19082 16352
rect 19146 16288 19162 16352
rect 19226 16288 19234 16352
rect 18914 16287 19234 16288
rect 2773 16284 2839 16285
rect 2773 16282 2820 16284
rect 2728 16280 2820 16282
rect 2728 16224 2778 16280
rect 2728 16222 2820 16224
rect 2773 16220 2820 16222
rect 2884 16220 2890 16284
rect 11329 16282 11395 16285
rect 18638 16282 18644 16284
rect 11329 16280 18644 16282
rect 11329 16224 11334 16280
rect 11390 16224 18644 16280
rect 11329 16222 18644 16224
rect 2773 16219 2839 16220
rect 11329 16219 11395 16222
rect 18638 16220 18644 16222
rect 18708 16220 18714 16284
rect 12525 16146 12591 16149
rect 12390 16144 12591 16146
rect 12390 16088 12530 16144
rect 12586 16088 12591 16144
rect 12390 16086 12591 16088
rect 12249 15874 12315 15877
rect 12390 15874 12450 16086
rect 12525 16083 12591 16086
rect 13353 16146 13419 16149
rect 13813 16146 13879 16149
rect 13353 16144 13879 16146
rect 13353 16088 13358 16144
rect 13414 16088 13818 16144
rect 13874 16088 13879 16144
rect 13353 16086 13879 16088
rect 13353 16083 13419 16086
rect 13813 16083 13879 16086
rect 16246 16084 16252 16148
rect 16316 16146 16322 16148
rect 17217 16146 17283 16149
rect 16316 16144 17283 16146
rect 16316 16088 17222 16144
rect 17278 16088 17283 16144
rect 16316 16086 17283 16088
rect 16316 16084 16322 16086
rect 17217 16083 17283 16086
rect 14365 16010 14431 16013
rect 16614 16010 16620 16012
rect 14365 16008 16620 16010
rect 14365 15952 14370 16008
rect 14426 15952 16620 16008
rect 14365 15950 16620 15952
rect 14365 15947 14431 15950
rect 16614 15948 16620 15950
rect 16684 15948 16690 16012
rect 12249 15872 12450 15874
rect 12249 15816 12254 15872
rect 12310 15816 12450 15872
rect 12249 15814 12450 15816
rect 12249 15811 12315 15814
rect 5436 15808 5756 15809
rect 5436 15744 5444 15808
rect 5508 15744 5524 15808
rect 5588 15744 5604 15808
rect 5668 15744 5684 15808
rect 5748 15744 5756 15808
rect 5436 15743 5756 15744
rect 14422 15808 14742 15809
rect 14422 15744 14430 15808
rect 14494 15744 14510 15808
rect 14574 15744 14590 15808
rect 14654 15744 14670 15808
rect 14734 15744 14742 15808
rect 14422 15743 14742 15744
rect 23407 15808 23727 15809
rect 23407 15744 23415 15808
rect 23479 15744 23495 15808
rect 23559 15744 23575 15808
rect 23639 15744 23655 15808
rect 23719 15744 23727 15808
rect 23407 15743 23727 15744
rect 2405 15738 2471 15741
rect 3734 15738 3740 15740
rect 2405 15736 3740 15738
rect 2405 15680 2410 15736
rect 2466 15680 3740 15736
rect 2405 15678 3740 15680
rect 2405 15675 2471 15678
rect 3734 15676 3740 15678
rect 3804 15676 3810 15740
rect 12617 15738 12683 15741
rect 12617 15736 13002 15738
rect 12617 15680 12622 15736
rect 12678 15680 13002 15736
rect 12617 15678 13002 15680
rect 12617 15675 12683 15678
rect 1853 15602 1919 15605
rect 1853 15600 2514 15602
rect 1853 15544 1858 15600
rect 1914 15544 2514 15600
rect 1853 15542 2514 15544
rect 1853 15539 1919 15542
rect 2454 15466 2514 15542
rect 6678 15540 6684 15604
rect 6748 15602 6754 15604
rect 6821 15602 6887 15605
rect 6748 15600 6887 15602
rect 6748 15544 6826 15600
rect 6882 15544 6887 15600
rect 6748 15542 6887 15544
rect 12942 15602 13002 15678
rect 15101 15736 15167 15741
rect 15101 15680 15106 15736
rect 15162 15680 15167 15736
rect 15101 15675 15167 15680
rect 13077 15602 13143 15605
rect 12942 15600 13143 15602
rect 12942 15544 13082 15600
rect 13138 15544 13143 15600
rect 12942 15542 13143 15544
rect 6748 15540 6754 15542
rect 6821 15539 6887 15542
rect 13077 15539 13143 15542
rect 14641 15602 14707 15605
rect 15104 15602 15164 15675
rect 14641 15600 15164 15602
rect 14641 15544 14646 15600
rect 14702 15544 15164 15600
rect 14641 15542 15164 15544
rect 21081 15602 21147 15605
rect 26785 15602 26851 15605
rect 21081 15600 26851 15602
rect 21081 15544 21086 15600
rect 21142 15544 26790 15600
rect 26846 15544 26851 15600
rect 21081 15542 26851 15544
rect 14641 15539 14707 15542
rect 21081 15539 21147 15542
rect 26785 15539 26851 15542
rect 2681 15466 2747 15469
rect 2454 15464 2747 15466
rect 2454 15408 2686 15464
rect 2742 15408 2747 15464
rect 2454 15406 2747 15408
rect 2681 15403 2747 15406
rect 14549 15466 14615 15469
rect 23197 15468 23263 15469
rect 23197 15466 23244 15468
rect 14549 15464 21834 15466
rect 14549 15408 14554 15464
rect 14610 15408 21834 15464
rect 14549 15406 21834 15408
rect 23152 15464 23244 15466
rect 23152 15408 23202 15464
rect 23152 15406 23244 15408
rect 14549 15403 14615 15406
rect 3877 15330 3943 15333
rect 6310 15330 6316 15332
rect 3877 15328 6316 15330
rect 3877 15272 3882 15328
rect 3938 15272 6316 15328
rect 3877 15270 6316 15272
rect 3877 15267 3943 15270
rect 6310 15268 6316 15270
rect 6380 15268 6386 15332
rect 12709 15330 12775 15333
rect 10918 15328 12775 15330
rect 10918 15272 12714 15328
rect 12770 15272 12775 15328
rect 10918 15270 12775 15272
rect 9929 15264 10249 15265
rect 9929 15200 9937 15264
rect 10001 15200 10017 15264
rect 10081 15200 10097 15264
rect 10161 15200 10177 15264
rect 10241 15200 10249 15264
rect 9929 15199 10249 15200
rect 7925 15058 7991 15061
rect 8569 15058 8635 15061
rect 10918 15058 10978 15270
rect 12709 15267 12775 15270
rect 15377 15330 15443 15333
rect 17125 15330 17191 15333
rect 21774 15332 21834 15406
rect 23197 15404 23244 15406
rect 23308 15404 23314 15468
rect 23197 15403 23263 15404
rect 15377 15328 17191 15330
rect 15377 15272 15382 15328
rect 15438 15272 17130 15328
rect 17186 15272 17191 15328
rect 15377 15270 17191 15272
rect 15377 15267 15443 15270
rect 17125 15267 17191 15270
rect 21766 15268 21772 15332
rect 21836 15330 21842 15332
rect 22185 15330 22251 15333
rect 21836 15328 22251 15330
rect 21836 15272 22190 15328
rect 22246 15272 22251 15328
rect 21836 15270 22251 15272
rect 21836 15268 21842 15270
rect 22185 15267 22251 15270
rect 18914 15264 19234 15265
rect 18914 15200 18922 15264
rect 18986 15200 19002 15264
rect 19066 15200 19082 15264
rect 19146 15200 19162 15264
rect 19226 15200 19234 15264
rect 18914 15199 19234 15200
rect 15653 15194 15719 15197
rect 16205 15194 16271 15197
rect 15653 15192 16271 15194
rect 15653 15136 15658 15192
rect 15714 15136 16210 15192
rect 16266 15136 16271 15192
rect 15653 15134 16271 15136
rect 15653 15131 15719 15134
rect 16205 15131 16271 15134
rect 20713 15194 20779 15197
rect 23105 15194 23171 15197
rect 23657 15194 23723 15197
rect 20713 15192 23723 15194
rect 20713 15136 20718 15192
rect 20774 15136 23110 15192
rect 23166 15136 23662 15192
rect 23718 15136 23723 15192
rect 20713 15134 23723 15136
rect 20713 15131 20779 15134
rect 23105 15131 23171 15134
rect 23657 15131 23723 15134
rect 17585 15058 17651 15061
rect 7925 15056 10978 15058
rect 7925 15000 7930 15056
rect 7986 15000 8574 15056
rect 8630 15000 10978 15056
rect 7925 14998 10978 15000
rect 13356 15056 17651 15058
rect 13356 15000 17590 15056
rect 17646 15000 17651 15056
rect 13356 14998 17651 15000
rect 7925 14995 7991 14998
rect 8569 14995 8635 14998
rect 11329 14922 11395 14925
rect 11646 14922 11652 14924
rect 11329 14920 11652 14922
rect 11329 14864 11334 14920
rect 11390 14864 11652 14920
rect 11329 14862 11652 14864
rect 11329 14859 11395 14862
rect 11646 14860 11652 14862
rect 11716 14860 11722 14924
rect 8845 14786 8911 14789
rect 9070 14786 9076 14788
rect 8845 14784 9076 14786
rect 8845 14728 8850 14784
rect 8906 14728 9076 14784
rect 8845 14726 9076 14728
rect 8845 14723 8911 14726
rect 9070 14724 9076 14726
rect 9140 14724 9146 14788
rect 12157 14786 12223 14789
rect 13356 14786 13416 14998
rect 17585 14995 17651 14998
rect 19885 15058 19951 15061
rect 22185 15058 22251 15061
rect 19885 15056 22251 15058
rect 19885 15000 19890 15056
rect 19946 15000 22190 15056
rect 22246 15000 22251 15056
rect 19885 14998 22251 15000
rect 19885 14995 19951 14998
rect 22185 14995 22251 14998
rect 24526 14996 24532 15060
rect 24596 15058 24602 15060
rect 25129 15058 25195 15061
rect 24596 15056 25195 15058
rect 24596 15000 25134 15056
rect 25190 15000 25195 15056
rect 24596 14998 25195 15000
rect 24596 14996 24602 14998
rect 25129 14995 25195 14998
rect 13537 14922 13603 14925
rect 15469 14922 15535 14925
rect 13537 14920 15535 14922
rect 13537 14864 13542 14920
rect 13598 14864 15474 14920
rect 15530 14864 15535 14920
rect 13537 14862 15535 14864
rect 13537 14859 13603 14862
rect 15469 14859 15535 14862
rect 17350 14860 17356 14924
rect 17420 14922 17426 14924
rect 23473 14922 23539 14925
rect 17420 14920 23539 14922
rect 17420 14864 23478 14920
rect 23534 14864 23539 14920
rect 17420 14862 23539 14864
rect 17420 14860 17426 14862
rect 23473 14859 23539 14862
rect 12157 14784 13416 14786
rect 12157 14728 12162 14784
rect 12218 14728 13416 14784
rect 12157 14726 13416 14728
rect 12157 14723 12223 14726
rect 5436 14720 5756 14721
rect 5436 14656 5444 14720
rect 5508 14656 5524 14720
rect 5588 14656 5604 14720
rect 5668 14656 5684 14720
rect 5748 14656 5756 14720
rect 5436 14655 5756 14656
rect 14422 14720 14742 14721
rect 14422 14656 14430 14720
rect 14494 14656 14510 14720
rect 14574 14656 14590 14720
rect 14654 14656 14670 14720
rect 14734 14656 14742 14720
rect 14422 14655 14742 14656
rect 23407 14720 23727 14721
rect 23407 14656 23415 14720
rect 23479 14656 23495 14720
rect 23559 14656 23575 14720
rect 23639 14656 23655 14720
rect 23719 14656 23727 14720
rect 23407 14655 23727 14656
rect 9857 14650 9923 14653
rect 11881 14650 11947 14653
rect 9857 14648 11947 14650
rect 9857 14592 9862 14648
rect 9918 14592 11886 14648
rect 11942 14592 11947 14648
rect 9857 14590 11947 14592
rect 9857 14587 9923 14590
rect 11881 14587 11947 14590
rect 15878 14588 15884 14652
rect 15948 14650 15954 14652
rect 16573 14650 16639 14653
rect 15948 14648 16639 14650
rect 15948 14592 16578 14648
rect 16634 14592 16639 14648
rect 15948 14590 16639 14592
rect 15948 14588 15954 14590
rect 16573 14587 16639 14590
rect 19885 14650 19951 14653
rect 22645 14650 22711 14653
rect 23197 14650 23263 14653
rect 19885 14648 21788 14650
rect 19885 14592 19890 14648
rect 19946 14592 21788 14648
rect 19885 14590 21788 14592
rect 19885 14587 19951 14590
rect 12709 14514 12775 14517
rect 16665 14514 16731 14517
rect 12709 14512 16731 14514
rect 12709 14456 12714 14512
rect 12770 14456 16670 14512
rect 16726 14456 16731 14512
rect 12709 14454 16731 14456
rect 12709 14451 12775 14454
rect 16665 14451 16731 14454
rect 20529 14514 20595 14517
rect 21541 14514 21607 14517
rect 20529 14512 21607 14514
rect 20529 14456 20534 14512
rect 20590 14456 21546 14512
rect 21602 14456 21607 14512
rect 20529 14454 21607 14456
rect 21728 14514 21788 14590
rect 22645 14648 23263 14650
rect 22645 14592 22650 14648
rect 22706 14592 23202 14648
rect 23258 14592 23263 14648
rect 22645 14590 23263 14592
rect 22645 14587 22711 14590
rect 23197 14587 23263 14590
rect 23657 14514 23723 14517
rect 24158 14514 24164 14516
rect 21728 14512 24164 14514
rect 21728 14456 23662 14512
rect 23718 14456 24164 14512
rect 21728 14454 24164 14456
rect 20529 14451 20595 14454
rect 21541 14451 21607 14454
rect 23657 14451 23723 14454
rect 24158 14452 24164 14454
rect 24228 14514 24234 14516
rect 26509 14514 26575 14517
rect 24228 14512 26575 14514
rect 24228 14456 26514 14512
rect 26570 14456 26575 14512
rect 24228 14454 26575 14456
rect 24228 14452 24234 14454
rect 26509 14451 26575 14454
rect 3877 14380 3943 14381
rect 3877 14376 3924 14380
rect 3988 14378 3994 14380
rect 10685 14378 10751 14381
rect 13486 14378 13492 14380
rect 3877 14320 3882 14376
rect 3877 14316 3924 14320
rect 3988 14318 4034 14378
rect 10685 14376 13492 14378
rect 10685 14320 10690 14376
rect 10746 14320 13492 14376
rect 10685 14318 13492 14320
rect 3988 14316 3994 14318
rect 3877 14315 3943 14316
rect 10685 14315 10751 14318
rect 13486 14316 13492 14318
rect 13556 14316 13562 14380
rect 13721 14378 13787 14381
rect 18505 14378 18571 14381
rect 13721 14376 18571 14378
rect 13721 14320 13726 14376
rect 13782 14320 18510 14376
rect 18566 14320 18571 14376
rect 13721 14318 18571 14320
rect 13721 14315 13787 14318
rect 18505 14315 18571 14318
rect 18638 14316 18644 14380
rect 18708 14378 18714 14380
rect 20662 14378 20668 14380
rect 18708 14318 20668 14378
rect 18708 14316 18714 14318
rect 20662 14316 20668 14318
rect 20732 14378 20738 14380
rect 22093 14378 22159 14381
rect 22645 14378 22711 14381
rect 20732 14318 21880 14378
rect 20732 14316 20738 14318
rect 3141 14242 3207 14245
rect 3141 14240 3250 14242
rect 3141 14184 3146 14240
rect 3202 14184 3250 14240
rect 3141 14179 3250 14184
rect 11278 14180 11284 14244
rect 11348 14242 11354 14244
rect 11513 14242 11579 14245
rect 11348 14240 11579 14242
rect 11348 14184 11518 14240
rect 11574 14184 11579 14240
rect 11348 14182 11579 14184
rect 11348 14180 11354 14182
rect 11513 14179 11579 14182
rect 15009 14242 15075 14245
rect 16246 14242 16252 14244
rect 15009 14240 16252 14242
rect 15009 14184 15014 14240
rect 15070 14184 16252 14240
rect 15009 14182 16252 14184
rect 15009 14179 15075 14182
rect 16246 14180 16252 14182
rect 16316 14180 16322 14244
rect 21449 14242 21515 14245
rect 21406 14240 21515 14242
rect 21406 14184 21454 14240
rect 21510 14184 21515 14240
rect 21406 14179 21515 14184
rect 21820 14242 21880 14318
rect 22093 14376 22711 14378
rect 22093 14320 22098 14376
rect 22154 14320 22650 14376
rect 22706 14320 22711 14376
rect 22093 14318 22711 14320
rect 22093 14315 22159 14318
rect 22645 14315 22711 14318
rect 23105 14378 23171 14381
rect 25313 14378 25379 14381
rect 23105 14376 25379 14378
rect 23105 14320 23110 14376
rect 23166 14320 25318 14376
rect 25374 14320 25379 14376
rect 23105 14318 25379 14320
rect 23105 14315 23171 14318
rect 25313 14315 25379 14318
rect 22185 14242 22251 14245
rect 21820 14240 22251 14242
rect 21820 14184 22190 14240
rect 22246 14184 22251 14240
rect 21820 14182 22251 14184
rect 22185 14179 22251 14182
rect 3190 13834 3250 14179
rect 9929 14176 10249 14177
rect 9929 14112 9937 14176
rect 10001 14112 10017 14176
rect 10081 14112 10097 14176
rect 10161 14112 10177 14176
rect 10241 14112 10249 14176
rect 9929 14111 10249 14112
rect 18914 14176 19234 14177
rect 18914 14112 18922 14176
rect 18986 14112 19002 14176
rect 19066 14112 19082 14176
rect 19146 14112 19162 14176
rect 19226 14112 19234 14176
rect 18914 14111 19234 14112
rect 10869 14106 10935 14109
rect 14641 14106 14707 14109
rect 10869 14104 14707 14106
rect 10869 14048 10874 14104
rect 10930 14048 14646 14104
rect 14702 14048 14707 14104
rect 10869 14046 14707 14048
rect 10869 14043 10935 14046
rect 14641 14043 14707 14046
rect 21406 13973 21466 14179
rect 3550 13908 3556 13972
rect 3620 13970 3626 13972
rect 6821 13970 6887 13973
rect 3620 13968 6887 13970
rect 3620 13912 6826 13968
rect 6882 13912 6887 13968
rect 3620 13910 6887 13912
rect 3620 13908 3626 13910
rect 6821 13907 6887 13910
rect 11513 13970 11579 13973
rect 11646 13970 11652 13972
rect 11513 13968 11652 13970
rect 11513 13912 11518 13968
rect 11574 13912 11652 13968
rect 11513 13910 11652 13912
rect 11513 13907 11579 13910
rect 11646 13908 11652 13910
rect 11716 13908 11722 13972
rect 13169 13970 13235 13973
rect 15009 13970 15075 13973
rect 13169 13968 15075 13970
rect 13169 13912 13174 13968
rect 13230 13912 15014 13968
rect 15070 13912 15075 13968
rect 13169 13910 15075 13912
rect 13169 13907 13235 13910
rect 15009 13907 15075 13910
rect 15469 13972 15535 13973
rect 15469 13968 15516 13972
rect 15580 13970 15586 13972
rect 18413 13970 18479 13973
rect 19149 13970 19215 13973
rect 15469 13912 15474 13968
rect 15469 13908 15516 13912
rect 15580 13910 15626 13970
rect 18413 13968 19215 13970
rect 18413 13912 18418 13968
rect 18474 13912 19154 13968
rect 19210 13912 19215 13968
rect 18413 13910 19215 13912
rect 15580 13908 15586 13910
rect 15469 13907 15535 13908
rect 18413 13907 18479 13910
rect 19149 13907 19215 13910
rect 19517 13970 19583 13973
rect 19517 13968 21282 13970
rect 19517 13912 19522 13968
rect 19578 13912 21282 13968
rect 19517 13910 21282 13912
rect 21406 13968 21515 13973
rect 21406 13912 21454 13968
rect 21510 13912 21515 13968
rect 21406 13910 21515 13912
rect 19517 13907 19583 13910
rect 3877 13834 3943 13837
rect 3190 13832 3943 13834
rect 3190 13776 3882 13832
rect 3938 13776 3943 13832
rect 3190 13774 3943 13776
rect 3877 13771 3943 13774
rect 15837 13834 15903 13837
rect 16062 13834 16068 13836
rect 15837 13832 16068 13834
rect 15837 13776 15842 13832
rect 15898 13776 16068 13832
rect 15837 13774 16068 13776
rect 15837 13771 15903 13774
rect 16062 13772 16068 13774
rect 16132 13772 16138 13836
rect 17718 13772 17724 13836
rect 17788 13834 17794 13836
rect 19885 13834 19951 13837
rect 17788 13832 19951 13834
rect 17788 13776 19890 13832
rect 19946 13776 19951 13832
rect 17788 13774 19951 13776
rect 21222 13834 21282 13910
rect 21449 13907 21515 13910
rect 21725 13970 21791 13973
rect 22001 13970 22067 13973
rect 21725 13968 22067 13970
rect 21725 13912 21730 13968
rect 21786 13912 22006 13968
rect 22062 13912 22067 13968
rect 21725 13910 22067 13912
rect 21725 13907 21791 13910
rect 22001 13907 22067 13910
rect 23473 13970 23539 13973
rect 24209 13970 24275 13973
rect 23473 13968 24275 13970
rect 23473 13912 23478 13968
rect 23534 13912 24214 13968
rect 24270 13912 24275 13968
rect 23473 13910 24275 13912
rect 23473 13907 23539 13910
rect 24209 13907 24275 13910
rect 22277 13834 22343 13837
rect 21222 13832 22343 13834
rect 21222 13776 22282 13832
rect 22338 13776 22343 13832
rect 21222 13774 22343 13776
rect 17788 13772 17794 13774
rect 19885 13771 19951 13774
rect 22277 13771 22343 13774
rect 22645 13834 22711 13837
rect 25221 13834 25287 13837
rect 22645 13832 25287 13834
rect 22645 13776 22650 13832
rect 22706 13776 25226 13832
rect 25282 13776 25287 13832
rect 22645 13774 25287 13776
rect 22645 13771 22711 13774
rect 25221 13771 25287 13774
rect 2957 13698 3023 13701
rect 17585 13700 17651 13701
rect 4102 13698 4108 13700
rect 2957 13696 4108 13698
rect 2957 13640 2962 13696
rect 3018 13640 4108 13696
rect 2957 13638 4108 13640
rect 2957 13635 3023 13638
rect 4102 13636 4108 13638
rect 4172 13636 4178 13700
rect 17534 13698 17540 13700
rect 17494 13638 17540 13698
rect 17604 13696 17651 13700
rect 17646 13640 17651 13696
rect 17534 13636 17540 13638
rect 17604 13636 17651 13640
rect 19888 13698 19948 13771
rect 21541 13698 21607 13701
rect 19888 13696 21607 13698
rect 19888 13640 21546 13696
rect 21602 13640 21607 13696
rect 19888 13638 21607 13640
rect 17585 13635 17651 13636
rect 21541 13635 21607 13638
rect 5436 13632 5756 13633
rect 5436 13568 5444 13632
rect 5508 13568 5524 13632
rect 5588 13568 5604 13632
rect 5668 13568 5684 13632
rect 5748 13568 5756 13632
rect 5436 13567 5756 13568
rect 14422 13632 14742 13633
rect 14422 13568 14430 13632
rect 14494 13568 14510 13632
rect 14574 13568 14590 13632
rect 14654 13568 14670 13632
rect 14734 13568 14742 13632
rect 14422 13567 14742 13568
rect 23407 13632 23727 13633
rect 23407 13568 23415 13632
rect 23479 13568 23495 13632
rect 23559 13568 23575 13632
rect 23639 13568 23655 13632
rect 23719 13568 23727 13632
rect 23407 13567 23727 13568
rect 3233 13564 3299 13565
rect 3182 13500 3188 13564
rect 3252 13562 3299 13564
rect 19149 13562 19215 13565
rect 3252 13560 3344 13562
rect 3294 13504 3344 13560
rect 3252 13502 3344 13504
rect 16990 13560 19215 13562
rect 16990 13504 19154 13560
rect 19210 13504 19215 13560
rect 16990 13502 19215 13504
rect 3252 13500 3299 13502
rect 3233 13499 3299 13500
rect 13261 13426 13327 13429
rect 16990 13426 17050 13502
rect 19149 13499 19215 13502
rect 13261 13424 17050 13426
rect 13261 13368 13266 13424
rect 13322 13368 17050 13424
rect 13261 13366 17050 13368
rect 17125 13426 17191 13429
rect 17902 13426 17908 13428
rect 17125 13424 17908 13426
rect 17125 13368 17130 13424
rect 17186 13368 17908 13424
rect 17125 13366 17908 13368
rect 13261 13363 13327 13366
rect 17125 13363 17191 13366
rect 17902 13364 17908 13366
rect 17972 13364 17978 13428
rect 20529 13426 20595 13429
rect 26417 13426 26483 13429
rect 20529 13424 26483 13426
rect 20529 13368 20534 13424
rect 20590 13368 26422 13424
rect 26478 13368 26483 13424
rect 20529 13366 26483 13368
rect 20529 13363 20595 13366
rect 26417 13363 26483 13366
rect 4889 13290 4955 13293
rect 5165 13292 5231 13293
rect 5165 13290 5212 13292
rect 4294 13288 4955 13290
rect 4294 13232 4894 13288
rect 4950 13232 4955 13288
rect 4294 13230 4955 13232
rect 5120 13288 5212 13290
rect 5120 13232 5170 13288
rect 5120 13230 5212 13232
rect 3601 13020 3667 13021
rect 3550 12956 3556 13020
rect 3620 13018 3667 13020
rect 3620 13016 3712 13018
rect 3662 12960 3712 13016
rect 3620 12958 3712 12960
rect 3620 12956 3667 12958
rect 3601 12955 3667 12956
rect 3182 12820 3188 12884
rect 3252 12882 3258 12884
rect 3417 12882 3483 12885
rect 3252 12880 3483 12882
rect 3252 12824 3422 12880
rect 3478 12824 3483 12880
rect 3252 12822 3483 12824
rect 3252 12820 3258 12822
rect 3417 12819 3483 12822
rect 2681 12744 2747 12749
rect 2681 12688 2686 12744
rect 2742 12688 2747 12744
rect 2681 12683 2747 12688
rect 2684 12202 2744 12683
rect 4294 12610 4354 13230
rect 4889 13227 4955 13230
rect 5165 13228 5212 13230
rect 5276 13228 5282 13292
rect 7925 13290 7991 13293
rect 8702 13290 8708 13292
rect 7925 13288 8708 13290
rect 7925 13232 7930 13288
rect 7986 13232 8708 13288
rect 7925 13230 8708 13232
rect 5165 13227 5231 13228
rect 7925 13227 7991 13230
rect 8702 13228 8708 13230
rect 8772 13228 8778 13292
rect 18045 13288 18111 13293
rect 18045 13232 18050 13288
rect 18106 13232 18111 13288
rect 18045 13227 18111 13232
rect 22093 13290 22159 13293
rect 24025 13290 24091 13293
rect 22093 13288 24091 13290
rect 22093 13232 22098 13288
rect 22154 13232 24030 13288
rect 24086 13232 24091 13288
rect 22093 13230 24091 13232
rect 22093 13227 22159 13230
rect 24025 13227 24091 13230
rect 9121 13154 9187 13157
rect 9438 13154 9444 13156
rect 9121 13152 9444 13154
rect 9121 13096 9126 13152
rect 9182 13096 9444 13152
rect 9121 13094 9444 13096
rect 9121 13091 9187 13094
rect 9438 13092 9444 13094
rect 9508 13092 9514 13156
rect 17769 13154 17835 13157
rect 18048 13154 18108 13227
rect 18505 13156 18571 13157
rect 17769 13152 18108 13154
rect 17769 13096 17774 13152
rect 17830 13096 18108 13152
rect 17769 13094 18108 13096
rect 17769 13091 17835 13094
rect 18454 13092 18460 13156
rect 18524 13154 18571 13156
rect 19517 13154 19583 13157
rect 20621 13154 20687 13157
rect 18524 13152 18616 13154
rect 18566 13096 18616 13152
rect 18524 13094 18616 13096
rect 19517 13152 20687 13154
rect 19517 13096 19522 13152
rect 19578 13096 20626 13152
rect 20682 13096 20687 13152
rect 19517 13094 20687 13096
rect 18524 13092 18571 13094
rect 18505 13091 18571 13092
rect 19517 13091 19583 13094
rect 20621 13091 20687 13094
rect 23238 13092 23244 13156
rect 23308 13154 23314 13156
rect 23381 13154 23447 13157
rect 23308 13152 23447 13154
rect 23308 13096 23386 13152
rect 23442 13096 23447 13152
rect 23308 13094 23447 13096
rect 23308 13092 23314 13094
rect 23381 13091 23447 13094
rect 9929 13088 10249 13089
rect 9929 13024 9937 13088
rect 10001 13024 10017 13088
rect 10081 13024 10097 13088
rect 10161 13024 10177 13088
rect 10241 13024 10249 13088
rect 9929 13023 10249 13024
rect 18914 13088 19234 13089
rect 18914 13024 18922 13088
rect 18986 13024 19002 13088
rect 19066 13024 19082 13088
rect 19146 13024 19162 13088
rect 19226 13024 19234 13088
rect 18914 13023 19234 13024
rect 4654 12956 4660 13020
rect 4724 13018 4730 13020
rect 9213 13018 9279 13021
rect 4724 13016 9279 13018
rect 4724 12960 9218 13016
rect 9274 12960 9279 13016
rect 4724 12958 9279 12960
rect 4724 12956 4730 12958
rect 9213 12955 9279 12958
rect 15142 12956 15148 13020
rect 15212 13018 15218 13020
rect 15469 13018 15535 13021
rect 15212 13016 15535 13018
rect 15212 12960 15474 13016
rect 15530 12960 15535 13016
rect 15212 12958 15535 12960
rect 15212 12956 15218 12958
rect 15469 12955 15535 12958
rect 17953 13018 18019 13021
rect 18321 13018 18387 13021
rect 17953 13016 18387 13018
rect 17953 12960 17958 13016
rect 18014 12960 18326 13016
rect 18382 12960 18387 13016
rect 17953 12958 18387 12960
rect 17953 12955 18019 12958
rect 18321 12955 18387 12958
rect 18505 13018 18571 13021
rect 18689 13018 18755 13021
rect 18505 13016 18755 13018
rect 18505 12960 18510 13016
rect 18566 12960 18694 13016
rect 18750 12960 18755 13016
rect 18505 12958 18755 12960
rect 18505 12955 18571 12958
rect 18689 12955 18755 12958
rect 20989 13018 21055 13021
rect 20989 13016 21098 13018
rect 20989 12960 20994 13016
rect 21050 12960 21098 13016
rect 20989 12955 21098 12960
rect 4654 12820 4660 12884
rect 4724 12882 4730 12884
rect 5533 12882 5599 12885
rect 8569 12884 8635 12885
rect 8518 12882 8524 12884
rect 4724 12880 5599 12882
rect 4724 12824 5538 12880
rect 5594 12824 5599 12880
rect 4724 12822 5599 12824
rect 8478 12822 8524 12882
rect 8588 12880 8635 12884
rect 8630 12824 8635 12880
rect 4724 12820 4730 12822
rect 5533 12819 5599 12822
rect 8518 12820 8524 12822
rect 8588 12820 8635 12824
rect 8569 12819 8635 12820
rect 13997 12882 14063 12885
rect 14958 12882 14964 12884
rect 13997 12880 14964 12882
rect 13997 12824 14002 12880
rect 14058 12824 14964 12880
rect 13997 12822 14964 12824
rect 13997 12819 14063 12822
rect 14958 12820 14964 12822
rect 15028 12820 15034 12884
rect 15837 12882 15903 12885
rect 17861 12882 17927 12885
rect 15837 12880 17927 12882
rect 15837 12824 15842 12880
rect 15898 12824 17866 12880
rect 17922 12824 17927 12880
rect 15837 12822 17927 12824
rect 15837 12819 15903 12822
rect 17861 12819 17927 12822
rect 7833 12748 7899 12749
rect 4470 12684 4476 12748
rect 4540 12746 4546 12748
rect 7782 12746 7788 12748
rect 4540 12686 5044 12746
rect 7742 12686 7788 12746
rect 7852 12744 7899 12748
rect 7894 12688 7899 12744
rect 4540 12684 4546 12686
rect 4470 12610 4476 12612
rect 4294 12550 4476 12610
rect 4470 12548 4476 12550
rect 4540 12548 4546 12612
rect 2998 12412 3004 12476
rect 3068 12474 3074 12476
rect 4153 12474 4219 12477
rect 3068 12472 4219 12474
rect 3068 12416 4158 12472
rect 4214 12416 4219 12472
rect 3068 12414 4219 12416
rect 3068 12412 3074 12414
rect 4153 12411 4219 12414
rect 4705 12474 4771 12477
rect 4838 12474 4844 12476
rect 4705 12472 4844 12474
rect 4705 12416 4710 12472
rect 4766 12416 4844 12472
rect 4705 12414 4844 12416
rect 4705 12411 4771 12414
rect 4838 12412 4844 12414
rect 4908 12412 4914 12476
rect 4984 12474 5044 12686
rect 7782 12684 7788 12686
rect 7852 12684 7899 12688
rect 7966 12684 7972 12748
rect 8036 12746 8042 12748
rect 10409 12746 10475 12749
rect 8036 12744 10475 12746
rect 8036 12688 10414 12744
rect 10470 12688 10475 12744
rect 8036 12686 10475 12688
rect 8036 12684 8042 12686
rect 7833 12683 7899 12684
rect 10409 12683 10475 12686
rect 5257 12612 5323 12613
rect 6545 12612 6611 12613
rect 5206 12610 5212 12612
rect 5166 12550 5212 12610
rect 5276 12608 5323 12612
rect 5318 12552 5323 12608
rect 5206 12548 5212 12550
rect 5276 12548 5323 12552
rect 6494 12548 6500 12612
rect 6564 12610 6611 12612
rect 7373 12610 7439 12613
rect 6564 12608 6656 12610
rect 6606 12552 6656 12608
rect 6564 12550 6656 12552
rect 7373 12608 7712 12610
rect 7373 12552 7378 12608
rect 7434 12552 7712 12608
rect 7373 12550 7712 12552
rect 6564 12548 6611 12550
rect 5257 12547 5323 12548
rect 6545 12547 6611 12548
rect 7373 12547 7439 12550
rect 5436 12544 5756 12545
rect 5436 12480 5444 12544
rect 5508 12480 5524 12544
rect 5588 12480 5604 12544
rect 5668 12480 5684 12544
rect 5748 12480 5756 12544
rect 5436 12479 5756 12480
rect 7652 12477 7712 12550
rect 8702 12548 8708 12612
rect 8772 12610 8778 12612
rect 8845 12610 8911 12613
rect 9397 12610 9463 12613
rect 8772 12608 8911 12610
rect 8772 12552 8850 12608
rect 8906 12552 8911 12608
rect 8772 12550 8911 12552
rect 8772 12548 8778 12550
rect 8845 12547 8911 12550
rect 9078 12608 9463 12610
rect 9078 12552 9402 12608
rect 9458 12552 9463 12608
rect 9078 12550 9463 12552
rect 5257 12474 5323 12477
rect 4984 12472 5323 12474
rect 4984 12416 5262 12472
rect 5318 12416 5323 12472
rect 4984 12414 5323 12416
rect 5257 12411 5323 12414
rect 7005 12476 7071 12477
rect 7005 12472 7052 12476
rect 7116 12474 7122 12476
rect 7005 12416 7010 12472
rect 7005 12412 7052 12416
rect 7116 12414 7162 12474
rect 7116 12412 7122 12414
rect 7230 12412 7236 12476
rect 7300 12474 7306 12476
rect 7373 12474 7439 12477
rect 7300 12472 7439 12474
rect 7300 12416 7378 12472
rect 7434 12416 7439 12472
rect 7300 12414 7439 12416
rect 7300 12412 7306 12414
rect 7005 12411 7071 12412
rect 7373 12411 7439 12414
rect 7649 12472 7715 12477
rect 7649 12416 7654 12472
rect 7710 12416 7715 12472
rect 7649 12411 7715 12416
rect 8661 12474 8727 12477
rect 9078 12474 9138 12550
rect 9397 12547 9463 12550
rect 14422 12544 14742 12545
rect 14422 12480 14430 12544
rect 14494 12480 14510 12544
rect 14574 12480 14590 12544
rect 14654 12480 14670 12544
rect 14734 12480 14742 12544
rect 14422 12479 14742 12480
rect 8661 12472 9138 12474
rect 8661 12416 8666 12472
rect 8722 12416 9138 12472
rect 8661 12414 9138 12416
rect 8661 12411 8727 12414
rect 9254 12412 9260 12476
rect 9324 12474 9330 12476
rect 9397 12474 9463 12477
rect 9324 12472 9463 12474
rect 9324 12416 9402 12472
rect 9458 12416 9463 12472
rect 9324 12414 9463 12416
rect 9324 12412 9330 12414
rect 9397 12411 9463 12414
rect 13077 12474 13143 12477
rect 13721 12474 13787 12477
rect 13077 12472 13787 12474
rect 13077 12416 13082 12472
rect 13138 12416 13726 12472
rect 13782 12416 13787 12472
rect 13077 12414 13787 12416
rect 21038 12474 21098 12955
rect 26601 12882 26667 12885
rect 26558 12880 26667 12882
rect 26558 12824 26606 12880
rect 26662 12824 26667 12880
rect 26558 12819 26667 12824
rect 22870 12684 22876 12748
rect 22940 12746 22946 12748
rect 24117 12746 24183 12749
rect 22940 12744 24183 12746
rect 22940 12688 24122 12744
rect 24178 12688 24183 12744
rect 22940 12686 24183 12688
rect 22940 12684 22946 12686
rect 24117 12683 24183 12686
rect 26141 12746 26207 12749
rect 26558 12746 26618 12819
rect 26141 12744 26618 12746
rect 26141 12688 26146 12744
rect 26202 12688 26618 12744
rect 26141 12686 26618 12688
rect 27061 12746 27127 12749
rect 27061 12744 27584 12746
rect 27061 12688 27066 12744
rect 27122 12688 27584 12744
rect 27061 12686 27584 12688
rect 26141 12683 26207 12686
rect 27061 12683 27127 12686
rect 21265 12610 21331 12613
rect 21398 12610 21404 12612
rect 21265 12608 21404 12610
rect 21265 12552 21270 12608
rect 21326 12552 21404 12608
rect 21265 12550 21404 12552
rect 21265 12547 21331 12550
rect 21398 12548 21404 12550
rect 21468 12548 21474 12612
rect 23407 12544 23727 12545
rect 23407 12480 23415 12544
rect 23479 12480 23495 12544
rect 23559 12480 23575 12544
rect 23639 12480 23655 12544
rect 23719 12480 23727 12544
rect 23407 12479 23727 12480
rect 27524 12477 27584 12686
rect 21265 12474 21331 12477
rect 24117 12476 24183 12477
rect 24117 12474 24164 12476
rect 21038 12472 21331 12474
rect 21038 12416 21270 12472
rect 21326 12416 21331 12472
rect 21038 12414 21331 12416
rect 24072 12472 24164 12474
rect 24072 12416 24122 12472
rect 24072 12414 24164 12416
rect 13077 12411 13143 12414
rect 13721 12411 13787 12414
rect 21265 12411 21331 12414
rect 24117 12412 24164 12414
rect 24228 12412 24234 12476
rect 27521 12472 27587 12477
rect 27521 12416 27526 12472
rect 27582 12416 27587 12472
rect 24117 12411 24183 12412
rect 27521 12411 27587 12416
rect 4521 12340 4587 12341
rect 6545 12340 6611 12341
rect 4470 12338 4476 12340
rect 4430 12278 4476 12338
rect 4540 12336 4587 12340
rect 6494 12338 6500 12340
rect 4582 12280 4587 12336
rect 4470 12276 4476 12278
rect 4540 12276 4587 12280
rect 6454 12278 6500 12338
rect 6564 12336 6611 12340
rect 6606 12280 6611 12336
rect 6494 12276 6500 12278
rect 6564 12276 6611 12280
rect 4521 12275 4587 12276
rect 6545 12275 6611 12276
rect 6729 12338 6795 12341
rect 6862 12338 6868 12340
rect 6729 12336 6868 12338
rect 6729 12280 6734 12336
rect 6790 12280 6868 12336
rect 6729 12278 6868 12280
rect 6729 12275 6795 12278
rect 6862 12276 6868 12278
rect 6932 12276 6938 12340
rect 7046 12276 7052 12340
rect 7116 12338 7122 12340
rect 7189 12338 7255 12341
rect 7373 12340 7439 12341
rect 7741 12340 7807 12341
rect 7373 12338 7420 12340
rect 7116 12336 7255 12338
rect 7116 12280 7194 12336
rect 7250 12280 7255 12336
rect 7116 12278 7255 12280
rect 7328 12336 7420 12338
rect 7328 12280 7378 12336
rect 7328 12278 7420 12280
rect 7116 12276 7122 12278
rect 7189 12275 7255 12278
rect 7373 12276 7420 12278
rect 7484 12276 7490 12340
rect 7741 12336 7788 12340
rect 7852 12338 7858 12340
rect 7741 12280 7746 12336
rect 7741 12276 7788 12280
rect 7852 12278 7898 12338
rect 7852 12276 7858 12278
rect 8518 12276 8524 12340
rect 8588 12338 8594 12340
rect 8661 12338 8727 12341
rect 8588 12336 8727 12338
rect 8588 12280 8666 12336
rect 8722 12280 8727 12336
rect 8588 12278 8727 12280
rect 8588 12276 8594 12278
rect 7373 12275 7439 12276
rect 7741 12275 7807 12276
rect 8661 12275 8727 12278
rect 9581 12338 9647 12341
rect 10869 12340 10935 12341
rect 9581 12336 10196 12338
rect 9581 12280 9586 12336
rect 9642 12280 10196 12336
rect 9581 12278 10196 12280
rect 9581 12275 9647 12278
rect 10136 12202 10196 12278
rect 10869 12336 10916 12340
rect 10980 12338 10986 12340
rect 15929 12338 15995 12341
rect 16430 12338 16436 12340
rect 10869 12280 10874 12336
rect 10869 12276 10916 12280
rect 10980 12278 11026 12338
rect 15929 12336 16436 12338
rect 15929 12280 15934 12336
rect 15990 12280 16436 12336
rect 15929 12278 16436 12280
rect 10980 12276 10986 12278
rect 10869 12275 10935 12276
rect 15929 12275 15995 12278
rect 16430 12276 16436 12278
rect 16500 12276 16506 12340
rect 17585 12338 17651 12341
rect 19701 12338 19767 12341
rect 25865 12338 25931 12341
rect 17585 12336 17970 12338
rect 17585 12280 17590 12336
rect 17646 12280 17970 12336
rect 17585 12278 17970 12280
rect 17585 12275 17651 12278
rect 10593 12202 10659 12205
rect 10777 12204 10843 12205
rect 2684 12142 8218 12202
rect 10136 12200 10659 12202
rect 10136 12144 10598 12200
rect 10654 12144 10659 12200
rect 10136 12142 10659 12144
rect 8158 12069 8218 12142
rect 10593 12139 10659 12142
rect 10726 12140 10732 12204
rect 10796 12202 10843 12204
rect 16941 12202 17007 12205
rect 17910 12204 17970 12278
rect 19701 12336 25931 12338
rect 19701 12280 19706 12336
rect 19762 12280 25870 12336
rect 25926 12280 25931 12336
rect 19701 12278 25931 12280
rect 19701 12275 19767 12278
rect 25865 12275 25931 12278
rect 17350 12202 17356 12204
rect 10796 12200 10888 12202
rect 10838 12144 10888 12200
rect 10796 12142 10888 12144
rect 16941 12200 17356 12202
rect 16941 12144 16946 12200
rect 17002 12144 17356 12200
rect 16941 12142 17356 12144
rect 10796 12140 10843 12142
rect 10777 12139 10843 12140
rect 16941 12139 17007 12142
rect 17350 12140 17356 12142
rect 17420 12140 17426 12204
rect 17902 12140 17908 12204
rect 17972 12140 17978 12204
rect 18965 12202 19031 12205
rect 18692 12200 19031 12202
rect 18692 12144 18970 12200
rect 19026 12144 19031 12200
rect 18692 12142 19031 12144
rect 2957 12068 3023 12069
rect 2957 12064 3004 12068
rect 3068 12066 3074 12068
rect 4061 12066 4127 12069
rect 4705 12068 4771 12069
rect 4286 12066 4292 12068
rect 2957 12008 2962 12064
rect 2957 12004 3004 12008
rect 3068 12006 3114 12066
rect 4061 12064 4292 12066
rect 4061 12008 4066 12064
rect 4122 12008 4292 12064
rect 4061 12006 4292 12008
rect 3068 12004 3074 12006
rect 2957 12003 3023 12004
rect 4061 12003 4127 12006
rect 4286 12004 4292 12006
rect 4356 12004 4362 12068
rect 4654 12066 4660 12068
rect 4614 12006 4660 12066
rect 4724 12064 4771 12068
rect 4766 12008 4771 12064
rect 4654 12004 4660 12006
rect 4724 12004 4771 12008
rect 6678 12004 6684 12068
rect 6748 12066 6754 12068
rect 6821 12066 6887 12069
rect 6748 12064 6887 12066
rect 6748 12008 6826 12064
rect 6882 12008 6887 12064
rect 6748 12006 6887 12008
rect 6748 12004 6754 12006
rect 4705 12003 4771 12004
rect 6821 12003 6887 12006
rect 7189 12066 7255 12069
rect 7598 12066 7604 12068
rect 7189 12064 7604 12066
rect 7189 12008 7194 12064
rect 7250 12008 7604 12064
rect 7189 12006 7604 12008
rect 7189 12003 7255 12006
rect 7598 12004 7604 12006
rect 7668 12004 7674 12068
rect 8158 12064 8267 12069
rect 8158 12008 8206 12064
rect 8262 12008 8267 12064
rect 8158 12006 8267 12008
rect 8201 12003 8267 12006
rect 14038 12004 14044 12068
rect 14108 12066 14114 12068
rect 14181 12066 14247 12069
rect 14108 12064 14247 12066
rect 14108 12008 14186 12064
rect 14242 12008 14247 12064
rect 14108 12006 14247 12008
rect 14108 12004 14114 12006
rect 14181 12003 14247 12006
rect 17350 12004 17356 12068
rect 17420 12066 17426 12068
rect 17585 12066 17651 12069
rect 17420 12064 17651 12066
rect 17420 12008 17590 12064
rect 17646 12008 17651 12064
rect 17420 12006 17651 12008
rect 17420 12004 17426 12006
rect 17585 12003 17651 12006
rect 9929 12000 10249 12001
rect 9929 11936 9937 12000
rect 10001 11936 10017 12000
rect 10081 11936 10097 12000
rect 10161 11936 10177 12000
rect 10241 11936 10249 12000
rect 9929 11935 10249 11936
rect 5942 11868 5948 11932
rect 6012 11930 6018 11932
rect 6361 11930 6427 11933
rect 6012 11928 6427 11930
rect 6012 11872 6366 11928
rect 6422 11872 6427 11928
rect 6012 11870 6427 11872
rect 6012 11868 6018 11870
rect 6361 11867 6427 11870
rect 14641 11930 14707 11933
rect 16982 11930 16988 11932
rect 14641 11928 16988 11930
rect 14641 11872 14646 11928
rect 14702 11872 16988 11928
rect 14641 11870 16988 11872
rect 14641 11867 14707 11870
rect 16982 11868 16988 11870
rect 17052 11868 17058 11932
rect 17585 11930 17651 11933
rect 18270 11930 18276 11932
rect 17585 11928 18276 11930
rect 17585 11872 17590 11928
rect 17646 11872 18276 11928
rect 17585 11870 18276 11872
rect 17585 11867 17651 11870
rect 18270 11868 18276 11870
rect 18340 11868 18346 11932
rect 9438 11732 9444 11796
rect 9508 11794 9514 11796
rect 9581 11794 9647 11797
rect 9508 11792 9647 11794
rect 9508 11736 9586 11792
rect 9642 11736 9647 11792
rect 9508 11734 9647 11736
rect 9508 11732 9514 11734
rect 9581 11731 9647 11734
rect 9765 11794 9831 11797
rect 12014 11794 12020 11796
rect 9765 11792 12020 11794
rect 9765 11736 9770 11792
rect 9826 11736 12020 11792
rect 9765 11734 12020 11736
rect 9765 11731 9831 11734
rect 12014 11732 12020 11734
rect 12084 11732 12090 11796
rect 17534 11732 17540 11796
rect 17604 11794 17610 11796
rect 17677 11794 17743 11797
rect 17604 11792 17743 11794
rect 17604 11736 17682 11792
rect 17738 11736 17743 11792
rect 17604 11734 17743 11736
rect 18692 11794 18752 12142
rect 18965 12139 19031 12142
rect 21398 12004 21404 12068
rect 21468 12066 21474 12068
rect 21725 12066 21791 12069
rect 21468 12064 21791 12066
rect 21468 12008 21730 12064
rect 21786 12008 21791 12064
rect 21468 12006 21791 12008
rect 21468 12004 21474 12006
rect 21725 12003 21791 12006
rect 18914 12000 19234 12001
rect 18914 11936 18922 12000
rect 18986 11936 19002 12000
rect 19066 11936 19082 12000
rect 19146 11936 19162 12000
rect 19226 11936 19234 12000
rect 18914 11935 19234 11936
rect 21173 11932 21239 11933
rect 21173 11928 21220 11932
rect 21284 11930 21290 11932
rect 21173 11872 21178 11928
rect 21173 11868 21220 11872
rect 21284 11870 21330 11930
rect 21284 11868 21290 11870
rect 21173 11867 21239 11868
rect 18873 11794 18939 11797
rect 18692 11792 18939 11794
rect 18692 11736 18878 11792
rect 18934 11736 18939 11792
rect 18692 11734 18939 11736
rect 17604 11732 17610 11734
rect 17677 11731 17743 11734
rect 18873 11731 18939 11734
rect 3918 11596 3924 11660
rect 3988 11658 3994 11660
rect 5073 11658 5139 11661
rect 3988 11656 5139 11658
rect 3988 11600 5078 11656
rect 5134 11600 5139 11656
rect 3988 11598 5139 11600
rect 3988 11596 3994 11598
rect 5073 11595 5139 11598
rect 17309 11658 17375 11661
rect 17718 11658 17724 11660
rect 17309 11656 17724 11658
rect 17309 11600 17314 11656
rect 17370 11600 17724 11656
rect 17309 11598 17724 11600
rect 17309 11595 17375 11598
rect 17718 11596 17724 11598
rect 17788 11596 17794 11660
rect 21766 11596 21772 11660
rect 21836 11658 21842 11660
rect 22001 11658 22067 11661
rect 21836 11656 22067 11658
rect 21836 11600 22006 11656
rect 22062 11600 22067 11656
rect 21836 11598 22067 11600
rect 21836 11596 21842 11598
rect 22001 11595 22067 11598
rect 23749 11658 23815 11661
rect 24526 11658 24532 11660
rect 23749 11656 24532 11658
rect 23749 11600 23754 11656
rect 23810 11600 24532 11656
rect 23749 11598 24532 11600
rect 23749 11595 23815 11598
rect 24526 11596 24532 11598
rect 24596 11596 24602 11660
rect 27245 11658 27311 11661
rect 28373 11658 29173 11688
rect 27245 11656 29173 11658
rect 27245 11600 27250 11656
rect 27306 11600 29173 11656
rect 27245 11598 29173 11600
rect 27245 11595 27311 11598
rect 28373 11568 29173 11598
rect 15193 11522 15259 11525
rect 15326 11522 15332 11524
rect 15193 11520 15332 11522
rect 15193 11464 15198 11520
rect 15254 11464 15332 11520
rect 15193 11462 15332 11464
rect 15193 11459 15259 11462
rect 15326 11460 15332 11462
rect 15396 11460 15402 11524
rect 15929 11522 15995 11525
rect 18454 11522 18460 11524
rect 15929 11520 18460 11522
rect 15929 11464 15934 11520
rect 15990 11464 18460 11520
rect 15929 11462 18460 11464
rect 15929 11459 15995 11462
rect 18454 11460 18460 11462
rect 18524 11460 18530 11524
rect 5436 11456 5756 11457
rect 5436 11392 5444 11456
rect 5508 11392 5524 11456
rect 5588 11392 5604 11456
rect 5668 11392 5684 11456
rect 5748 11392 5756 11456
rect 5436 11391 5756 11392
rect 14422 11456 14742 11457
rect 14422 11392 14430 11456
rect 14494 11392 14510 11456
rect 14574 11392 14590 11456
rect 14654 11392 14670 11456
rect 14734 11392 14742 11456
rect 14422 11391 14742 11392
rect 23407 11456 23727 11457
rect 23407 11392 23415 11456
rect 23479 11392 23495 11456
rect 23559 11392 23575 11456
rect 23639 11392 23655 11456
rect 23719 11392 23727 11456
rect 23407 11391 23727 11392
rect 9070 11188 9076 11252
rect 9140 11250 9146 11252
rect 9305 11250 9371 11253
rect 9140 11248 9371 11250
rect 9140 11192 9310 11248
rect 9366 11192 9371 11248
rect 9140 11190 9371 11192
rect 9140 11188 9146 11190
rect 9305 11187 9371 11190
rect 13077 11250 13143 11253
rect 19885 11250 19951 11253
rect 13077 11248 19951 11250
rect 13077 11192 13082 11248
rect 13138 11192 19890 11248
rect 19946 11192 19951 11248
rect 13077 11190 19951 11192
rect 13077 11187 13143 11190
rect 19885 11187 19951 11190
rect 7649 11116 7715 11117
rect 7598 11052 7604 11116
rect 7668 11114 7715 11116
rect 7668 11112 7760 11114
rect 7710 11056 7760 11112
rect 7668 11054 7760 11056
rect 7668 11052 7715 11054
rect 15878 11052 15884 11116
rect 15948 11114 15954 11116
rect 17309 11114 17375 11117
rect 18045 11116 18111 11117
rect 18045 11114 18092 11116
rect 15948 11112 17375 11114
rect 15948 11056 17314 11112
rect 17370 11056 17375 11112
rect 15948 11054 17375 11056
rect 18000 11112 18092 11114
rect 18000 11056 18050 11112
rect 18000 11054 18092 11056
rect 15948 11052 15954 11054
rect 7649 11051 7715 11052
rect 17309 11051 17375 11054
rect 18045 11052 18092 11054
rect 18156 11052 18162 11116
rect 21950 11114 21956 11116
rect 20900 11054 21956 11114
rect 18045 11051 18111 11052
rect 20900 10981 20960 11054
rect 21950 11052 21956 11054
rect 22020 11052 22026 11116
rect 6310 10916 6316 10980
rect 6380 10978 6386 10980
rect 8937 10978 9003 10981
rect 6380 10976 9003 10978
rect 6380 10920 8942 10976
rect 8998 10920 9003 10976
rect 6380 10918 9003 10920
rect 6380 10916 6386 10918
rect 8937 10915 9003 10918
rect 11421 10978 11487 10981
rect 11830 10978 11836 10980
rect 11421 10976 11836 10978
rect 11421 10920 11426 10976
rect 11482 10920 11836 10976
rect 11421 10918 11836 10920
rect 11421 10915 11487 10918
rect 11830 10916 11836 10918
rect 11900 10916 11906 10980
rect 12525 10978 12591 10981
rect 13445 10978 13511 10981
rect 12525 10976 13511 10978
rect 12525 10920 12530 10976
rect 12586 10920 13450 10976
rect 13506 10920 13511 10976
rect 12525 10918 13511 10920
rect 12525 10915 12591 10918
rect 13445 10915 13511 10918
rect 20897 10976 20963 10981
rect 20897 10920 20902 10976
rect 20958 10920 20963 10976
rect 20897 10915 20963 10920
rect 9929 10912 10249 10913
rect 9929 10848 9937 10912
rect 10001 10848 10017 10912
rect 10081 10848 10097 10912
rect 10161 10848 10177 10912
rect 10241 10848 10249 10912
rect 9929 10847 10249 10848
rect 18914 10912 19234 10913
rect 18914 10848 18922 10912
rect 18986 10848 19002 10912
rect 19066 10848 19082 10912
rect 19146 10848 19162 10912
rect 19226 10848 19234 10912
rect 18914 10847 19234 10848
rect 8150 10780 8156 10844
rect 8220 10842 8226 10844
rect 8845 10842 8911 10845
rect 8220 10840 8911 10842
rect 8220 10784 8850 10840
rect 8906 10784 8911 10840
rect 8220 10782 8911 10784
rect 8220 10780 8226 10782
rect 8845 10779 8911 10782
rect 10961 10842 11027 10845
rect 17861 10842 17927 10845
rect 20713 10844 20779 10845
rect 10961 10840 17927 10842
rect 10961 10784 10966 10840
rect 11022 10784 17866 10840
rect 17922 10784 17927 10840
rect 10961 10782 17927 10784
rect 10961 10779 11027 10782
rect 17861 10779 17927 10782
rect 20662 10780 20668 10844
rect 20732 10842 20779 10844
rect 20732 10840 20824 10842
rect 20774 10784 20824 10840
rect 20732 10782 20824 10784
rect 20732 10780 20779 10782
rect 20713 10779 20779 10780
rect 9949 10706 10015 10709
rect 11329 10706 11395 10709
rect 9949 10704 11395 10706
rect 9949 10648 9954 10704
rect 10010 10648 11334 10704
rect 11390 10648 11395 10704
rect 9949 10646 11395 10648
rect 9949 10643 10015 10646
rect 11329 10643 11395 10646
rect 16021 10706 16087 10709
rect 19241 10706 19307 10709
rect 16021 10704 19307 10706
rect 16021 10648 16026 10704
rect 16082 10648 19246 10704
rect 19302 10648 19307 10704
rect 16021 10646 19307 10648
rect 16021 10643 16087 10646
rect 19241 10643 19307 10646
rect 10358 10508 10364 10572
rect 10428 10570 10434 10572
rect 10685 10570 10751 10573
rect 10428 10568 10751 10570
rect 10428 10512 10690 10568
rect 10746 10512 10751 10568
rect 10428 10510 10751 10512
rect 10428 10508 10434 10510
rect 10685 10507 10751 10510
rect 17166 10508 17172 10572
rect 17236 10570 17242 10572
rect 19425 10570 19491 10573
rect 17236 10568 19491 10570
rect 17236 10512 19430 10568
rect 19486 10512 19491 10568
rect 17236 10510 19491 10512
rect 17236 10508 17242 10510
rect 19425 10507 19491 10510
rect 21173 10570 21239 10573
rect 22134 10570 22140 10572
rect 21173 10568 22140 10570
rect 21173 10512 21178 10568
rect 21234 10512 22140 10568
rect 21173 10510 22140 10512
rect 21173 10507 21239 10510
rect 22134 10508 22140 10510
rect 22204 10508 22210 10572
rect 10133 10434 10199 10437
rect 13077 10434 13143 10437
rect 10133 10432 13143 10434
rect 10133 10376 10138 10432
rect 10194 10376 13082 10432
rect 13138 10376 13143 10432
rect 10133 10374 13143 10376
rect 10133 10371 10199 10374
rect 13077 10371 13143 10374
rect 5436 10368 5756 10369
rect 5436 10304 5444 10368
rect 5508 10304 5524 10368
rect 5588 10304 5604 10368
rect 5668 10304 5684 10368
rect 5748 10304 5756 10368
rect 5436 10303 5756 10304
rect 14422 10368 14742 10369
rect 14422 10304 14430 10368
rect 14494 10304 14510 10368
rect 14574 10304 14590 10368
rect 14654 10304 14670 10368
rect 14734 10304 14742 10368
rect 14422 10303 14742 10304
rect 23407 10368 23727 10369
rect 23407 10304 23415 10368
rect 23479 10304 23495 10368
rect 23559 10304 23575 10368
rect 23639 10304 23655 10368
rect 23719 10304 23727 10368
rect 23407 10303 23727 10304
rect 3734 10100 3740 10164
rect 3804 10162 3810 10164
rect 9254 10162 9260 10164
rect 3804 10102 9260 10162
rect 3804 10100 3810 10102
rect 9254 10100 9260 10102
rect 9324 10100 9330 10164
rect 10133 10162 10199 10165
rect 11697 10162 11763 10165
rect 10133 10160 11763 10162
rect 10133 10104 10138 10160
rect 10194 10104 11702 10160
rect 11758 10104 11763 10160
rect 10133 10102 11763 10104
rect 10133 10099 10199 10102
rect 11697 10099 11763 10102
rect 14089 10162 14155 10165
rect 14825 10162 14891 10165
rect 14089 10160 14891 10162
rect 14089 10104 14094 10160
rect 14150 10104 14830 10160
rect 14886 10104 14891 10160
rect 14089 10102 14891 10104
rect 14089 10099 14155 10102
rect 14825 10099 14891 10102
rect 16665 10162 16731 10165
rect 19333 10162 19399 10165
rect 16665 10160 19399 10162
rect 16665 10104 16670 10160
rect 16726 10104 19338 10160
rect 19394 10104 19399 10160
rect 16665 10102 19399 10104
rect 16665 10099 16731 10102
rect 19333 10099 19399 10102
rect 21909 10162 21975 10165
rect 24485 10162 24551 10165
rect 21909 10160 24551 10162
rect 21909 10104 21914 10160
rect 21970 10104 24490 10160
rect 24546 10104 24551 10160
rect 21909 10102 24551 10104
rect 21909 10099 21975 10102
rect 24485 10099 24551 10102
rect 2814 9964 2820 10028
rect 2884 10026 2890 10028
rect 3049 10026 3115 10029
rect 2884 10024 3115 10026
rect 2884 9968 3054 10024
rect 3110 9968 3115 10024
rect 2884 9966 3115 9968
rect 2884 9964 2890 9966
rect 3049 9963 3115 9966
rect 6126 9964 6132 10028
rect 6196 10026 6202 10028
rect 6269 10026 6335 10029
rect 6196 10024 6335 10026
rect 6196 9968 6274 10024
rect 6330 9968 6335 10024
rect 6196 9966 6335 9968
rect 6196 9964 6202 9966
rect 6269 9963 6335 9966
rect 6913 10026 6979 10029
rect 7046 10026 7052 10028
rect 6913 10024 7052 10026
rect 6913 9968 6918 10024
rect 6974 9968 7052 10024
rect 6913 9966 7052 9968
rect 6913 9963 6979 9966
rect 7046 9964 7052 9966
rect 7116 9964 7122 10028
rect 12341 10026 12407 10029
rect 13537 10026 13603 10029
rect 14181 10026 14247 10029
rect 12341 10024 14247 10026
rect 12341 9968 12346 10024
rect 12402 9968 13542 10024
rect 13598 9968 14186 10024
rect 14242 9968 14247 10024
rect 12341 9966 14247 9968
rect 12341 9963 12407 9966
rect 13537 9963 13603 9966
rect 14181 9963 14247 9966
rect 17769 10026 17835 10029
rect 19425 10026 19491 10029
rect 17769 10024 19491 10026
rect 17769 9968 17774 10024
rect 17830 9968 19430 10024
rect 19486 9968 19491 10024
rect 17769 9966 19491 9968
rect 17769 9963 17835 9966
rect 19425 9963 19491 9966
rect 4797 9890 4863 9893
rect 5206 9890 5212 9892
rect 4797 9888 5212 9890
rect 4797 9832 4802 9888
rect 4858 9832 5212 9888
rect 4797 9830 5212 9832
rect 4797 9827 4863 9830
rect 5206 9828 5212 9830
rect 5276 9828 5282 9892
rect 7966 9828 7972 9892
rect 8036 9890 8042 9892
rect 8109 9890 8175 9893
rect 8036 9888 8175 9890
rect 8036 9832 8114 9888
rect 8170 9832 8175 9888
rect 8036 9830 8175 9832
rect 8036 9828 8042 9830
rect 8109 9827 8175 9830
rect 10317 9892 10383 9893
rect 10317 9888 10364 9892
rect 10428 9890 10434 9892
rect 10317 9832 10322 9888
rect 10317 9828 10364 9832
rect 10428 9830 10474 9890
rect 10428 9828 10434 9830
rect 14038 9828 14044 9892
rect 14108 9890 14114 9892
rect 14549 9890 14615 9893
rect 14108 9888 14615 9890
rect 14108 9832 14554 9888
rect 14610 9832 14615 9888
rect 14108 9830 14615 9832
rect 14108 9828 14114 9830
rect 10317 9827 10383 9828
rect 14549 9827 14615 9830
rect 9929 9824 10249 9825
rect 9929 9760 9937 9824
rect 10001 9760 10017 9824
rect 10081 9760 10097 9824
rect 10161 9760 10177 9824
rect 10241 9760 10249 9824
rect 9929 9759 10249 9760
rect 18914 9824 19234 9825
rect 18914 9760 18922 9824
rect 18986 9760 19002 9824
rect 19066 9760 19082 9824
rect 19146 9760 19162 9824
rect 19226 9760 19234 9824
rect 18914 9759 19234 9760
rect 5073 9756 5139 9757
rect 5022 9754 5028 9756
rect 4982 9694 5028 9754
rect 5092 9752 5139 9756
rect 5134 9696 5139 9752
rect 5022 9692 5028 9694
rect 5092 9692 5139 9696
rect 5073 9691 5139 9692
rect 10317 9754 10383 9757
rect 11094 9754 11100 9756
rect 10317 9752 11100 9754
rect 10317 9696 10322 9752
rect 10378 9696 11100 9752
rect 10317 9694 11100 9696
rect 10317 9691 10383 9694
rect 11094 9692 11100 9694
rect 11164 9692 11170 9756
rect 20437 9754 20503 9757
rect 25865 9754 25931 9757
rect 20437 9752 25931 9754
rect 20437 9696 20442 9752
rect 20498 9696 25870 9752
rect 25926 9696 25931 9752
rect 20437 9694 25931 9696
rect 20437 9691 20503 9694
rect 25865 9691 25931 9694
rect 18638 9556 18644 9620
rect 18708 9618 18714 9620
rect 22369 9618 22435 9621
rect 18708 9616 22435 9618
rect 18708 9560 22374 9616
rect 22430 9560 22435 9616
rect 18708 9558 22435 9560
rect 18708 9556 18714 9558
rect 22369 9555 22435 9558
rect 23289 9618 23355 9621
rect 23974 9618 23980 9620
rect 23289 9616 23980 9618
rect 23289 9560 23294 9616
rect 23350 9560 23980 9616
rect 23289 9558 23980 9560
rect 23289 9555 23355 9558
rect 23974 9556 23980 9558
rect 24044 9556 24050 9620
rect 10225 9482 10291 9485
rect 11513 9482 11579 9485
rect 10225 9480 11579 9482
rect 10225 9424 10230 9480
rect 10286 9424 11518 9480
rect 11574 9424 11579 9480
rect 10225 9422 11579 9424
rect 10225 9419 10291 9422
rect 11513 9419 11579 9422
rect 21950 9420 21956 9484
rect 22020 9482 22026 9484
rect 23749 9482 23815 9485
rect 22020 9480 23815 9482
rect 22020 9424 23754 9480
rect 23810 9424 23815 9480
rect 22020 9422 23815 9424
rect 22020 9420 22026 9422
rect 23749 9419 23815 9422
rect 9857 9346 9923 9349
rect 11789 9346 11855 9349
rect 9857 9344 11855 9346
rect 9857 9288 9862 9344
rect 9918 9288 11794 9344
rect 11850 9288 11855 9344
rect 9857 9286 11855 9288
rect 9857 9283 9923 9286
rect 11789 9283 11855 9286
rect 5436 9280 5756 9281
rect 5436 9216 5444 9280
rect 5508 9216 5524 9280
rect 5588 9216 5604 9280
rect 5668 9216 5684 9280
rect 5748 9216 5756 9280
rect 5436 9215 5756 9216
rect 14422 9280 14742 9281
rect 14422 9216 14430 9280
rect 14494 9216 14510 9280
rect 14574 9216 14590 9280
rect 14654 9216 14670 9280
rect 14734 9216 14742 9280
rect 14422 9215 14742 9216
rect 23407 9280 23727 9281
rect 23407 9216 23415 9280
rect 23479 9216 23495 9280
rect 23559 9216 23575 9280
rect 23639 9216 23655 9280
rect 23719 9216 23727 9280
rect 23407 9215 23727 9216
rect 12341 9074 12407 9077
rect 12525 9074 12591 9077
rect 12341 9072 12591 9074
rect 12341 9016 12346 9072
rect 12402 9016 12530 9072
rect 12586 9016 12591 9072
rect 12341 9014 12591 9016
rect 12341 9011 12407 9014
rect 12525 9011 12591 9014
rect 15694 9012 15700 9076
rect 15764 9074 15770 9076
rect 15837 9074 15903 9077
rect 15764 9072 15903 9074
rect 15764 9016 15842 9072
rect 15898 9016 15903 9072
rect 15764 9014 15903 9016
rect 15764 9012 15770 9014
rect 15837 9011 15903 9014
rect 19241 9074 19307 9077
rect 21633 9074 21699 9077
rect 19241 9072 21699 9074
rect 19241 9016 19246 9072
rect 19302 9016 21638 9072
rect 21694 9016 21699 9072
rect 19241 9014 21699 9016
rect 19241 9011 19307 9014
rect 21633 9011 21699 9014
rect 1669 8938 1735 8941
rect 2221 8938 2287 8941
rect 9581 8938 9647 8941
rect 1669 8936 9647 8938
rect 1669 8880 1674 8936
rect 1730 8880 2226 8936
rect 2282 8880 9586 8936
rect 9642 8880 9647 8936
rect 1669 8878 9647 8880
rect 1669 8875 1735 8878
rect 2221 8875 2287 8878
rect 9581 8875 9647 8878
rect 11789 8938 11855 8941
rect 16798 8938 16804 8940
rect 11789 8936 16804 8938
rect 11789 8880 11794 8936
rect 11850 8880 16804 8936
rect 11789 8878 16804 8880
rect 11789 8875 11855 8878
rect 16798 8876 16804 8878
rect 16868 8876 16874 8940
rect 18454 8876 18460 8940
rect 18524 8938 18530 8940
rect 18689 8938 18755 8941
rect 18524 8936 18755 8938
rect 18524 8880 18694 8936
rect 18750 8880 18755 8936
rect 18524 8878 18755 8880
rect 18524 8876 18530 8878
rect 18689 8875 18755 8878
rect 20437 8802 20503 8805
rect 24117 8802 24183 8805
rect 20437 8800 24183 8802
rect 20437 8744 20442 8800
rect 20498 8744 24122 8800
rect 24178 8744 24183 8800
rect 20437 8742 24183 8744
rect 20437 8739 20503 8742
rect 24117 8739 24183 8742
rect 9929 8736 10249 8737
rect 9929 8672 9937 8736
rect 10001 8672 10017 8736
rect 10081 8672 10097 8736
rect 10161 8672 10177 8736
rect 10241 8672 10249 8736
rect 9929 8671 10249 8672
rect 18914 8736 19234 8737
rect 18914 8672 18922 8736
rect 18986 8672 19002 8736
rect 19066 8672 19082 8736
rect 19146 8672 19162 8736
rect 19226 8672 19234 8736
rect 18914 8671 19234 8672
rect 11053 8666 11119 8669
rect 13905 8666 13971 8669
rect 11053 8664 13971 8666
rect 11053 8608 11058 8664
rect 11114 8608 13910 8664
rect 13966 8608 13971 8664
rect 11053 8606 13971 8608
rect 11053 8603 11119 8606
rect 13905 8603 13971 8606
rect 23657 8666 23723 8669
rect 25313 8666 25379 8669
rect 23657 8664 25379 8666
rect 23657 8608 23662 8664
rect 23718 8608 25318 8664
rect 25374 8608 25379 8664
rect 23657 8606 25379 8608
rect 23657 8603 23723 8606
rect 25313 8603 25379 8606
rect 2814 8468 2820 8532
rect 2884 8530 2890 8532
rect 3734 8530 3740 8532
rect 2884 8470 3740 8530
rect 2884 8468 2890 8470
rect 3734 8468 3740 8470
rect 3804 8530 3810 8532
rect 3969 8530 4035 8533
rect 6361 8530 6427 8533
rect 6545 8530 6611 8533
rect 3804 8528 4538 8530
rect 3804 8472 3974 8528
rect 4030 8472 4538 8528
rect 3804 8470 4538 8472
rect 3804 8468 3810 8470
rect 3969 8467 4035 8470
rect 4245 8394 4311 8397
rect 4110 8392 4311 8394
rect 4110 8336 4250 8392
rect 4306 8336 4311 8392
rect 4110 8334 4311 8336
rect 4478 8394 4538 8470
rect 6361 8528 6611 8530
rect 6361 8472 6366 8528
rect 6422 8472 6550 8528
rect 6606 8472 6611 8528
rect 6361 8470 6611 8472
rect 6361 8467 6427 8470
rect 6545 8467 6611 8470
rect 6913 8530 6979 8533
rect 7557 8530 7623 8533
rect 6913 8528 7623 8530
rect 6913 8472 6918 8528
rect 6974 8472 7562 8528
rect 7618 8472 7623 8528
rect 6913 8470 7623 8472
rect 6913 8467 6979 8470
rect 7557 8467 7623 8470
rect 9254 8468 9260 8532
rect 9324 8530 9330 8532
rect 10133 8530 10199 8533
rect 9324 8528 10199 8530
rect 9324 8472 10138 8528
rect 10194 8472 10199 8528
rect 9324 8470 10199 8472
rect 9324 8468 9330 8470
rect 10133 8467 10199 8470
rect 9489 8394 9555 8397
rect 4478 8392 9555 8394
rect 4478 8336 9494 8392
rect 9550 8336 9555 8392
rect 4478 8334 9555 8336
rect 4110 7173 4170 8334
rect 4245 8331 4311 8334
rect 9489 8331 9555 8334
rect 10041 8394 10107 8397
rect 10358 8394 10364 8396
rect 10041 8392 10364 8394
rect 10041 8336 10046 8392
rect 10102 8336 10364 8392
rect 10041 8334 10364 8336
rect 10041 8331 10107 8334
rect 10358 8332 10364 8334
rect 10428 8332 10434 8396
rect 11462 8332 11468 8396
rect 11532 8394 11538 8396
rect 11605 8394 11671 8397
rect 11532 8392 11671 8394
rect 11532 8336 11610 8392
rect 11666 8336 11671 8392
rect 11532 8334 11671 8336
rect 11532 8332 11538 8334
rect 11605 8331 11671 8334
rect 12341 8394 12407 8397
rect 13169 8394 13235 8397
rect 15837 8394 15903 8397
rect 12341 8392 15903 8394
rect 12341 8336 12346 8392
rect 12402 8336 13174 8392
rect 13230 8336 15842 8392
rect 15898 8336 15903 8392
rect 12341 8334 15903 8336
rect 12341 8331 12407 8334
rect 13169 8331 13235 8334
rect 13169 8258 13235 8261
rect 14089 8258 14155 8261
rect 13169 8256 14155 8258
rect 13169 8200 13174 8256
rect 13230 8200 14094 8256
rect 14150 8200 14155 8256
rect 13169 8198 14155 8200
rect 13169 8195 13235 8198
rect 14089 8195 14155 8198
rect 5436 8192 5756 8193
rect 5436 8128 5444 8192
rect 5508 8128 5524 8192
rect 5588 8128 5604 8192
rect 5668 8128 5684 8192
rect 5748 8128 5756 8192
rect 5436 8127 5756 8128
rect 14230 8125 14290 8334
rect 15837 8331 15903 8334
rect 23381 8394 23447 8397
rect 25313 8394 25379 8397
rect 23381 8392 25379 8394
rect 23381 8336 23386 8392
rect 23442 8336 25318 8392
rect 25374 8336 25379 8392
rect 23381 8334 25379 8336
rect 23381 8331 23447 8334
rect 25313 8331 25379 8334
rect 19425 8258 19491 8261
rect 19558 8258 19564 8260
rect 19425 8256 19564 8258
rect 19425 8200 19430 8256
rect 19486 8200 19564 8256
rect 19425 8198 19564 8200
rect 19425 8195 19491 8198
rect 19558 8196 19564 8198
rect 19628 8196 19634 8260
rect 20662 8196 20668 8260
rect 20732 8258 20738 8260
rect 22318 8258 22324 8260
rect 20732 8198 22324 8258
rect 20732 8196 20738 8198
rect 22318 8196 22324 8198
rect 22388 8196 22394 8260
rect 14422 8192 14742 8193
rect 14422 8128 14430 8192
rect 14494 8128 14510 8192
rect 14574 8128 14590 8192
rect 14654 8128 14670 8192
rect 14734 8128 14742 8192
rect 14422 8127 14742 8128
rect 23407 8192 23727 8193
rect 23407 8128 23415 8192
rect 23479 8128 23495 8192
rect 23559 8128 23575 8192
rect 23639 8128 23655 8192
rect 23719 8128 23727 8192
rect 23407 8127 23727 8128
rect 14181 8120 14290 8125
rect 14181 8064 14186 8120
rect 14242 8064 14290 8120
rect 14181 8062 14290 8064
rect 14181 8059 14247 8062
rect 14222 7924 14228 7988
rect 14292 7986 14298 7988
rect 14365 7986 14431 7989
rect 14292 7984 14431 7986
rect 14292 7928 14370 7984
rect 14426 7928 14431 7984
rect 14292 7926 14431 7928
rect 14292 7924 14298 7926
rect 14365 7923 14431 7926
rect 22001 7986 22067 7989
rect 22870 7986 22876 7988
rect 22001 7984 22876 7986
rect 22001 7928 22006 7984
rect 22062 7928 22876 7984
rect 22001 7926 22876 7928
rect 22001 7923 22067 7926
rect 22870 7924 22876 7926
rect 22940 7924 22946 7988
rect 23657 7986 23723 7989
rect 26233 7986 26299 7989
rect 23657 7984 26299 7986
rect 23657 7928 23662 7984
rect 23718 7928 26238 7984
rect 26294 7928 26299 7984
rect 23657 7926 26299 7928
rect 23657 7923 23723 7926
rect 26233 7923 26299 7926
rect 16849 7714 16915 7717
rect 16806 7712 16915 7714
rect 16806 7656 16854 7712
rect 16910 7656 16915 7712
rect 16806 7651 16915 7656
rect 21725 7714 21791 7717
rect 25957 7714 26023 7717
rect 21725 7712 26023 7714
rect 21725 7656 21730 7712
rect 21786 7656 25962 7712
rect 26018 7656 26023 7712
rect 21725 7654 26023 7656
rect 21725 7651 21791 7654
rect 25957 7651 26023 7654
rect 9929 7648 10249 7649
rect 9929 7584 9937 7648
rect 10001 7584 10017 7648
rect 10081 7584 10097 7648
rect 10161 7584 10177 7648
rect 10241 7584 10249 7648
rect 9929 7583 10249 7584
rect 16806 7445 16866 7651
rect 18914 7648 19234 7649
rect 18914 7584 18922 7648
rect 18986 7584 19002 7648
rect 19066 7584 19082 7648
rect 19146 7584 19162 7648
rect 19226 7584 19234 7648
rect 18914 7583 19234 7584
rect 27337 7578 27403 7581
rect 27337 7576 27584 7578
rect 27337 7520 27342 7576
rect 27398 7520 27584 7576
rect 27337 7518 27584 7520
rect 27337 7515 27403 7518
rect 6862 7380 6868 7444
rect 6932 7442 6938 7444
rect 7281 7442 7347 7445
rect 6932 7440 7347 7442
rect 6932 7384 7286 7440
rect 7342 7384 7347 7440
rect 6932 7382 7347 7384
rect 6932 7380 6938 7382
rect 7281 7379 7347 7382
rect 16757 7440 16866 7445
rect 16757 7384 16762 7440
rect 16818 7384 16866 7440
rect 16757 7382 16866 7384
rect 16757 7379 16823 7382
rect 19926 7380 19932 7444
rect 19996 7442 20002 7444
rect 20345 7442 20411 7445
rect 19996 7440 20411 7442
rect 19996 7384 20350 7440
rect 20406 7384 20411 7440
rect 19996 7382 20411 7384
rect 19996 7380 20002 7382
rect 20345 7379 20411 7382
rect 20805 7442 20871 7445
rect 24945 7442 25011 7445
rect 25262 7442 25268 7444
rect 20805 7440 21328 7442
rect 20805 7384 20810 7440
rect 20866 7384 21328 7440
rect 20805 7382 21328 7384
rect 20805 7379 20871 7382
rect 7598 7244 7604 7308
rect 7668 7306 7674 7308
rect 7741 7306 7807 7309
rect 7668 7304 7807 7306
rect 7668 7248 7746 7304
rect 7802 7248 7807 7304
rect 7668 7246 7807 7248
rect 7668 7244 7674 7246
rect 7741 7243 7807 7246
rect 16941 7306 17007 7309
rect 17902 7306 17908 7308
rect 16941 7304 17908 7306
rect 16941 7248 16946 7304
rect 17002 7248 17908 7304
rect 16941 7246 17908 7248
rect 16941 7243 17007 7246
rect 17902 7244 17908 7246
rect 17972 7244 17978 7308
rect 21268 7306 21328 7382
rect 24945 7440 25268 7442
rect 24945 7384 24950 7440
rect 25006 7384 25268 7440
rect 24945 7382 25268 7384
rect 24945 7379 25011 7382
rect 25262 7380 25268 7382
rect 25332 7380 25338 7444
rect 27524 7309 27584 7518
rect 21541 7306 21607 7309
rect 21268 7304 21607 7306
rect 21268 7248 21546 7304
rect 21602 7248 21607 7304
rect 21268 7246 21607 7248
rect 21541 7243 21607 7246
rect 21725 7306 21791 7309
rect 25497 7306 25563 7309
rect 21725 7304 25563 7306
rect 21725 7248 21730 7304
rect 21786 7248 25502 7304
rect 25558 7248 25563 7304
rect 21725 7246 25563 7248
rect 21725 7243 21791 7246
rect 25497 7243 25563 7246
rect 27521 7304 27587 7309
rect 27521 7248 27526 7304
rect 27582 7248 27587 7304
rect 27521 7243 27587 7248
rect 4061 7168 4170 7173
rect 4061 7112 4066 7168
rect 4122 7112 4170 7168
rect 4061 7110 4170 7112
rect 24301 7170 24367 7173
rect 24669 7170 24735 7173
rect 24301 7168 24735 7170
rect 24301 7112 24306 7168
rect 24362 7112 24674 7168
rect 24730 7112 24735 7168
rect 24301 7110 24735 7112
rect 4061 7107 4127 7110
rect 24301 7107 24367 7110
rect 24669 7107 24735 7110
rect 5436 7104 5756 7105
rect 5436 7040 5444 7104
rect 5508 7040 5524 7104
rect 5588 7040 5604 7104
rect 5668 7040 5684 7104
rect 5748 7040 5756 7104
rect 5436 7039 5756 7040
rect 14422 7104 14742 7105
rect 14422 7040 14430 7104
rect 14494 7040 14510 7104
rect 14574 7040 14590 7104
rect 14654 7040 14670 7104
rect 14734 7040 14742 7104
rect 14422 7039 14742 7040
rect 23407 7104 23727 7105
rect 23407 7040 23415 7104
rect 23479 7040 23495 7104
rect 23559 7040 23575 7104
rect 23639 7040 23655 7104
rect 23719 7040 23727 7104
rect 23407 7039 23727 7040
rect 24577 7034 24643 7037
rect 24396 7032 24643 7034
rect 24396 6976 24582 7032
rect 24638 6976 24643 7032
rect 24396 6974 24643 6976
rect 24396 6901 24456 6974
rect 24577 6971 24643 6974
rect 3049 6898 3115 6901
rect 3006 6896 3115 6898
rect 3006 6840 3054 6896
rect 3110 6840 3115 6896
rect 3006 6835 3115 6840
rect 3233 6898 3299 6901
rect 3366 6898 3372 6900
rect 3233 6896 3372 6898
rect 3233 6840 3238 6896
rect 3294 6840 3372 6896
rect 3233 6838 3372 6840
rect 3233 6835 3299 6838
rect 3366 6836 3372 6838
rect 3436 6836 3442 6900
rect 3601 6898 3667 6901
rect 3734 6898 3740 6900
rect 3601 6896 3740 6898
rect 3601 6840 3606 6896
rect 3662 6840 3740 6896
rect 3601 6838 3740 6840
rect 3601 6835 3667 6838
rect 3734 6836 3740 6838
rect 3804 6836 3810 6900
rect 5073 6898 5139 6901
rect 11145 6898 11211 6901
rect 5073 6896 11211 6898
rect 5073 6840 5078 6896
rect 5134 6840 11150 6896
rect 11206 6840 11211 6896
rect 5073 6838 11211 6840
rect 5073 6835 5139 6838
rect 11145 6835 11211 6838
rect 24393 6896 24459 6901
rect 24393 6840 24398 6896
rect 24454 6840 24459 6896
rect 24393 6835 24459 6840
rect 3006 6490 3066 6835
rect 5901 6762 5967 6765
rect 7005 6762 7071 6765
rect 5901 6760 7071 6762
rect 5901 6704 5906 6760
rect 5962 6704 7010 6760
rect 7066 6704 7071 6760
rect 5901 6702 7071 6704
rect 5901 6699 5967 6702
rect 7005 6699 7071 6702
rect 11697 6762 11763 6765
rect 17861 6762 17927 6765
rect 11697 6760 17927 6762
rect 11697 6704 11702 6760
rect 11758 6704 17866 6760
rect 17922 6704 17927 6760
rect 11697 6702 17927 6704
rect 11697 6699 11763 6702
rect 17861 6699 17927 6702
rect 18229 6762 18295 6765
rect 24761 6762 24827 6765
rect 25037 6762 25103 6765
rect 18229 6760 22110 6762
rect 18229 6704 18234 6760
rect 18290 6704 22110 6760
rect 18229 6702 22110 6704
rect 18229 6699 18295 6702
rect 16665 6626 16731 6629
rect 17861 6626 17927 6629
rect 16665 6624 17927 6626
rect 16665 6568 16670 6624
rect 16726 6568 17866 6624
rect 17922 6568 17927 6624
rect 16665 6566 17927 6568
rect 22050 6626 22110 6702
rect 24761 6760 25103 6762
rect 24761 6704 24766 6760
rect 24822 6704 25042 6760
rect 25098 6704 25103 6760
rect 24761 6702 25103 6704
rect 24761 6699 24827 6702
rect 25037 6699 25103 6702
rect 24393 6626 24459 6629
rect 22050 6624 24459 6626
rect 22050 6568 24398 6624
rect 24454 6568 24459 6624
rect 22050 6566 24459 6568
rect 16665 6563 16731 6566
rect 17861 6563 17927 6566
rect 24393 6563 24459 6566
rect 9929 6560 10249 6561
rect 9929 6496 9937 6560
rect 10001 6496 10017 6560
rect 10081 6496 10097 6560
rect 10161 6496 10177 6560
rect 10241 6496 10249 6560
rect 9929 6495 10249 6496
rect 18914 6560 19234 6561
rect 18914 6496 18922 6560
rect 18986 6496 19002 6560
rect 19066 6496 19082 6560
rect 19146 6496 19162 6560
rect 19226 6496 19234 6560
rect 18914 6495 19234 6496
rect 3325 6490 3391 6493
rect 3006 6488 3391 6490
rect 3006 6432 3330 6488
rect 3386 6432 3391 6488
rect 3006 6430 3391 6432
rect 3325 6427 3391 6430
rect 21357 6490 21423 6493
rect 23289 6490 23355 6493
rect 25037 6492 25103 6493
rect 25037 6490 25084 6492
rect 21357 6488 23355 6490
rect 21357 6432 21362 6488
rect 21418 6432 23294 6488
rect 23350 6432 23355 6488
rect 21357 6430 23355 6432
rect 24992 6488 25084 6490
rect 24992 6432 25042 6488
rect 24992 6430 25084 6432
rect 21357 6427 21423 6430
rect 23289 6427 23355 6430
rect 25037 6428 25084 6430
rect 25148 6428 25154 6492
rect 27337 6490 27403 6493
rect 27470 6490 27476 6492
rect 27337 6488 27476 6490
rect 27337 6432 27342 6488
rect 27398 6432 27476 6488
rect 27337 6430 27476 6432
rect 25037 6427 25103 6428
rect 27337 6427 27403 6430
rect 27470 6428 27476 6430
rect 27540 6428 27546 6492
rect 1393 6354 1459 6357
rect 8937 6354 9003 6357
rect 1393 6352 9003 6354
rect 1393 6296 1398 6352
rect 1454 6296 8942 6352
rect 8998 6296 9003 6352
rect 1393 6294 9003 6296
rect 1393 6291 1459 6294
rect 8937 6291 9003 6294
rect 12985 6354 13051 6357
rect 15561 6354 15627 6357
rect 17861 6354 17927 6357
rect 12985 6352 15627 6354
rect 12985 6296 12990 6352
rect 13046 6296 15566 6352
rect 15622 6296 15627 6352
rect 12985 6294 15627 6296
rect 12985 6291 13051 6294
rect 15561 6291 15627 6294
rect 16622 6352 17927 6354
rect 16622 6296 17866 6352
rect 17922 6296 17927 6352
rect 16622 6294 17927 6296
rect 10225 6218 10291 6221
rect 14733 6218 14799 6221
rect 15929 6218 15995 6221
rect 16622 6218 16682 6294
rect 17861 6291 17927 6294
rect 18137 6354 18203 6357
rect 20989 6354 21055 6357
rect 18137 6352 21055 6354
rect 18137 6296 18142 6352
rect 18198 6296 20994 6352
rect 21050 6296 21055 6352
rect 18137 6294 21055 6296
rect 18137 6291 18203 6294
rect 20989 6291 21055 6294
rect 22645 6354 22711 6357
rect 26049 6354 26115 6357
rect 22645 6352 26115 6354
rect 22645 6296 22650 6352
rect 22706 6296 26054 6352
rect 26110 6296 26115 6352
rect 22645 6294 26115 6296
rect 22645 6291 22711 6294
rect 26049 6291 26115 6294
rect 10225 6216 16682 6218
rect 10225 6160 10230 6216
rect 10286 6160 14738 6216
rect 14794 6160 15934 6216
rect 15990 6160 16682 6216
rect 10225 6158 16682 6160
rect 16757 6218 16823 6221
rect 23790 6218 23796 6220
rect 16757 6216 23796 6218
rect 16757 6160 16762 6216
rect 16818 6160 23796 6216
rect 16757 6158 23796 6160
rect 10225 6155 10291 6158
rect 14733 6155 14799 6158
rect 15929 6155 15995 6158
rect 16757 6155 16823 6158
rect 23790 6156 23796 6158
rect 23860 6156 23866 6220
rect 17953 6082 18019 6085
rect 18086 6082 18092 6084
rect 17953 6080 18092 6082
rect 17953 6024 17958 6080
rect 18014 6024 18092 6080
rect 17953 6022 18092 6024
rect 17953 6019 18019 6022
rect 18086 6020 18092 6022
rect 18156 6020 18162 6084
rect 20110 6020 20116 6084
rect 20180 6082 20186 6084
rect 22277 6082 22343 6085
rect 20180 6080 22343 6082
rect 20180 6024 22282 6080
rect 22338 6024 22343 6080
rect 20180 6022 22343 6024
rect 20180 6020 20186 6022
rect 22277 6019 22343 6022
rect 5436 6016 5756 6017
rect 5436 5952 5444 6016
rect 5508 5952 5524 6016
rect 5588 5952 5604 6016
rect 5668 5952 5684 6016
rect 5748 5952 5756 6016
rect 5436 5951 5756 5952
rect 14422 6016 14742 6017
rect 14422 5952 14430 6016
rect 14494 5952 14510 6016
rect 14574 5952 14590 6016
rect 14654 5952 14670 6016
rect 14734 5952 14742 6016
rect 14422 5951 14742 5952
rect 23407 6016 23727 6017
rect 23407 5952 23415 6016
rect 23479 5952 23495 6016
rect 23559 5952 23575 6016
rect 23639 5952 23655 6016
rect 23719 5952 23727 6016
rect 23407 5951 23727 5952
rect 20989 5948 21055 5949
rect 22461 5948 22527 5949
rect 20989 5946 21036 5948
rect 20944 5944 21036 5946
rect 20944 5888 20994 5944
rect 20944 5886 21036 5888
rect 20989 5884 21036 5886
rect 21100 5884 21106 5948
rect 22461 5946 22508 5948
rect 22416 5944 22508 5946
rect 22416 5888 22466 5944
rect 22416 5886 22508 5888
rect 22461 5884 22508 5886
rect 22572 5884 22578 5948
rect 20989 5883 21055 5884
rect 22461 5883 22527 5884
rect 14365 5810 14431 5813
rect 15101 5810 15167 5813
rect 14365 5808 15167 5810
rect 14365 5752 14370 5808
rect 14426 5752 15106 5808
rect 15162 5752 15167 5808
rect 14365 5750 15167 5752
rect 14365 5747 14431 5750
rect 15101 5747 15167 5750
rect 21357 5810 21423 5813
rect 23105 5810 23171 5813
rect 21357 5808 23171 5810
rect 21357 5752 21362 5808
rect 21418 5752 23110 5808
rect 23166 5752 23171 5808
rect 21357 5750 23171 5752
rect 21357 5747 21423 5750
rect 23105 5747 23171 5750
rect 2957 5676 3023 5677
rect 2957 5674 3004 5676
rect 2912 5672 3004 5674
rect 2912 5616 2962 5672
rect 2912 5614 3004 5616
rect 2957 5612 3004 5614
rect 3068 5612 3074 5676
rect 3550 5612 3556 5676
rect 3620 5674 3626 5676
rect 9673 5674 9739 5677
rect 3620 5672 9739 5674
rect 3620 5616 9678 5672
rect 9734 5616 9739 5672
rect 3620 5614 9739 5616
rect 3620 5612 3626 5614
rect 2957 5611 3023 5612
rect 9673 5611 9739 5614
rect 9949 5674 10015 5677
rect 15653 5674 15719 5677
rect 18270 5674 18276 5676
rect 9949 5672 10426 5674
rect 9949 5616 9954 5672
rect 10010 5616 10426 5672
rect 9949 5614 10426 5616
rect 9949 5611 10015 5614
rect 9929 5472 10249 5473
rect 9929 5408 9937 5472
rect 10001 5408 10017 5472
rect 10081 5408 10097 5472
rect 10161 5408 10177 5472
rect 10241 5408 10249 5472
rect 9929 5407 10249 5408
rect 2773 5402 2839 5405
rect 7281 5402 7347 5405
rect 2773 5400 7347 5402
rect 2773 5344 2778 5400
rect 2834 5344 7286 5400
rect 7342 5344 7347 5400
rect 2773 5342 7347 5344
rect 2773 5339 2839 5342
rect 7281 5339 7347 5342
rect 3785 5266 3851 5269
rect 3742 5264 3851 5266
rect 3742 5208 3790 5264
rect 3846 5208 3851 5264
rect 3742 5203 3851 5208
rect 10225 5266 10291 5269
rect 10366 5266 10426 5614
rect 15653 5672 18276 5674
rect 15653 5616 15658 5672
rect 15714 5616 18276 5672
rect 15653 5614 18276 5616
rect 15653 5611 15719 5614
rect 18270 5612 18276 5614
rect 18340 5612 18346 5676
rect 21817 5674 21883 5677
rect 21950 5674 21956 5676
rect 21817 5672 21956 5674
rect 21817 5616 21822 5672
rect 21878 5616 21956 5672
rect 21817 5614 21956 5616
rect 21817 5611 21883 5614
rect 21950 5612 21956 5614
rect 22020 5612 22026 5676
rect 17033 5538 17099 5541
rect 17350 5538 17356 5540
rect 17033 5536 17356 5538
rect 17033 5480 17038 5536
rect 17094 5480 17356 5536
rect 17033 5478 17356 5480
rect 17033 5475 17099 5478
rect 17350 5476 17356 5478
rect 17420 5476 17426 5540
rect 20253 5538 20319 5541
rect 20662 5538 20668 5540
rect 20253 5536 20668 5538
rect 20253 5480 20258 5536
rect 20314 5480 20668 5536
rect 20253 5478 20668 5480
rect 20253 5475 20319 5478
rect 20662 5476 20668 5478
rect 20732 5476 20738 5540
rect 23473 5538 23539 5541
rect 25405 5538 25471 5541
rect 23473 5536 25471 5538
rect 23473 5480 23478 5536
rect 23534 5480 25410 5536
rect 25466 5480 25471 5536
rect 23473 5478 25471 5480
rect 23473 5475 23539 5478
rect 25405 5475 25471 5478
rect 18914 5472 19234 5473
rect 18914 5408 18922 5472
rect 18986 5408 19002 5472
rect 19066 5408 19082 5472
rect 19146 5408 19162 5472
rect 19226 5408 19234 5472
rect 18914 5407 19234 5408
rect 20478 5340 20484 5404
rect 20548 5402 20554 5404
rect 20621 5402 20687 5405
rect 20548 5400 20687 5402
rect 20548 5344 20626 5400
rect 20682 5344 20687 5400
rect 20548 5342 20687 5344
rect 20548 5340 20554 5342
rect 20621 5339 20687 5342
rect 21909 5402 21975 5405
rect 25681 5402 25747 5405
rect 21909 5400 25747 5402
rect 21909 5344 21914 5400
rect 21970 5344 25686 5400
rect 25742 5344 25747 5400
rect 21909 5342 25747 5344
rect 21909 5339 21975 5342
rect 25681 5339 25747 5342
rect 10225 5264 10426 5266
rect 10225 5208 10230 5264
rect 10286 5208 10426 5264
rect 10225 5206 10426 5208
rect 10225 5203 10291 5206
rect 10542 5204 10548 5268
rect 10612 5266 10618 5268
rect 10777 5266 10843 5269
rect 10612 5264 10843 5266
rect 10612 5208 10782 5264
rect 10838 5208 10843 5264
rect 10612 5206 10843 5208
rect 10612 5204 10618 5206
rect 10777 5203 10843 5206
rect 19977 5266 20043 5269
rect 22277 5266 22343 5269
rect 19977 5264 22343 5266
rect 19977 5208 19982 5264
rect 20038 5208 22282 5264
rect 22338 5208 22343 5264
rect 19977 5206 22343 5208
rect 19977 5203 20043 5206
rect 22277 5203 22343 5206
rect 3601 5130 3667 5133
rect 3742 5130 3802 5203
rect 3601 5128 3802 5130
rect 3601 5072 3606 5128
rect 3662 5072 3802 5128
rect 3601 5070 3802 5072
rect 3601 5067 3667 5070
rect 7414 5068 7420 5132
rect 7484 5130 7490 5132
rect 11053 5130 11119 5133
rect 7484 5128 11119 5130
rect 7484 5072 11058 5128
rect 11114 5072 11119 5128
rect 7484 5070 11119 5072
rect 7484 5068 7490 5070
rect 11053 5067 11119 5070
rect 20345 5130 20411 5133
rect 20621 5130 20687 5133
rect 20345 5128 20687 5130
rect 20345 5072 20350 5128
rect 20406 5072 20626 5128
rect 20682 5072 20687 5128
rect 20345 5070 20687 5072
rect 20345 5067 20411 5070
rect 20621 5067 20687 5070
rect 24209 5130 24275 5133
rect 24669 5130 24735 5133
rect 24209 5128 24735 5130
rect 24209 5072 24214 5128
rect 24270 5072 24674 5128
rect 24730 5072 24735 5128
rect 24209 5070 24735 5072
rect 24209 5067 24275 5070
rect 24669 5067 24735 5070
rect 5436 4928 5756 4929
rect 5436 4864 5444 4928
rect 5508 4864 5524 4928
rect 5588 4864 5604 4928
rect 5668 4864 5684 4928
rect 5748 4864 5756 4928
rect 5436 4863 5756 4864
rect 14422 4928 14742 4929
rect 14422 4864 14430 4928
rect 14494 4864 14510 4928
rect 14574 4864 14590 4928
rect 14654 4864 14670 4928
rect 14734 4864 14742 4928
rect 14422 4863 14742 4864
rect 23407 4928 23727 4929
rect 23407 4864 23415 4928
rect 23479 4864 23495 4928
rect 23559 4864 23575 4928
rect 23639 4864 23655 4928
rect 23719 4864 23727 4928
rect 23407 4863 23727 4864
rect 8017 4724 8083 4725
rect 7966 4660 7972 4724
rect 8036 4722 8083 4724
rect 22553 4722 22619 4725
rect 23381 4722 23447 4725
rect 8036 4720 8128 4722
rect 8078 4664 8128 4720
rect 8036 4662 8128 4664
rect 22553 4720 23447 4722
rect 22553 4664 22558 4720
rect 22614 4664 23386 4720
rect 23442 4664 23447 4720
rect 22553 4662 23447 4664
rect 8036 4660 8083 4662
rect 8017 4659 8083 4660
rect 22553 4659 22619 4662
rect 23381 4659 23447 4662
rect 3182 4388 3188 4452
rect 3252 4450 3258 4452
rect 6545 4450 6611 4453
rect 3252 4448 6611 4450
rect 3252 4392 6550 4448
rect 6606 4392 6611 4448
rect 3252 4390 6611 4392
rect 3252 4388 3258 4390
rect 6545 4387 6611 4390
rect 9929 4384 10249 4385
rect 9929 4320 9937 4384
rect 10001 4320 10017 4384
rect 10081 4320 10097 4384
rect 10161 4320 10177 4384
rect 10241 4320 10249 4384
rect 9929 4319 10249 4320
rect 18914 4384 19234 4385
rect 18914 4320 18922 4384
rect 18986 4320 19002 4384
rect 19066 4320 19082 4384
rect 19146 4320 19162 4384
rect 19226 4320 19234 4384
rect 18914 4319 19234 4320
rect 2037 4314 2103 4317
rect 2037 4312 6194 4314
rect 2037 4256 2042 4312
rect 2098 4256 6194 4312
rect 2037 4254 6194 4256
rect 2037 4251 2103 4254
rect 6134 3909 6194 4254
rect 19333 4042 19399 4045
rect 20110 4042 20116 4044
rect 19333 4040 20116 4042
rect 19333 3984 19338 4040
rect 19394 3984 20116 4040
rect 19333 3982 20116 3984
rect 19333 3979 19399 3982
rect 20110 3980 20116 3982
rect 20180 3980 20186 4044
rect 6134 3904 6243 3909
rect 6134 3848 6182 3904
rect 6238 3848 6243 3904
rect 6134 3846 6243 3848
rect 6177 3843 6243 3846
rect 19425 3906 19491 3909
rect 19926 3906 19932 3908
rect 19425 3904 19932 3906
rect 19425 3848 19430 3904
rect 19486 3848 19932 3904
rect 19425 3846 19932 3848
rect 19425 3843 19491 3846
rect 19926 3844 19932 3846
rect 19996 3844 20002 3908
rect 26233 3906 26299 3909
rect 28373 3906 29173 3936
rect 26233 3904 29173 3906
rect 26233 3848 26238 3904
rect 26294 3848 29173 3904
rect 26233 3846 29173 3848
rect 26233 3843 26299 3846
rect 5436 3840 5756 3841
rect 5436 3776 5444 3840
rect 5508 3776 5524 3840
rect 5588 3776 5604 3840
rect 5668 3776 5684 3840
rect 5748 3776 5756 3840
rect 5436 3775 5756 3776
rect 14422 3840 14742 3841
rect 14422 3776 14430 3840
rect 14494 3776 14510 3840
rect 14574 3776 14590 3840
rect 14654 3776 14670 3840
rect 14734 3776 14742 3840
rect 14422 3775 14742 3776
rect 23407 3840 23727 3841
rect 23407 3776 23415 3840
rect 23479 3776 23495 3840
rect 23559 3776 23575 3840
rect 23639 3776 23655 3840
rect 23719 3776 23727 3840
rect 28373 3816 29173 3846
rect 23407 3775 23727 3776
rect 3693 3770 3759 3773
rect 5257 3770 5323 3773
rect 3693 3768 5323 3770
rect 3693 3712 3698 3768
rect 3754 3712 5262 3768
rect 5318 3712 5323 3768
rect 3693 3710 5323 3712
rect 3693 3707 3759 3710
rect 5257 3707 5323 3710
rect 1117 3634 1183 3637
rect 5441 3634 5507 3637
rect 1117 3632 5507 3634
rect 1117 3576 1122 3632
rect 1178 3576 5446 3632
rect 5502 3576 5507 3632
rect 1117 3574 5507 3576
rect 1117 3571 1183 3574
rect 5441 3571 5507 3574
rect 105 3498 171 3501
rect 16614 3498 16620 3500
rect 105 3496 16620 3498
rect 105 3440 110 3496
rect 166 3440 16620 3496
rect 105 3438 16620 3440
rect 105 3435 171 3438
rect 16614 3436 16620 3438
rect 16684 3436 16690 3500
rect 9929 3296 10249 3297
rect 9929 3232 9937 3296
rect 10001 3232 10017 3296
rect 10081 3232 10097 3296
rect 10161 3232 10177 3296
rect 10241 3232 10249 3296
rect 9929 3231 10249 3232
rect 18914 3296 19234 3297
rect 18914 3232 18922 3296
rect 18986 3232 19002 3296
rect 19066 3232 19082 3296
rect 19146 3232 19162 3296
rect 19226 3232 19234 3296
rect 18914 3231 19234 3232
rect 2865 3226 2931 3229
rect 3325 3226 3391 3229
rect 2865 3224 3391 3226
rect 2865 3168 2870 3224
rect 2926 3168 3330 3224
rect 3386 3168 3391 3224
rect 2865 3166 3391 3168
rect 2865 3163 2931 3166
rect 3325 3163 3391 3166
rect 5257 3226 5323 3229
rect 6269 3226 6335 3229
rect 6821 3226 6887 3229
rect 5257 3224 6887 3226
rect 5257 3168 5262 3224
rect 5318 3168 6274 3224
rect 6330 3168 6826 3224
rect 6882 3168 6887 3224
rect 5257 3166 6887 3168
rect 5257 3163 5323 3166
rect 6269 3163 6335 3166
rect 6821 3163 6887 3166
rect 18638 3164 18644 3228
rect 18708 3226 18714 3228
rect 18781 3226 18847 3229
rect 18708 3224 18847 3226
rect 18708 3168 18786 3224
rect 18842 3168 18847 3224
rect 18708 3166 18847 3168
rect 18708 3164 18714 3166
rect 18781 3163 18847 3166
rect 4102 3028 4108 3092
rect 4172 3090 4178 3092
rect 12617 3090 12683 3093
rect 4172 3088 12683 3090
rect 4172 3032 12622 3088
rect 12678 3032 12683 3088
rect 4172 3030 12683 3032
rect 4172 3028 4178 3030
rect 12617 3027 12683 3030
rect 7005 2954 7071 2957
rect 7373 2954 7439 2957
rect 7005 2952 7439 2954
rect 7005 2896 7010 2952
rect 7066 2896 7378 2952
rect 7434 2896 7439 2952
rect 7005 2894 7439 2896
rect 7005 2891 7071 2894
rect 7373 2891 7439 2894
rect 20069 2954 20135 2957
rect 20989 2954 21055 2957
rect 20069 2952 21055 2954
rect 20069 2896 20074 2952
rect 20130 2896 20994 2952
rect 21050 2896 21055 2952
rect 20069 2894 21055 2896
rect 20069 2891 20135 2894
rect 20989 2891 21055 2894
rect 1301 2818 1367 2821
rect 11053 2818 11119 2821
rect 12157 2818 12223 2821
rect 1301 2816 5274 2818
rect 1301 2760 1306 2816
rect 1362 2760 5274 2816
rect 1301 2758 5274 2760
rect 1301 2755 1367 2758
rect 5214 2546 5274 2758
rect 11053 2816 12223 2818
rect 11053 2760 11058 2816
rect 11114 2760 12162 2816
rect 12218 2760 12223 2816
rect 11053 2758 12223 2760
rect 11053 2755 11119 2758
rect 12157 2755 12223 2758
rect 5436 2752 5756 2753
rect 5436 2688 5444 2752
rect 5508 2688 5524 2752
rect 5588 2688 5604 2752
rect 5668 2688 5684 2752
rect 5748 2688 5756 2752
rect 5436 2687 5756 2688
rect 14422 2752 14742 2753
rect 14422 2688 14430 2752
rect 14494 2688 14510 2752
rect 14574 2688 14590 2752
rect 14654 2688 14670 2752
rect 14734 2688 14742 2752
rect 14422 2687 14742 2688
rect 23407 2752 23727 2753
rect 23407 2688 23415 2752
rect 23479 2688 23495 2752
rect 23559 2688 23575 2752
rect 23639 2688 23655 2752
rect 23719 2688 23727 2752
rect 23407 2687 23727 2688
rect 5717 2546 5783 2549
rect 5214 2544 5783 2546
rect 5214 2488 5722 2544
rect 5778 2488 5783 2544
rect 5214 2486 5783 2488
rect 5717 2483 5783 2486
rect 10961 2546 11027 2549
rect 12198 2546 12204 2548
rect 10961 2544 12204 2546
rect 10961 2488 10966 2544
rect 11022 2488 12204 2544
rect 10961 2486 12204 2488
rect 10961 2483 11027 2486
rect 12198 2484 12204 2486
rect 12268 2484 12274 2548
rect 9929 2208 10249 2209
rect 9929 2144 9937 2208
rect 10001 2144 10017 2208
rect 10081 2144 10097 2208
rect 10161 2144 10177 2208
rect 10241 2144 10249 2208
rect 9929 2143 10249 2144
rect 18914 2208 19234 2209
rect 18914 2144 18922 2208
rect 18986 2144 19002 2208
rect 19066 2144 19082 2208
rect 19146 2144 19162 2208
rect 19226 2144 19234 2208
rect 18914 2143 19234 2144
<< via3 >>
rect 5444 28860 5508 28864
rect 5444 28804 5448 28860
rect 5448 28804 5504 28860
rect 5504 28804 5508 28860
rect 5444 28800 5508 28804
rect 5524 28860 5588 28864
rect 5524 28804 5528 28860
rect 5528 28804 5584 28860
rect 5584 28804 5588 28860
rect 5524 28800 5588 28804
rect 5604 28860 5668 28864
rect 5604 28804 5608 28860
rect 5608 28804 5664 28860
rect 5664 28804 5668 28860
rect 5604 28800 5668 28804
rect 5684 28860 5748 28864
rect 5684 28804 5688 28860
rect 5688 28804 5744 28860
rect 5744 28804 5748 28860
rect 5684 28800 5748 28804
rect 14430 28860 14494 28864
rect 14430 28804 14434 28860
rect 14434 28804 14490 28860
rect 14490 28804 14494 28860
rect 14430 28800 14494 28804
rect 14510 28860 14574 28864
rect 14510 28804 14514 28860
rect 14514 28804 14570 28860
rect 14570 28804 14574 28860
rect 14510 28800 14574 28804
rect 14590 28860 14654 28864
rect 14590 28804 14594 28860
rect 14594 28804 14650 28860
rect 14650 28804 14654 28860
rect 14590 28800 14654 28804
rect 14670 28860 14734 28864
rect 14670 28804 14674 28860
rect 14674 28804 14730 28860
rect 14730 28804 14734 28860
rect 14670 28800 14734 28804
rect 23415 28860 23479 28864
rect 23415 28804 23419 28860
rect 23419 28804 23475 28860
rect 23475 28804 23479 28860
rect 23415 28800 23479 28804
rect 23495 28860 23559 28864
rect 23495 28804 23499 28860
rect 23499 28804 23555 28860
rect 23555 28804 23559 28860
rect 23495 28800 23559 28804
rect 23575 28860 23639 28864
rect 23575 28804 23579 28860
rect 23579 28804 23635 28860
rect 23635 28804 23639 28860
rect 23575 28800 23639 28804
rect 23655 28860 23719 28864
rect 23655 28804 23659 28860
rect 23659 28804 23715 28860
rect 23715 28804 23719 28860
rect 23655 28800 23719 28804
rect 9937 28316 10001 28320
rect 9937 28260 9941 28316
rect 9941 28260 9997 28316
rect 9997 28260 10001 28316
rect 9937 28256 10001 28260
rect 10017 28316 10081 28320
rect 10017 28260 10021 28316
rect 10021 28260 10077 28316
rect 10077 28260 10081 28316
rect 10017 28256 10081 28260
rect 10097 28316 10161 28320
rect 10097 28260 10101 28316
rect 10101 28260 10157 28316
rect 10157 28260 10161 28316
rect 10097 28256 10161 28260
rect 10177 28316 10241 28320
rect 10177 28260 10181 28316
rect 10181 28260 10237 28316
rect 10237 28260 10241 28316
rect 10177 28256 10241 28260
rect 18922 28316 18986 28320
rect 18922 28260 18926 28316
rect 18926 28260 18982 28316
rect 18982 28260 18986 28316
rect 18922 28256 18986 28260
rect 19002 28316 19066 28320
rect 19002 28260 19006 28316
rect 19006 28260 19062 28316
rect 19062 28260 19066 28316
rect 19002 28256 19066 28260
rect 19082 28316 19146 28320
rect 19082 28260 19086 28316
rect 19086 28260 19142 28316
rect 19142 28260 19146 28316
rect 19082 28256 19146 28260
rect 19162 28316 19226 28320
rect 19162 28260 19166 28316
rect 19166 28260 19222 28316
rect 19222 28260 19226 28316
rect 19162 28256 19226 28260
rect 14228 27916 14292 27980
rect 5444 27772 5508 27776
rect 5444 27716 5448 27772
rect 5448 27716 5504 27772
rect 5504 27716 5508 27772
rect 5444 27712 5508 27716
rect 5524 27772 5588 27776
rect 5524 27716 5528 27772
rect 5528 27716 5584 27772
rect 5584 27716 5588 27772
rect 5524 27712 5588 27716
rect 5604 27772 5668 27776
rect 5604 27716 5608 27772
rect 5608 27716 5664 27772
rect 5664 27716 5668 27772
rect 5604 27712 5668 27716
rect 5684 27772 5748 27776
rect 5684 27716 5688 27772
rect 5688 27716 5744 27772
rect 5744 27716 5748 27772
rect 5684 27712 5748 27716
rect 14430 27772 14494 27776
rect 14430 27716 14434 27772
rect 14434 27716 14490 27772
rect 14490 27716 14494 27772
rect 14430 27712 14494 27716
rect 14510 27772 14574 27776
rect 14510 27716 14514 27772
rect 14514 27716 14570 27772
rect 14570 27716 14574 27772
rect 14510 27712 14574 27716
rect 14590 27772 14654 27776
rect 14590 27716 14594 27772
rect 14594 27716 14650 27772
rect 14650 27716 14654 27772
rect 14590 27712 14654 27716
rect 14670 27772 14734 27776
rect 14670 27716 14674 27772
rect 14674 27716 14730 27772
rect 14730 27716 14734 27772
rect 14670 27712 14734 27716
rect 23415 27772 23479 27776
rect 23415 27716 23419 27772
rect 23419 27716 23475 27772
rect 23475 27716 23479 27772
rect 23415 27712 23479 27716
rect 23495 27772 23559 27776
rect 23495 27716 23499 27772
rect 23499 27716 23555 27772
rect 23555 27716 23559 27772
rect 23495 27712 23559 27716
rect 23575 27772 23639 27776
rect 23575 27716 23579 27772
rect 23579 27716 23635 27772
rect 23635 27716 23639 27772
rect 23575 27712 23639 27716
rect 23655 27772 23719 27776
rect 23655 27716 23659 27772
rect 23659 27716 23715 27772
rect 23715 27716 23719 27772
rect 23655 27712 23719 27716
rect 12204 27704 12268 27708
rect 12204 27648 12218 27704
rect 12218 27648 12268 27704
rect 12204 27644 12268 27648
rect 23796 27704 23860 27708
rect 23796 27648 23846 27704
rect 23846 27648 23860 27704
rect 23796 27644 23860 27648
rect 9937 27228 10001 27232
rect 9937 27172 9941 27228
rect 9941 27172 9997 27228
rect 9997 27172 10001 27228
rect 9937 27168 10001 27172
rect 10017 27228 10081 27232
rect 10017 27172 10021 27228
rect 10021 27172 10077 27228
rect 10077 27172 10081 27228
rect 10017 27168 10081 27172
rect 10097 27228 10161 27232
rect 10097 27172 10101 27228
rect 10101 27172 10157 27228
rect 10157 27172 10161 27228
rect 10097 27168 10161 27172
rect 10177 27228 10241 27232
rect 10177 27172 10181 27228
rect 10181 27172 10237 27228
rect 10237 27172 10241 27228
rect 10177 27168 10241 27172
rect 18922 27228 18986 27232
rect 18922 27172 18926 27228
rect 18926 27172 18982 27228
rect 18982 27172 18986 27228
rect 18922 27168 18986 27172
rect 19002 27228 19066 27232
rect 19002 27172 19006 27228
rect 19006 27172 19062 27228
rect 19062 27172 19066 27228
rect 19002 27168 19066 27172
rect 19082 27228 19146 27232
rect 19082 27172 19086 27228
rect 19086 27172 19142 27228
rect 19142 27172 19146 27228
rect 19082 27168 19146 27172
rect 19162 27228 19226 27232
rect 19162 27172 19166 27228
rect 19166 27172 19222 27228
rect 19222 27172 19226 27228
rect 19162 27168 19226 27172
rect 6500 26828 6564 26892
rect 5444 26684 5508 26688
rect 5444 26628 5448 26684
rect 5448 26628 5504 26684
rect 5504 26628 5508 26684
rect 5444 26624 5508 26628
rect 5524 26684 5588 26688
rect 5524 26628 5528 26684
rect 5528 26628 5584 26684
rect 5584 26628 5588 26684
rect 5524 26624 5588 26628
rect 5604 26684 5668 26688
rect 5604 26628 5608 26684
rect 5608 26628 5664 26684
rect 5664 26628 5668 26684
rect 5604 26624 5668 26628
rect 5684 26684 5748 26688
rect 5684 26628 5688 26684
rect 5688 26628 5744 26684
rect 5744 26628 5748 26684
rect 5684 26624 5748 26628
rect 14430 26684 14494 26688
rect 14430 26628 14434 26684
rect 14434 26628 14490 26684
rect 14490 26628 14494 26684
rect 14430 26624 14494 26628
rect 14510 26684 14574 26688
rect 14510 26628 14514 26684
rect 14514 26628 14570 26684
rect 14570 26628 14574 26684
rect 14510 26624 14574 26628
rect 14590 26684 14654 26688
rect 14590 26628 14594 26684
rect 14594 26628 14650 26684
rect 14650 26628 14654 26684
rect 14590 26624 14654 26628
rect 14670 26684 14734 26688
rect 14670 26628 14674 26684
rect 14674 26628 14730 26684
rect 14730 26628 14734 26684
rect 14670 26624 14734 26628
rect 23415 26684 23479 26688
rect 23415 26628 23419 26684
rect 23419 26628 23475 26684
rect 23475 26628 23479 26684
rect 23415 26624 23479 26628
rect 23495 26684 23559 26688
rect 23495 26628 23499 26684
rect 23499 26628 23555 26684
rect 23555 26628 23559 26684
rect 23495 26624 23559 26628
rect 23575 26684 23639 26688
rect 23575 26628 23579 26684
rect 23579 26628 23635 26684
rect 23635 26628 23639 26684
rect 23575 26624 23639 26628
rect 23655 26684 23719 26688
rect 23655 26628 23659 26684
rect 23659 26628 23715 26684
rect 23715 26628 23719 26684
rect 23655 26624 23719 26628
rect 11468 26420 11532 26484
rect 3372 26284 3436 26348
rect 15332 26284 15396 26348
rect 18276 26284 18340 26348
rect 19564 26284 19628 26348
rect 23244 26344 23308 26348
rect 23244 26288 23258 26344
rect 23258 26288 23308 26344
rect 23244 26284 23308 26288
rect 9937 26140 10001 26144
rect 9937 26084 9941 26140
rect 9941 26084 9997 26140
rect 9997 26084 10001 26140
rect 9937 26080 10001 26084
rect 10017 26140 10081 26144
rect 10017 26084 10021 26140
rect 10021 26084 10077 26140
rect 10077 26084 10081 26140
rect 10017 26080 10081 26084
rect 10097 26140 10161 26144
rect 10097 26084 10101 26140
rect 10101 26084 10157 26140
rect 10157 26084 10161 26140
rect 10097 26080 10161 26084
rect 10177 26140 10241 26144
rect 10177 26084 10181 26140
rect 10181 26084 10237 26140
rect 10237 26084 10241 26140
rect 10177 26080 10241 26084
rect 18922 26140 18986 26144
rect 18922 26084 18926 26140
rect 18926 26084 18982 26140
rect 18982 26084 18986 26140
rect 18922 26080 18986 26084
rect 19002 26140 19066 26144
rect 19002 26084 19006 26140
rect 19006 26084 19062 26140
rect 19062 26084 19066 26140
rect 19002 26080 19066 26084
rect 19082 26140 19146 26144
rect 19082 26084 19086 26140
rect 19086 26084 19142 26140
rect 19142 26084 19146 26140
rect 19082 26080 19146 26084
rect 19162 26140 19226 26144
rect 19162 26084 19166 26140
rect 19166 26084 19222 26140
rect 19222 26084 19226 26140
rect 19162 26080 19226 26084
rect 5444 25596 5508 25600
rect 5444 25540 5448 25596
rect 5448 25540 5504 25596
rect 5504 25540 5508 25596
rect 5444 25536 5508 25540
rect 5524 25596 5588 25600
rect 5524 25540 5528 25596
rect 5528 25540 5584 25596
rect 5584 25540 5588 25596
rect 5524 25536 5588 25540
rect 5604 25596 5668 25600
rect 5604 25540 5608 25596
rect 5608 25540 5664 25596
rect 5664 25540 5668 25596
rect 5604 25536 5668 25540
rect 5684 25596 5748 25600
rect 5684 25540 5688 25596
rect 5688 25540 5744 25596
rect 5744 25540 5748 25596
rect 5684 25536 5748 25540
rect 14430 25596 14494 25600
rect 14430 25540 14434 25596
rect 14434 25540 14490 25596
rect 14490 25540 14494 25596
rect 14430 25536 14494 25540
rect 14510 25596 14574 25600
rect 14510 25540 14514 25596
rect 14514 25540 14570 25596
rect 14570 25540 14574 25596
rect 14510 25536 14574 25540
rect 14590 25596 14654 25600
rect 14590 25540 14594 25596
rect 14594 25540 14650 25596
rect 14650 25540 14654 25596
rect 14590 25536 14654 25540
rect 14670 25596 14734 25600
rect 14670 25540 14674 25596
rect 14674 25540 14730 25596
rect 14730 25540 14734 25596
rect 14670 25536 14734 25540
rect 23415 25596 23479 25600
rect 23415 25540 23419 25596
rect 23419 25540 23475 25596
rect 23475 25540 23479 25596
rect 23415 25536 23479 25540
rect 23495 25596 23559 25600
rect 23495 25540 23499 25596
rect 23499 25540 23555 25596
rect 23555 25540 23559 25596
rect 23495 25536 23559 25540
rect 23575 25596 23639 25600
rect 23575 25540 23579 25596
rect 23579 25540 23635 25596
rect 23635 25540 23639 25596
rect 23575 25536 23639 25540
rect 23655 25596 23719 25600
rect 23655 25540 23659 25596
rect 23659 25540 23715 25596
rect 23715 25540 23719 25596
rect 23655 25536 23719 25540
rect 27476 25332 27540 25396
rect 25084 25060 25148 25124
rect 9937 25052 10001 25056
rect 9937 24996 9941 25052
rect 9941 24996 9997 25052
rect 9997 24996 10001 25052
rect 9937 24992 10001 24996
rect 10017 25052 10081 25056
rect 10017 24996 10021 25052
rect 10021 24996 10077 25052
rect 10077 24996 10081 25052
rect 10017 24992 10081 24996
rect 10097 25052 10161 25056
rect 10097 24996 10101 25052
rect 10101 24996 10157 25052
rect 10157 24996 10161 25052
rect 10097 24992 10161 24996
rect 10177 25052 10241 25056
rect 10177 24996 10181 25052
rect 10181 24996 10237 25052
rect 10237 24996 10241 25052
rect 10177 24992 10241 24996
rect 18922 25052 18986 25056
rect 18922 24996 18926 25052
rect 18926 24996 18982 25052
rect 18982 24996 18986 25052
rect 18922 24992 18986 24996
rect 19002 25052 19066 25056
rect 19002 24996 19006 25052
rect 19006 24996 19062 25052
rect 19062 24996 19066 25052
rect 19002 24992 19066 24996
rect 19082 25052 19146 25056
rect 19082 24996 19086 25052
rect 19086 24996 19142 25052
rect 19142 24996 19146 25052
rect 19082 24992 19146 24996
rect 19162 25052 19226 25056
rect 19162 24996 19166 25052
rect 19166 24996 19222 25052
rect 19222 24996 19226 25052
rect 19162 24992 19226 24996
rect 25268 24924 25332 24988
rect 15700 24788 15764 24852
rect 5444 24508 5508 24512
rect 5444 24452 5448 24508
rect 5448 24452 5504 24508
rect 5504 24452 5508 24508
rect 5444 24448 5508 24452
rect 5524 24508 5588 24512
rect 5524 24452 5528 24508
rect 5528 24452 5584 24508
rect 5584 24452 5588 24508
rect 5524 24448 5588 24452
rect 5604 24508 5668 24512
rect 5604 24452 5608 24508
rect 5608 24452 5664 24508
rect 5664 24452 5668 24508
rect 5604 24448 5668 24452
rect 5684 24508 5748 24512
rect 5684 24452 5688 24508
rect 5688 24452 5744 24508
rect 5744 24452 5748 24508
rect 5684 24448 5748 24452
rect 14430 24508 14494 24512
rect 14430 24452 14434 24508
rect 14434 24452 14490 24508
rect 14490 24452 14494 24508
rect 14430 24448 14494 24452
rect 14510 24508 14574 24512
rect 14510 24452 14514 24508
rect 14514 24452 14570 24508
rect 14570 24452 14574 24508
rect 14510 24448 14574 24452
rect 14590 24508 14654 24512
rect 14590 24452 14594 24508
rect 14594 24452 14650 24508
rect 14650 24452 14654 24508
rect 14590 24448 14654 24452
rect 14670 24508 14734 24512
rect 14670 24452 14674 24508
rect 14674 24452 14730 24508
rect 14730 24452 14734 24508
rect 14670 24448 14734 24452
rect 23415 24508 23479 24512
rect 23415 24452 23419 24508
rect 23419 24452 23475 24508
rect 23475 24452 23479 24508
rect 23415 24448 23479 24452
rect 23495 24508 23559 24512
rect 23495 24452 23499 24508
rect 23499 24452 23555 24508
rect 23555 24452 23559 24508
rect 23495 24448 23559 24452
rect 23575 24508 23639 24512
rect 23575 24452 23579 24508
rect 23579 24452 23635 24508
rect 23635 24452 23639 24508
rect 23575 24448 23639 24452
rect 23655 24508 23719 24512
rect 23655 24452 23659 24508
rect 23659 24452 23715 24508
rect 23715 24452 23719 24508
rect 23655 24448 23719 24452
rect 22692 23972 22756 24036
rect 9937 23964 10001 23968
rect 9937 23908 9941 23964
rect 9941 23908 9997 23964
rect 9997 23908 10001 23964
rect 9937 23904 10001 23908
rect 10017 23964 10081 23968
rect 10017 23908 10021 23964
rect 10021 23908 10077 23964
rect 10077 23908 10081 23964
rect 10017 23904 10081 23908
rect 10097 23964 10161 23968
rect 10097 23908 10101 23964
rect 10101 23908 10157 23964
rect 10157 23908 10161 23964
rect 10097 23904 10161 23908
rect 10177 23964 10241 23968
rect 10177 23908 10181 23964
rect 10181 23908 10237 23964
rect 10237 23908 10241 23964
rect 10177 23904 10241 23908
rect 18922 23964 18986 23968
rect 18922 23908 18926 23964
rect 18926 23908 18982 23964
rect 18982 23908 18986 23964
rect 18922 23904 18986 23908
rect 19002 23964 19066 23968
rect 19002 23908 19006 23964
rect 19006 23908 19062 23964
rect 19062 23908 19066 23964
rect 19002 23904 19066 23908
rect 19082 23964 19146 23968
rect 19082 23908 19086 23964
rect 19086 23908 19142 23964
rect 19142 23908 19146 23964
rect 19082 23904 19146 23908
rect 19162 23964 19226 23968
rect 19162 23908 19166 23964
rect 19166 23908 19222 23964
rect 19222 23908 19226 23964
rect 19162 23904 19226 23908
rect 23980 23700 24044 23764
rect 21220 23428 21284 23492
rect 22324 23488 22388 23492
rect 22324 23432 22338 23488
rect 22338 23432 22388 23488
rect 22324 23428 22388 23432
rect 5444 23420 5508 23424
rect 5444 23364 5448 23420
rect 5448 23364 5504 23420
rect 5504 23364 5508 23420
rect 5444 23360 5508 23364
rect 5524 23420 5588 23424
rect 5524 23364 5528 23420
rect 5528 23364 5584 23420
rect 5584 23364 5588 23420
rect 5524 23360 5588 23364
rect 5604 23420 5668 23424
rect 5604 23364 5608 23420
rect 5608 23364 5664 23420
rect 5664 23364 5668 23420
rect 5604 23360 5668 23364
rect 5684 23420 5748 23424
rect 5684 23364 5688 23420
rect 5688 23364 5744 23420
rect 5744 23364 5748 23420
rect 5684 23360 5748 23364
rect 14430 23420 14494 23424
rect 14430 23364 14434 23420
rect 14434 23364 14490 23420
rect 14490 23364 14494 23420
rect 14430 23360 14494 23364
rect 14510 23420 14574 23424
rect 14510 23364 14514 23420
rect 14514 23364 14570 23420
rect 14570 23364 14574 23420
rect 14510 23360 14574 23364
rect 14590 23420 14654 23424
rect 14590 23364 14594 23420
rect 14594 23364 14650 23420
rect 14650 23364 14654 23420
rect 14590 23360 14654 23364
rect 14670 23420 14734 23424
rect 14670 23364 14674 23420
rect 14674 23364 14730 23420
rect 14730 23364 14734 23420
rect 14670 23360 14734 23364
rect 23415 23420 23479 23424
rect 23415 23364 23419 23420
rect 23419 23364 23475 23420
rect 23475 23364 23479 23420
rect 23415 23360 23479 23364
rect 23495 23420 23559 23424
rect 23495 23364 23499 23420
rect 23499 23364 23555 23420
rect 23555 23364 23559 23420
rect 23495 23360 23559 23364
rect 23575 23420 23639 23424
rect 23575 23364 23579 23420
rect 23579 23364 23635 23420
rect 23635 23364 23639 23420
rect 23575 23360 23639 23364
rect 23655 23420 23719 23424
rect 23655 23364 23659 23420
rect 23659 23364 23715 23420
rect 23715 23364 23719 23420
rect 23655 23360 23719 23364
rect 4476 22884 4540 22948
rect 20484 23020 20548 23084
rect 23244 23156 23308 23220
rect 9937 22876 10001 22880
rect 9937 22820 9941 22876
rect 9941 22820 9997 22876
rect 9997 22820 10001 22876
rect 9937 22816 10001 22820
rect 10017 22876 10081 22880
rect 10017 22820 10021 22876
rect 10021 22820 10077 22876
rect 10077 22820 10081 22876
rect 10017 22816 10081 22820
rect 10097 22876 10161 22880
rect 10097 22820 10101 22876
rect 10101 22820 10157 22876
rect 10157 22820 10161 22876
rect 10097 22816 10161 22820
rect 10177 22876 10241 22880
rect 10177 22820 10181 22876
rect 10181 22820 10237 22876
rect 10237 22820 10241 22876
rect 10177 22816 10241 22820
rect 18922 22876 18986 22880
rect 18922 22820 18926 22876
rect 18926 22820 18982 22876
rect 18982 22820 18986 22876
rect 18922 22816 18986 22820
rect 19002 22876 19066 22880
rect 19002 22820 19006 22876
rect 19006 22820 19062 22876
rect 19062 22820 19066 22876
rect 19002 22816 19066 22820
rect 19082 22876 19146 22880
rect 19082 22820 19086 22876
rect 19086 22820 19142 22876
rect 19142 22820 19146 22876
rect 19082 22816 19146 22820
rect 19162 22876 19226 22880
rect 19162 22820 19166 22876
rect 19166 22820 19222 22876
rect 19222 22820 19226 22876
rect 19162 22816 19226 22820
rect 4108 22672 4172 22676
rect 4108 22616 4158 22672
rect 4158 22616 4172 22672
rect 4108 22612 4172 22616
rect 4844 22536 4908 22540
rect 4844 22480 4894 22536
rect 4894 22480 4908 22536
rect 4844 22476 4908 22480
rect 5212 22536 5276 22540
rect 5212 22480 5262 22536
rect 5262 22480 5276 22536
rect 5212 22476 5276 22480
rect 5444 22332 5508 22336
rect 5444 22276 5448 22332
rect 5448 22276 5504 22332
rect 5504 22276 5508 22332
rect 5444 22272 5508 22276
rect 5524 22332 5588 22336
rect 5524 22276 5528 22332
rect 5528 22276 5584 22332
rect 5584 22276 5588 22332
rect 5524 22272 5588 22276
rect 5604 22332 5668 22336
rect 5604 22276 5608 22332
rect 5608 22276 5664 22332
rect 5664 22276 5668 22332
rect 5604 22272 5668 22276
rect 5684 22332 5748 22336
rect 5684 22276 5688 22332
rect 5688 22276 5744 22332
rect 5744 22276 5748 22332
rect 5684 22272 5748 22276
rect 14430 22332 14494 22336
rect 14430 22276 14434 22332
rect 14434 22276 14490 22332
rect 14490 22276 14494 22332
rect 14430 22272 14494 22276
rect 14510 22332 14574 22336
rect 14510 22276 14514 22332
rect 14514 22276 14570 22332
rect 14570 22276 14574 22332
rect 14510 22272 14574 22276
rect 14590 22332 14654 22336
rect 14590 22276 14594 22332
rect 14594 22276 14650 22332
rect 14650 22276 14654 22332
rect 14590 22272 14654 22276
rect 14670 22332 14734 22336
rect 14670 22276 14674 22332
rect 14674 22276 14730 22332
rect 14730 22276 14734 22332
rect 14670 22272 14734 22276
rect 22508 22884 22572 22948
rect 23415 22332 23479 22336
rect 23415 22276 23419 22332
rect 23419 22276 23475 22332
rect 23475 22276 23479 22332
rect 23415 22272 23479 22276
rect 23495 22332 23559 22336
rect 23495 22276 23499 22332
rect 23499 22276 23555 22332
rect 23555 22276 23559 22332
rect 23495 22272 23559 22276
rect 23575 22332 23639 22336
rect 23575 22276 23579 22332
rect 23579 22276 23635 22332
rect 23635 22276 23639 22332
rect 23575 22272 23639 22276
rect 23655 22332 23719 22336
rect 23655 22276 23659 22332
rect 23659 22276 23715 22332
rect 23715 22276 23719 22332
rect 23655 22272 23719 22276
rect 6316 21796 6380 21860
rect 18276 21856 18340 21860
rect 18276 21800 18290 21856
rect 18290 21800 18340 21856
rect 18276 21796 18340 21800
rect 9937 21788 10001 21792
rect 9937 21732 9941 21788
rect 9941 21732 9997 21788
rect 9997 21732 10001 21788
rect 9937 21728 10001 21732
rect 10017 21788 10081 21792
rect 10017 21732 10021 21788
rect 10021 21732 10077 21788
rect 10077 21732 10081 21788
rect 10017 21728 10081 21732
rect 10097 21788 10161 21792
rect 10097 21732 10101 21788
rect 10101 21732 10157 21788
rect 10157 21732 10161 21788
rect 10097 21728 10161 21732
rect 10177 21788 10241 21792
rect 10177 21732 10181 21788
rect 10181 21732 10237 21788
rect 10237 21732 10241 21788
rect 10177 21728 10241 21732
rect 18922 21788 18986 21792
rect 18922 21732 18926 21788
rect 18926 21732 18982 21788
rect 18982 21732 18986 21788
rect 18922 21728 18986 21732
rect 19002 21788 19066 21792
rect 19002 21732 19006 21788
rect 19006 21732 19062 21788
rect 19062 21732 19066 21788
rect 19002 21728 19066 21732
rect 19082 21788 19146 21792
rect 19082 21732 19086 21788
rect 19086 21732 19142 21788
rect 19142 21732 19146 21788
rect 19082 21728 19146 21732
rect 19162 21788 19226 21792
rect 19162 21732 19166 21788
rect 19166 21732 19222 21788
rect 19222 21732 19226 21788
rect 19162 21728 19226 21732
rect 5212 21388 5276 21452
rect 7236 21388 7300 21452
rect 14964 21448 15028 21452
rect 14964 21392 15014 21448
rect 15014 21392 15028 21448
rect 14964 21388 15028 21392
rect 5212 21252 5276 21316
rect 5444 21244 5508 21248
rect 5444 21188 5448 21244
rect 5448 21188 5504 21244
rect 5504 21188 5508 21244
rect 5444 21184 5508 21188
rect 5524 21244 5588 21248
rect 5524 21188 5528 21244
rect 5528 21188 5584 21244
rect 5584 21188 5588 21244
rect 5524 21184 5588 21188
rect 5604 21244 5668 21248
rect 5604 21188 5608 21244
rect 5608 21188 5664 21244
rect 5664 21188 5668 21244
rect 5604 21184 5668 21188
rect 5684 21244 5748 21248
rect 5684 21188 5688 21244
rect 5688 21188 5744 21244
rect 5744 21188 5748 21244
rect 5684 21184 5748 21188
rect 14430 21244 14494 21248
rect 14430 21188 14434 21244
rect 14434 21188 14490 21244
rect 14490 21188 14494 21244
rect 14430 21184 14494 21188
rect 14510 21244 14574 21248
rect 14510 21188 14514 21244
rect 14514 21188 14570 21244
rect 14570 21188 14574 21244
rect 14510 21184 14574 21188
rect 14590 21244 14654 21248
rect 14590 21188 14594 21244
rect 14594 21188 14650 21244
rect 14650 21188 14654 21244
rect 14590 21184 14654 21188
rect 14670 21244 14734 21248
rect 14670 21188 14674 21244
rect 14674 21188 14730 21244
rect 14730 21188 14734 21244
rect 14670 21184 14734 21188
rect 23415 21244 23479 21248
rect 23415 21188 23419 21244
rect 23419 21188 23475 21244
rect 23475 21188 23479 21244
rect 23415 21184 23479 21188
rect 23495 21244 23559 21248
rect 23495 21188 23499 21244
rect 23499 21188 23555 21244
rect 23555 21188 23559 21244
rect 23495 21184 23559 21188
rect 23575 21244 23639 21248
rect 23575 21188 23579 21244
rect 23579 21188 23635 21244
rect 23635 21188 23639 21244
rect 23575 21184 23639 21188
rect 23655 21244 23719 21248
rect 23655 21188 23659 21244
rect 23659 21188 23715 21244
rect 23715 21188 23719 21244
rect 23655 21184 23719 21188
rect 6132 20980 6196 21044
rect 13676 20980 13740 21044
rect 14044 21040 14108 21044
rect 14044 20984 14058 21040
rect 14058 20984 14108 21040
rect 14044 20980 14108 20984
rect 9628 20844 9692 20908
rect 11284 20844 11348 20908
rect 9260 20708 9324 20772
rect 21956 20708 22020 20772
rect 22140 20708 22204 20772
rect 9937 20700 10001 20704
rect 9937 20644 9941 20700
rect 9941 20644 9997 20700
rect 9997 20644 10001 20700
rect 9937 20640 10001 20644
rect 10017 20700 10081 20704
rect 10017 20644 10021 20700
rect 10021 20644 10077 20700
rect 10077 20644 10081 20700
rect 10017 20640 10081 20644
rect 10097 20700 10161 20704
rect 10097 20644 10101 20700
rect 10101 20644 10157 20700
rect 10157 20644 10161 20700
rect 10097 20640 10161 20644
rect 10177 20700 10241 20704
rect 10177 20644 10181 20700
rect 10181 20644 10237 20700
rect 10237 20644 10241 20700
rect 10177 20640 10241 20644
rect 18922 20700 18986 20704
rect 18922 20644 18926 20700
rect 18926 20644 18982 20700
rect 18982 20644 18986 20700
rect 18922 20640 18986 20644
rect 19002 20700 19066 20704
rect 19002 20644 19006 20700
rect 19006 20644 19062 20700
rect 19062 20644 19066 20700
rect 19002 20640 19066 20644
rect 19082 20700 19146 20704
rect 19082 20644 19086 20700
rect 19086 20644 19142 20700
rect 19142 20644 19146 20700
rect 19082 20640 19146 20644
rect 19162 20700 19226 20704
rect 19162 20644 19166 20700
rect 19166 20644 19222 20700
rect 19222 20644 19226 20700
rect 19162 20640 19226 20644
rect 4844 20572 4908 20636
rect 7972 20436 8036 20500
rect 3556 20360 3620 20364
rect 3556 20304 3606 20360
rect 3606 20304 3620 20360
rect 3556 20300 3620 20304
rect 5444 20156 5508 20160
rect 5444 20100 5448 20156
rect 5448 20100 5504 20156
rect 5504 20100 5508 20156
rect 5444 20096 5508 20100
rect 5524 20156 5588 20160
rect 5524 20100 5528 20156
rect 5528 20100 5584 20156
rect 5584 20100 5588 20156
rect 5524 20096 5588 20100
rect 5604 20156 5668 20160
rect 5604 20100 5608 20156
rect 5608 20100 5664 20156
rect 5664 20100 5668 20156
rect 5604 20096 5668 20100
rect 5684 20156 5748 20160
rect 5684 20100 5688 20156
rect 5688 20100 5744 20156
rect 5744 20100 5748 20156
rect 5684 20096 5748 20100
rect 14430 20156 14494 20160
rect 14430 20100 14434 20156
rect 14434 20100 14490 20156
rect 14490 20100 14494 20156
rect 14430 20096 14494 20100
rect 14510 20156 14574 20160
rect 14510 20100 14514 20156
rect 14514 20100 14570 20156
rect 14570 20100 14574 20156
rect 14510 20096 14574 20100
rect 14590 20156 14654 20160
rect 14590 20100 14594 20156
rect 14594 20100 14650 20156
rect 14650 20100 14654 20156
rect 14590 20096 14654 20100
rect 14670 20156 14734 20160
rect 14670 20100 14674 20156
rect 14674 20100 14730 20156
rect 14730 20100 14734 20156
rect 14670 20096 14734 20100
rect 23415 20156 23479 20160
rect 23415 20100 23419 20156
rect 23419 20100 23475 20156
rect 23475 20100 23479 20156
rect 23415 20096 23479 20100
rect 23495 20156 23559 20160
rect 23495 20100 23499 20156
rect 23499 20100 23555 20156
rect 23555 20100 23559 20156
rect 23495 20096 23559 20100
rect 23575 20156 23639 20160
rect 23575 20100 23579 20156
rect 23579 20100 23635 20156
rect 23635 20100 23639 20156
rect 23575 20096 23639 20100
rect 23655 20156 23719 20160
rect 23655 20100 23659 20156
rect 23659 20100 23715 20156
rect 23715 20100 23719 20156
rect 23655 20096 23719 20100
rect 13492 20028 13556 20092
rect 7788 19892 7852 19956
rect 8156 19952 8220 19956
rect 8156 19896 8170 19952
rect 8170 19896 8220 19952
rect 8156 19892 8220 19896
rect 15884 19952 15948 19956
rect 15884 19896 15934 19952
rect 15934 19896 15948 19952
rect 15884 19892 15948 19896
rect 18460 19892 18524 19956
rect 5948 19620 6012 19684
rect 16436 19756 16500 19820
rect 15148 19620 15212 19684
rect 9937 19612 10001 19616
rect 9937 19556 9941 19612
rect 9941 19556 9997 19612
rect 9997 19556 10001 19612
rect 9937 19552 10001 19556
rect 10017 19612 10081 19616
rect 10017 19556 10021 19612
rect 10021 19556 10077 19612
rect 10077 19556 10081 19612
rect 10017 19552 10081 19556
rect 10097 19612 10161 19616
rect 10097 19556 10101 19612
rect 10101 19556 10157 19612
rect 10157 19556 10161 19612
rect 10097 19552 10161 19556
rect 10177 19612 10241 19616
rect 10177 19556 10181 19612
rect 10181 19556 10237 19612
rect 10237 19556 10241 19612
rect 10177 19552 10241 19556
rect 13492 19544 13556 19548
rect 13492 19488 13506 19544
rect 13506 19488 13556 19544
rect 13492 19484 13556 19488
rect 8156 19408 8220 19412
rect 8156 19352 8170 19408
rect 8170 19352 8220 19408
rect 8156 19348 8220 19352
rect 18922 19612 18986 19616
rect 18922 19556 18926 19612
rect 18926 19556 18982 19612
rect 18982 19556 18986 19612
rect 18922 19552 18986 19556
rect 19002 19612 19066 19616
rect 19002 19556 19006 19612
rect 19006 19556 19062 19612
rect 19062 19556 19066 19612
rect 19002 19552 19066 19556
rect 19082 19612 19146 19616
rect 19082 19556 19086 19612
rect 19086 19556 19142 19612
rect 19142 19556 19146 19612
rect 19082 19552 19146 19556
rect 19162 19612 19226 19616
rect 19162 19556 19166 19612
rect 19166 19556 19222 19612
rect 19222 19556 19226 19612
rect 19162 19552 19226 19556
rect 22876 19408 22940 19412
rect 22876 19352 22890 19408
rect 22890 19352 22940 19408
rect 22876 19348 22940 19352
rect 3004 19212 3068 19276
rect 11100 19212 11164 19276
rect 16252 19212 16316 19276
rect 16620 19212 16684 19276
rect 8156 19076 8220 19140
rect 15516 19076 15580 19140
rect 16804 19076 16868 19140
rect 5444 19068 5508 19072
rect 5444 19012 5448 19068
rect 5448 19012 5504 19068
rect 5504 19012 5508 19068
rect 5444 19008 5508 19012
rect 5524 19068 5588 19072
rect 5524 19012 5528 19068
rect 5528 19012 5584 19068
rect 5584 19012 5588 19068
rect 5524 19008 5588 19012
rect 5604 19068 5668 19072
rect 5604 19012 5608 19068
rect 5608 19012 5664 19068
rect 5664 19012 5668 19068
rect 5604 19008 5668 19012
rect 5684 19068 5748 19072
rect 5684 19012 5688 19068
rect 5688 19012 5744 19068
rect 5744 19012 5748 19068
rect 5684 19008 5748 19012
rect 14430 19068 14494 19072
rect 14430 19012 14434 19068
rect 14434 19012 14490 19068
rect 14490 19012 14494 19068
rect 14430 19008 14494 19012
rect 14510 19068 14574 19072
rect 14510 19012 14514 19068
rect 14514 19012 14570 19068
rect 14570 19012 14574 19068
rect 14510 19008 14574 19012
rect 14590 19068 14654 19072
rect 14590 19012 14594 19068
rect 14594 19012 14650 19068
rect 14650 19012 14654 19068
rect 14590 19008 14654 19012
rect 14670 19068 14734 19072
rect 14670 19012 14674 19068
rect 14674 19012 14730 19068
rect 14730 19012 14734 19068
rect 14670 19008 14734 19012
rect 23415 19068 23479 19072
rect 23415 19012 23419 19068
rect 23419 19012 23475 19068
rect 23475 19012 23479 19068
rect 23415 19008 23479 19012
rect 23495 19068 23559 19072
rect 23495 19012 23499 19068
rect 23499 19012 23555 19068
rect 23555 19012 23559 19068
rect 23495 19008 23559 19012
rect 23575 19068 23639 19072
rect 23575 19012 23579 19068
rect 23579 19012 23635 19068
rect 23635 19012 23639 19068
rect 23575 19008 23639 19012
rect 23655 19068 23719 19072
rect 23655 19012 23659 19068
rect 23659 19012 23715 19068
rect 23715 19012 23719 19068
rect 23655 19008 23719 19012
rect 4660 18940 4724 19004
rect 5948 18940 6012 19004
rect 9628 18940 9692 19004
rect 12020 18940 12084 19004
rect 17908 18940 17972 19004
rect 2636 18804 2700 18868
rect 10732 18804 10796 18868
rect 18092 18804 18156 18868
rect 2820 18668 2884 18732
rect 3188 18668 3252 18732
rect 15516 18668 15580 18732
rect 16068 18668 16132 18732
rect 3924 18532 3988 18596
rect 5948 18532 6012 18596
rect 6316 18532 6380 18596
rect 9937 18524 10001 18528
rect 9937 18468 9941 18524
rect 9941 18468 9997 18524
rect 9997 18468 10001 18524
rect 9937 18464 10001 18468
rect 10017 18524 10081 18528
rect 10017 18468 10021 18524
rect 10021 18468 10077 18524
rect 10077 18468 10081 18524
rect 10017 18464 10081 18468
rect 10097 18524 10161 18528
rect 10097 18468 10101 18524
rect 10101 18468 10157 18524
rect 10157 18468 10161 18524
rect 10097 18464 10161 18468
rect 10177 18524 10241 18528
rect 10177 18468 10181 18524
rect 10181 18468 10237 18524
rect 10237 18468 10241 18524
rect 10177 18464 10241 18468
rect 4292 18260 4356 18324
rect 5212 18396 5276 18460
rect 7788 18396 7852 18460
rect 10916 18396 10980 18460
rect 18276 18456 18340 18460
rect 18922 18524 18986 18528
rect 18922 18468 18926 18524
rect 18926 18468 18982 18524
rect 18982 18468 18986 18524
rect 18922 18464 18986 18468
rect 19002 18524 19066 18528
rect 19002 18468 19006 18524
rect 19006 18468 19062 18524
rect 19062 18468 19066 18524
rect 19002 18464 19066 18468
rect 19082 18524 19146 18528
rect 19082 18468 19086 18524
rect 19086 18468 19142 18524
rect 19142 18468 19146 18524
rect 19082 18464 19146 18468
rect 19162 18524 19226 18528
rect 19162 18468 19166 18524
rect 19166 18468 19222 18524
rect 19222 18468 19226 18524
rect 19162 18464 19226 18468
rect 18276 18400 18290 18456
rect 18290 18400 18340 18456
rect 18276 18396 18340 18400
rect 6500 18260 6564 18324
rect 5028 18124 5092 18188
rect 5212 18124 5276 18188
rect 10364 18124 10428 18188
rect 13676 18124 13740 18188
rect 16988 18124 17052 18188
rect 11468 17988 11532 18052
rect 16804 17988 16868 18052
rect 5444 17980 5508 17984
rect 5444 17924 5448 17980
rect 5448 17924 5504 17980
rect 5504 17924 5508 17980
rect 5444 17920 5508 17924
rect 5524 17980 5588 17984
rect 5524 17924 5528 17980
rect 5528 17924 5584 17980
rect 5584 17924 5588 17980
rect 5524 17920 5588 17924
rect 5604 17980 5668 17984
rect 5604 17924 5608 17980
rect 5608 17924 5664 17980
rect 5664 17924 5668 17980
rect 5604 17920 5668 17924
rect 5684 17980 5748 17984
rect 5684 17924 5688 17980
rect 5688 17924 5744 17980
rect 5744 17924 5748 17980
rect 5684 17920 5748 17924
rect 14430 17980 14494 17984
rect 14430 17924 14434 17980
rect 14434 17924 14490 17980
rect 14490 17924 14494 17980
rect 14430 17920 14494 17924
rect 14510 17980 14574 17984
rect 14510 17924 14514 17980
rect 14514 17924 14570 17980
rect 14570 17924 14574 17980
rect 14510 17920 14574 17924
rect 14590 17980 14654 17984
rect 14590 17924 14594 17980
rect 14594 17924 14650 17980
rect 14650 17924 14654 17980
rect 14590 17920 14654 17924
rect 14670 17980 14734 17984
rect 14670 17924 14674 17980
rect 14674 17924 14730 17980
rect 14730 17924 14734 17980
rect 14670 17920 14734 17924
rect 23415 17980 23479 17984
rect 23415 17924 23419 17980
rect 23419 17924 23475 17980
rect 23475 17924 23479 17980
rect 23415 17920 23479 17924
rect 23495 17980 23559 17984
rect 23495 17924 23499 17980
rect 23499 17924 23555 17980
rect 23555 17924 23559 17980
rect 23495 17920 23559 17924
rect 23575 17980 23639 17984
rect 23575 17924 23579 17980
rect 23579 17924 23635 17980
rect 23635 17924 23639 17980
rect 23575 17920 23639 17924
rect 23655 17980 23719 17984
rect 23655 17924 23659 17980
rect 23659 17924 23715 17980
rect 23715 17924 23719 17980
rect 23655 17920 23719 17924
rect 10548 17852 10612 17916
rect 2820 17716 2884 17780
rect 13492 17716 13556 17780
rect 21036 17716 21100 17780
rect 4844 17580 4908 17644
rect 15148 17580 15212 17644
rect 11468 17444 11532 17508
rect 9937 17436 10001 17440
rect 9937 17380 9941 17436
rect 9941 17380 9997 17436
rect 9997 17380 10001 17436
rect 9937 17376 10001 17380
rect 10017 17436 10081 17440
rect 10017 17380 10021 17436
rect 10021 17380 10077 17436
rect 10077 17380 10081 17436
rect 10017 17376 10081 17380
rect 10097 17436 10161 17440
rect 10097 17380 10101 17436
rect 10101 17380 10157 17436
rect 10157 17380 10161 17436
rect 10097 17376 10161 17380
rect 10177 17436 10241 17440
rect 10177 17380 10181 17436
rect 10181 17380 10237 17436
rect 10237 17380 10241 17436
rect 10177 17376 10241 17380
rect 7052 17308 7116 17372
rect 17356 17444 17420 17508
rect 18922 17436 18986 17440
rect 18922 17380 18926 17436
rect 18926 17380 18982 17436
rect 18982 17380 18986 17436
rect 18922 17376 18986 17380
rect 19002 17436 19066 17440
rect 19002 17380 19006 17436
rect 19006 17380 19062 17436
rect 19062 17380 19066 17436
rect 19002 17376 19066 17380
rect 19082 17436 19146 17440
rect 19082 17380 19086 17436
rect 19086 17380 19142 17436
rect 19142 17380 19146 17436
rect 19082 17376 19146 17380
rect 19162 17436 19226 17440
rect 19162 17380 19166 17436
rect 19166 17380 19222 17436
rect 19222 17380 19226 17436
rect 19162 17376 19226 17380
rect 14044 17172 14108 17236
rect 7420 17096 7484 17100
rect 7420 17040 7434 17096
rect 7434 17040 7484 17096
rect 7420 17036 7484 17040
rect 11836 17036 11900 17100
rect 17172 17036 17236 17100
rect 18276 17096 18340 17100
rect 18276 17040 18290 17096
rect 18290 17040 18340 17096
rect 18276 17036 18340 17040
rect 16804 16900 16868 16964
rect 18460 16960 18524 16964
rect 18460 16904 18474 16960
rect 18474 16904 18524 16960
rect 18460 16900 18524 16904
rect 5444 16892 5508 16896
rect 5444 16836 5448 16892
rect 5448 16836 5504 16892
rect 5504 16836 5508 16892
rect 5444 16832 5508 16836
rect 5524 16892 5588 16896
rect 5524 16836 5528 16892
rect 5528 16836 5584 16892
rect 5584 16836 5588 16892
rect 5524 16832 5588 16836
rect 5604 16892 5668 16896
rect 5604 16836 5608 16892
rect 5608 16836 5664 16892
rect 5664 16836 5668 16892
rect 5604 16832 5668 16836
rect 5684 16892 5748 16896
rect 5684 16836 5688 16892
rect 5688 16836 5744 16892
rect 5744 16836 5748 16892
rect 5684 16832 5748 16836
rect 14430 16892 14494 16896
rect 14430 16836 14434 16892
rect 14434 16836 14490 16892
rect 14490 16836 14494 16892
rect 14430 16832 14494 16836
rect 14510 16892 14574 16896
rect 14510 16836 14514 16892
rect 14514 16836 14570 16892
rect 14570 16836 14574 16892
rect 14510 16832 14574 16836
rect 14590 16892 14654 16896
rect 14590 16836 14594 16892
rect 14594 16836 14650 16892
rect 14650 16836 14654 16892
rect 14590 16832 14654 16836
rect 14670 16892 14734 16896
rect 14670 16836 14674 16892
rect 14674 16836 14730 16892
rect 14730 16836 14734 16892
rect 14670 16832 14734 16836
rect 23415 16892 23479 16896
rect 23415 16836 23419 16892
rect 23419 16836 23475 16892
rect 23475 16836 23479 16892
rect 23415 16832 23479 16836
rect 23495 16892 23559 16896
rect 23495 16836 23499 16892
rect 23499 16836 23555 16892
rect 23555 16836 23559 16892
rect 23495 16832 23559 16836
rect 23575 16892 23639 16896
rect 23575 16836 23579 16892
rect 23579 16836 23635 16892
rect 23635 16836 23639 16892
rect 23575 16832 23639 16836
rect 23655 16892 23719 16896
rect 23655 16836 23659 16892
rect 23659 16836 23715 16892
rect 23715 16836 23719 16892
rect 23655 16832 23719 16836
rect 16252 16764 16316 16828
rect 18276 16764 18340 16828
rect 15516 16628 15580 16692
rect 22692 16628 22756 16692
rect 16620 16356 16684 16420
rect 22876 16356 22940 16420
rect 9937 16348 10001 16352
rect 9937 16292 9941 16348
rect 9941 16292 9997 16348
rect 9997 16292 10001 16348
rect 9937 16288 10001 16292
rect 10017 16348 10081 16352
rect 10017 16292 10021 16348
rect 10021 16292 10077 16348
rect 10077 16292 10081 16348
rect 10017 16288 10081 16292
rect 10097 16348 10161 16352
rect 10097 16292 10101 16348
rect 10101 16292 10157 16348
rect 10157 16292 10161 16348
rect 10097 16288 10161 16292
rect 10177 16348 10241 16352
rect 10177 16292 10181 16348
rect 10181 16292 10237 16348
rect 10237 16292 10241 16348
rect 10177 16288 10241 16292
rect 18922 16348 18986 16352
rect 18922 16292 18926 16348
rect 18926 16292 18982 16348
rect 18982 16292 18986 16348
rect 18922 16288 18986 16292
rect 19002 16348 19066 16352
rect 19002 16292 19006 16348
rect 19006 16292 19062 16348
rect 19062 16292 19066 16348
rect 19002 16288 19066 16292
rect 19082 16348 19146 16352
rect 19082 16292 19086 16348
rect 19086 16292 19142 16348
rect 19142 16292 19146 16348
rect 19082 16288 19146 16292
rect 19162 16348 19226 16352
rect 19162 16292 19166 16348
rect 19166 16292 19222 16348
rect 19222 16292 19226 16348
rect 19162 16288 19226 16292
rect 2820 16280 2884 16284
rect 2820 16224 2834 16280
rect 2834 16224 2884 16280
rect 2820 16220 2884 16224
rect 18644 16220 18708 16284
rect 16252 16084 16316 16148
rect 16620 15948 16684 16012
rect 5444 15804 5508 15808
rect 5444 15748 5448 15804
rect 5448 15748 5504 15804
rect 5504 15748 5508 15804
rect 5444 15744 5508 15748
rect 5524 15804 5588 15808
rect 5524 15748 5528 15804
rect 5528 15748 5584 15804
rect 5584 15748 5588 15804
rect 5524 15744 5588 15748
rect 5604 15804 5668 15808
rect 5604 15748 5608 15804
rect 5608 15748 5664 15804
rect 5664 15748 5668 15804
rect 5604 15744 5668 15748
rect 5684 15804 5748 15808
rect 5684 15748 5688 15804
rect 5688 15748 5744 15804
rect 5744 15748 5748 15804
rect 5684 15744 5748 15748
rect 14430 15804 14494 15808
rect 14430 15748 14434 15804
rect 14434 15748 14490 15804
rect 14490 15748 14494 15804
rect 14430 15744 14494 15748
rect 14510 15804 14574 15808
rect 14510 15748 14514 15804
rect 14514 15748 14570 15804
rect 14570 15748 14574 15804
rect 14510 15744 14574 15748
rect 14590 15804 14654 15808
rect 14590 15748 14594 15804
rect 14594 15748 14650 15804
rect 14650 15748 14654 15804
rect 14590 15744 14654 15748
rect 14670 15804 14734 15808
rect 14670 15748 14674 15804
rect 14674 15748 14730 15804
rect 14730 15748 14734 15804
rect 14670 15744 14734 15748
rect 23415 15804 23479 15808
rect 23415 15748 23419 15804
rect 23419 15748 23475 15804
rect 23475 15748 23479 15804
rect 23415 15744 23479 15748
rect 23495 15804 23559 15808
rect 23495 15748 23499 15804
rect 23499 15748 23555 15804
rect 23555 15748 23559 15804
rect 23495 15744 23559 15748
rect 23575 15804 23639 15808
rect 23575 15748 23579 15804
rect 23579 15748 23635 15804
rect 23635 15748 23639 15804
rect 23575 15744 23639 15748
rect 23655 15804 23719 15808
rect 23655 15748 23659 15804
rect 23659 15748 23715 15804
rect 23715 15748 23719 15804
rect 23655 15744 23719 15748
rect 3740 15676 3804 15740
rect 6684 15540 6748 15604
rect 23244 15464 23308 15468
rect 23244 15408 23258 15464
rect 23258 15408 23308 15464
rect 6316 15268 6380 15332
rect 9937 15260 10001 15264
rect 9937 15204 9941 15260
rect 9941 15204 9997 15260
rect 9997 15204 10001 15260
rect 9937 15200 10001 15204
rect 10017 15260 10081 15264
rect 10017 15204 10021 15260
rect 10021 15204 10077 15260
rect 10077 15204 10081 15260
rect 10017 15200 10081 15204
rect 10097 15260 10161 15264
rect 10097 15204 10101 15260
rect 10101 15204 10157 15260
rect 10157 15204 10161 15260
rect 10097 15200 10161 15204
rect 10177 15260 10241 15264
rect 10177 15204 10181 15260
rect 10181 15204 10237 15260
rect 10237 15204 10241 15260
rect 10177 15200 10241 15204
rect 23244 15404 23308 15408
rect 21772 15268 21836 15332
rect 18922 15260 18986 15264
rect 18922 15204 18926 15260
rect 18926 15204 18982 15260
rect 18982 15204 18986 15260
rect 18922 15200 18986 15204
rect 19002 15260 19066 15264
rect 19002 15204 19006 15260
rect 19006 15204 19062 15260
rect 19062 15204 19066 15260
rect 19002 15200 19066 15204
rect 19082 15260 19146 15264
rect 19082 15204 19086 15260
rect 19086 15204 19142 15260
rect 19142 15204 19146 15260
rect 19082 15200 19146 15204
rect 19162 15260 19226 15264
rect 19162 15204 19166 15260
rect 19166 15204 19222 15260
rect 19222 15204 19226 15260
rect 19162 15200 19226 15204
rect 11652 14860 11716 14924
rect 9076 14724 9140 14788
rect 24532 14996 24596 15060
rect 17356 14860 17420 14924
rect 5444 14716 5508 14720
rect 5444 14660 5448 14716
rect 5448 14660 5504 14716
rect 5504 14660 5508 14716
rect 5444 14656 5508 14660
rect 5524 14716 5588 14720
rect 5524 14660 5528 14716
rect 5528 14660 5584 14716
rect 5584 14660 5588 14716
rect 5524 14656 5588 14660
rect 5604 14716 5668 14720
rect 5604 14660 5608 14716
rect 5608 14660 5664 14716
rect 5664 14660 5668 14716
rect 5604 14656 5668 14660
rect 5684 14716 5748 14720
rect 5684 14660 5688 14716
rect 5688 14660 5744 14716
rect 5744 14660 5748 14716
rect 5684 14656 5748 14660
rect 14430 14716 14494 14720
rect 14430 14660 14434 14716
rect 14434 14660 14490 14716
rect 14490 14660 14494 14716
rect 14430 14656 14494 14660
rect 14510 14716 14574 14720
rect 14510 14660 14514 14716
rect 14514 14660 14570 14716
rect 14570 14660 14574 14716
rect 14510 14656 14574 14660
rect 14590 14716 14654 14720
rect 14590 14660 14594 14716
rect 14594 14660 14650 14716
rect 14650 14660 14654 14716
rect 14590 14656 14654 14660
rect 14670 14716 14734 14720
rect 14670 14660 14674 14716
rect 14674 14660 14730 14716
rect 14730 14660 14734 14716
rect 14670 14656 14734 14660
rect 23415 14716 23479 14720
rect 23415 14660 23419 14716
rect 23419 14660 23475 14716
rect 23475 14660 23479 14716
rect 23415 14656 23479 14660
rect 23495 14716 23559 14720
rect 23495 14660 23499 14716
rect 23499 14660 23555 14716
rect 23555 14660 23559 14716
rect 23495 14656 23559 14660
rect 23575 14716 23639 14720
rect 23575 14660 23579 14716
rect 23579 14660 23635 14716
rect 23635 14660 23639 14716
rect 23575 14656 23639 14660
rect 23655 14716 23719 14720
rect 23655 14660 23659 14716
rect 23659 14660 23715 14716
rect 23715 14660 23719 14716
rect 23655 14656 23719 14660
rect 15884 14588 15948 14652
rect 24164 14452 24228 14516
rect 3924 14376 3988 14380
rect 3924 14320 3938 14376
rect 3938 14320 3988 14376
rect 3924 14316 3988 14320
rect 13492 14316 13556 14380
rect 18644 14316 18708 14380
rect 20668 14316 20732 14380
rect 11284 14180 11348 14244
rect 16252 14180 16316 14244
rect 9937 14172 10001 14176
rect 9937 14116 9941 14172
rect 9941 14116 9997 14172
rect 9997 14116 10001 14172
rect 9937 14112 10001 14116
rect 10017 14172 10081 14176
rect 10017 14116 10021 14172
rect 10021 14116 10077 14172
rect 10077 14116 10081 14172
rect 10017 14112 10081 14116
rect 10097 14172 10161 14176
rect 10097 14116 10101 14172
rect 10101 14116 10157 14172
rect 10157 14116 10161 14172
rect 10097 14112 10161 14116
rect 10177 14172 10241 14176
rect 10177 14116 10181 14172
rect 10181 14116 10237 14172
rect 10237 14116 10241 14172
rect 10177 14112 10241 14116
rect 18922 14172 18986 14176
rect 18922 14116 18926 14172
rect 18926 14116 18982 14172
rect 18982 14116 18986 14172
rect 18922 14112 18986 14116
rect 19002 14172 19066 14176
rect 19002 14116 19006 14172
rect 19006 14116 19062 14172
rect 19062 14116 19066 14172
rect 19002 14112 19066 14116
rect 19082 14172 19146 14176
rect 19082 14116 19086 14172
rect 19086 14116 19142 14172
rect 19142 14116 19146 14172
rect 19082 14112 19146 14116
rect 19162 14172 19226 14176
rect 19162 14116 19166 14172
rect 19166 14116 19222 14172
rect 19222 14116 19226 14172
rect 19162 14112 19226 14116
rect 3556 13908 3620 13972
rect 11652 13908 11716 13972
rect 15516 13968 15580 13972
rect 15516 13912 15530 13968
rect 15530 13912 15580 13968
rect 15516 13908 15580 13912
rect 16068 13772 16132 13836
rect 17724 13772 17788 13836
rect 4108 13636 4172 13700
rect 17540 13696 17604 13700
rect 17540 13640 17590 13696
rect 17590 13640 17604 13696
rect 17540 13636 17604 13640
rect 5444 13628 5508 13632
rect 5444 13572 5448 13628
rect 5448 13572 5504 13628
rect 5504 13572 5508 13628
rect 5444 13568 5508 13572
rect 5524 13628 5588 13632
rect 5524 13572 5528 13628
rect 5528 13572 5584 13628
rect 5584 13572 5588 13628
rect 5524 13568 5588 13572
rect 5604 13628 5668 13632
rect 5604 13572 5608 13628
rect 5608 13572 5664 13628
rect 5664 13572 5668 13628
rect 5604 13568 5668 13572
rect 5684 13628 5748 13632
rect 5684 13572 5688 13628
rect 5688 13572 5744 13628
rect 5744 13572 5748 13628
rect 5684 13568 5748 13572
rect 14430 13628 14494 13632
rect 14430 13572 14434 13628
rect 14434 13572 14490 13628
rect 14490 13572 14494 13628
rect 14430 13568 14494 13572
rect 14510 13628 14574 13632
rect 14510 13572 14514 13628
rect 14514 13572 14570 13628
rect 14570 13572 14574 13628
rect 14510 13568 14574 13572
rect 14590 13628 14654 13632
rect 14590 13572 14594 13628
rect 14594 13572 14650 13628
rect 14650 13572 14654 13628
rect 14590 13568 14654 13572
rect 14670 13628 14734 13632
rect 14670 13572 14674 13628
rect 14674 13572 14730 13628
rect 14730 13572 14734 13628
rect 14670 13568 14734 13572
rect 23415 13628 23479 13632
rect 23415 13572 23419 13628
rect 23419 13572 23475 13628
rect 23475 13572 23479 13628
rect 23415 13568 23479 13572
rect 23495 13628 23559 13632
rect 23495 13572 23499 13628
rect 23499 13572 23555 13628
rect 23555 13572 23559 13628
rect 23495 13568 23559 13572
rect 23575 13628 23639 13632
rect 23575 13572 23579 13628
rect 23579 13572 23635 13628
rect 23635 13572 23639 13628
rect 23575 13568 23639 13572
rect 23655 13628 23719 13632
rect 23655 13572 23659 13628
rect 23659 13572 23715 13628
rect 23715 13572 23719 13628
rect 23655 13568 23719 13572
rect 3188 13560 3252 13564
rect 3188 13504 3238 13560
rect 3238 13504 3252 13560
rect 3188 13500 3252 13504
rect 17908 13364 17972 13428
rect 5212 13288 5276 13292
rect 5212 13232 5226 13288
rect 5226 13232 5276 13288
rect 3556 13016 3620 13020
rect 3556 12960 3606 13016
rect 3606 12960 3620 13016
rect 3556 12956 3620 12960
rect 3188 12820 3252 12884
rect 5212 13228 5276 13232
rect 8708 13228 8772 13292
rect 9444 13092 9508 13156
rect 18460 13152 18524 13156
rect 18460 13096 18510 13152
rect 18510 13096 18524 13152
rect 18460 13092 18524 13096
rect 23244 13092 23308 13156
rect 9937 13084 10001 13088
rect 9937 13028 9941 13084
rect 9941 13028 9997 13084
rect 9997 13028 10001 13084
rect 9937 13024 10001 13028
rect 10017 13084 10081 13088
rect 10017 13028 10021 13084
rect 10021 13028 10077 13084
rect 10077 13028 10081 13084
rect 10017 13024 10081 13028
rect 10097 13084 10161 13088
rect 10097 13028 10101 13084
rect 10101 13028 10157 13084
rect 10157 13028 10161 13084
rect 10097 13024 10161 13028
rect 10177 13084 10241 13088
rect 10177 13028 10181 13084
rect 10181 13028 10237 13084
rect 10237 13028 10241 13084
rect 10177 13024 10241 13028
rect 18922 13084 18986 13088
rect 18922 13028 18926 13084
rect 18926 13028 18982 13084
rect 18982 13028 18986 13084
rect 18922 13024 18986 13028
rect 19002 13084 19066 13088
rect 19002 13028 19006 13084
rect 19006 13028 19062 13084
rect 19062 13028 19066 13084
rect 19002 13024 19066 13028
rect 19082 13084 19146 13088
rect 19082 13028 19086 13084
rect 19086 13028 19142 13084
rect 19142 13028 19146 13084
rect 19082 13024 19146 13028
rect 19162 13084 19226 13088
rect 19162 13028 19166 13084
rect 19166 13028 19222 13084
rect 19222 13028 19226 13084
rect 19162 13024 19226 13028
rect 4660 12956 4724 13020
rect 15148 12956 15212 13020
rect 4660 12820 4724 12884
rect 8524 12880 8588 12884
rect 8524 12824 8574 12880
rect 8574 12824 8588 12880
rect 8524 12820 8588 12824
rect 14964 12820 15028 12884
rect 4476 12684 4540 12748
rect 7788 12744 7852 12748
rect 7788 12688 7838 12744
rect 7838 12688 7852 12744
rect 4476 12548 4540 12612
rect 3004 12412 3068 12476
rect 4844 12412 4908 12476
rect 7788 12684 7852 12688
rect 7972 12684 8036 12748
rect 5212 12608 5276 12612
rect 5212 12552 5262 12608
rect 5262 12552 5276 12608
rect 5212 12548 5276 12552
rect 6500 12608 6564 12612
rect 6500 12552 6550 12608
rect 6550 12552 6564 12608
rect 6500 12548 6564 12552
rect 5444 12540 5508 12544
rect 5444 12484 5448 12540
rect 5448 12484 5504 12540
rect 5504 12484 5508 12540
rect 5444 12480 5508 12484
rect 5524 12540 5588 12544
rect 5524 12484 5528 12540
rect 5528 12484 5584 12540
rect 5584 12484 5588 12540
rect 5524 12480 5588 12484
rect 5604 12540 5668 12544
rect 5604 12484 5608 12540
rect 5608 12484 5664 12540
rect 5664 12484 5668 12540
rect 5604 12480 5668 12484
rect 5684 12540 5748 12544
rect 5684 12484 5688 12540
rect 5688 12484 5744 12540
rect 5744 12484 5748 12540
rect 5684 12480 5748 12484
rect 8708 12548 8772 12612
rect 7052 12472 7116 12476
rect 7052 12416 7066 12472
rect 7066 12416 7116 12472
rect 7052 12412 7116 12416
rect 7236 12412 7300 12476
rect 14430 12540 14494 12544
rect 14430 12484 14434 12540
rect 14434 12484 14490 12540
rect 14490 12484 14494 12540
rect 14430 12480 14494 12484
rect 14510 12540 14574 12544
rect 14510 12484 14514 12540
rect 14514 12484 14570 12540
rect 14570 12484 14574 12540
rect 14510 12480 14574 12484
rect 14590 12540 14654 12544
rect 14590 12484 14594 12540
rect 14594 12484 14650 12540
rect 14650 12484 14654 12540
rect 14590 12480 14654 12484
rect 14670 12540 14734 12544
rect 14670 12484 14674 12540
rect 14674 12484 14730 12540
rect 14730 12484 14734 12540
rect 14670 12480 14734 12484
rect 9260 12412 9324 12476
rect 22876 12684 22940 12748
rect 21404 12548 21468 12612
rect 23415 12540 23479 12544
rect 23415 12484 23419 12540
rect 23419 12484 23475 12540
rect 23475 12484 23479 12540
rect 23415 12480 23479 12484
rect 23495 12540 23559 12544
rect 23495 12484 23499 12540
rect 23499 12484 23555 12540
rect 23555 12484 23559 12540
rect 23495 12480 23559 12484
rect 23575 12540 23639 12544
rect 23575 12484 23579 12540
rect 23579 12484 23635 12540
rect 23635 12484 23639 12540
rect 23575 12480 23639 12484
rect 23655 12540 23719 12544
rect 23655 12484 23659 12540
rect 23659 12484 23715 12540
rect 23715 12484 23719 12540
rect 23655 12480 23719 12484
rect 24164 12472 24228 12476
rect 24164 12416 24178 12472
rect 24178 12416 24228 12472
rect 24164 12412 24228 12416
rect 4476 12336 4540 12340
rect 4476 12280 4526 12336
rect 4526 12280 4540 12336
rect 4476 12276 4540 12280
rect 6500 12336 6564 12340
rect 6500 12280 6550 12336
rect 6550 12280 6564 12336
rect 6500 12276 6564 12280
rect 6868 12276 6932 12340
rect 7052 12276 7116 12340
rect 7420 12336 7484 12340
rect 7420 12280 7434 12336
rect 7434 12280 7484 12336
rect 7420 12276 7484 12280
rect 7788 12336 7852 12340
rect 7788 12280 7802 12336
rect 7802 12280 7852 12336
rect 7788 12276 7852 12280
rect 8524 12276 8588 12340
rect 10916 12336 10980 12340
rect 10916 12280 10930 12336
rect 10930 12280 10980 12336
rect 10916 12276 10980 12280
rect 16436 12276 16500 12340
rect 10732 12200 10796 12204
rect 10732 12144 10782 12200
rect 10782 12144 10796 12200
rect 10732 12140 10796 12144
rect 17356 12140 17420 12204
rect 17908 12140 17972 12204
rect 3004 12064 3068 12068
rect 3004 12008 3018 12064
rect 3018 12008 3068 12064
rect 3004 12004 3068 12008
rect 4292 12004 4356 12068
rect 4660 12064 4724 12068
rect 4660 12008 4710 12064
rect 4710 12008 4724 12064
rect 4660 12004 4724 12008
rect 6684 12004 6748 12068
rect 7604 12004 7668 12068
rect 14044 12004 14108 12068
rect 17356 12004 17420 12068
rect 9937 11996 10001 12000
rect 9937 11940 9941 11996
rect 9941 11940 9997 11996
rect 9997 11940 10001 11996
rect 9937 11936 10001 11940
rect 10017 11996 10081 12000
rect 10017 11940 10021 11996
rect 10021 11940 10077 11996
rect 10077 11940 10081 11996
rect 10017 11936 10081 11940
rect 10097 11996 10161 12000
rect 10097 11940 10101 11996
rect 10101 11940 10157 11996
rect 10157 11940 10161 11996
rect 10097 11936 10161 11940
rect 10177 11996 10241 12000
rect 10177 11940 10181 11996
rect 10181 11940 10237 11996
rect 10237 11940 10241 11996
rect 10177 11936 10241 11940
rect 5948 11868 6012 11932
rect 16988 11868 17052 11932
rect 18276 11868 18340 11932
rect 9444 11732 9508 11796
rect 12020 11732 12084 11796
rect 17540 11732 17604 11796
rect 21404 12004 21468 12068
rect 18922 11996 18986 12000
rect 18922 11940 18926 11996
rect 18926 11940 18982 11996
rect 18982 11940 18986 11996
rect 18922 11936 18986 11940
rect 19002 11996 19066 12000
rect 19002 11940 19006 11996
rect 19006 11940 19062 11996
rect 19062 11940 19066 11996
rect 19002 11936 19066 11940
rect 19082 11996 19146 12000
rect 19082 11940 19086 11996
rect 19086 11940 19142 11996
rect 19142 11940 19146 11996
rect 19082 11936 19146 11940
rect 19162 11996 19226 12000
rect 19162 11940 19166 11996
rect 19166 11940 19222 11996
rect 19222 11940 19226 11996
rect 19162 11936 19226 11940
rect 21220 11928 21284 11932
rect 21220 11872 21234 11928
rect 21234 11872 21284 11928
rect 21220 11868 21284 11872
rect 3924 11596 3988 11660
rect 17724 11596 17788 11660
rect 21772 11596 21836 11660
rect 24532 11596 24596 11660
rect 15332 11460 15396 11524
rect 18460 11460 18524 11524
rect 5444 11452 5508 11456
rect 5444 11396 5448 11452
rect 5448 11396 5504 11452
rect 5504 11396 5508 11452
rect 5444 11392 5508 11396
rect 5524 11452 5588 11456
rect 5524 11396 5528 11452
rect 5528 11396 5584 11452
rect 5584 11396 5588 11452
rect 5524 11392 5588 11396
rect 5604 11452 5668 11456
rect 5604 11396 5608 11452
rect 5608 11396 5664 11452
rect 5664 11396 5668 11452
rect 5604 11392 5668 11396
rect 5684 11452 5748 11456
rect 5684 11396 5688 11452
rect 5688 11396 5744 11452
rect 5744 11396 5748 11452
rect 5684 11392 5748 11396
rect 14430 11452 14494 11456
rect 14430 11396 14434 11452
rect 14434 11396 14490 11452
rect 14490 11396 14494 11452
rect 14430 11392 14494 11396
rect 14510 11452 14574 11456
rect 14510 11396 14514 11452
rect 14514 11396 14570 11452
rect 14570 11396 14574 11452
rect 14510 11392 14574 11396
rect 14590 11452 14654 11456
rect 14590 11396 14594 11452
rect 14594 11396 14650 11452
rect 14650 11396 14654 11452
rect 14590 11392 14654 11396
rect 14670 11452 14734 11456
rect 14670 11396 14674 11452
rect 14674 11396 14730 11452
rect 14730 11396 14734 11452
rect 14670 11392 14734 11396
rect 23415 11452 23479 11456
rect 23415 11396 23419 11452
rect 23419 11396 23475 11452
rect 23475 11396 23479 11452
rect 23415 11392 23479 11396
rect 23495 11452 23559 11456
rect 23495 11396 23499 11452
rect 23499 11396 23555 11452
rect 23555 11396 23559 11452
rect 23495 11392 23559 11396
rect 23575 11452 23639 11456
rect 23575 11396 23579 11452
rect 23579 11396 23635 11452
rect 23635 11396 23639 11452
rect 23575 11392 23639 11396
rect 23655 11452 23719 11456
rect 23655 11396 23659 11452
rect 23659 11396 23715 11452
rect 23715 11396 23719 11452
rect 23655 11392 23719 11396
rect 9076 11188 9140 11252
rect 7604 11112 7668 11116
rect 7604 11056 7654 11112
rect 7654 11056 7668 11112
rect 7604 11052 7668 11056
rect 15884 11052 15948 11116
rect 18092 11112 18156 11116
rect 18092 11056 18106 11112
rect 18106 11056 18156 11112
rect 18092 11052 18156 11056
rect 21956 11052 22020 11116
rect 6316 10916 6380 10980
rect 11836 10916 11900 10980
rect 9937 10908 10001 10912
rect 9937 10852 9941 10908
rect 9941 10852 9997 10908
rect 9997 10852 10001 10908
rect 9937 10848 10001 10852
rect 10017 10908 10081 10912
rect 10017 10852 10021 10908
rect 10021 10852 10077 10908
rect 10077 10852 10081 10908
rect 10017 10848 10081 10852
rect 10097 10908 10161 10912
rect 10097 10852 10101 10908
rect 10101 10852 10157 10908
rect 10157 10852 10161 10908
rect 10097 10848 10161 10852
rect 10177 10908 10241 10912
rect 10177 10852 10181 10908
rect 10181 10852 10237 10908
rect 10237 10852 10241 10908
rect 10177 10848 10241 10852
rect 18922 10908 18986 10912
rect 18922 10852 18926 10908
rect 18926 10852 18982 10908
rect 18982 10852 18986 10908
rect 18922 10848 18986 10852
rect 19002 10908 19066 10912
rect 19002 10852 19006 10908
rect 19006 10852 19062 10908
rect 19062 10852 19066 10908
rect 19002 10848 19066 10852
rect 19082 10908 19146 10912
rect 19082 10852 19086 10908
rect 19086 10852 19142 10908
rect 19142 10852 19146 10908
rect 19082 10848 19146 10852
rect 19162 10908 19226 10912
rect 19162 10852 19166 10908
rect 19166 10852 19222 10908
rect 19222 10852 19226 10908
rect 19162 10848 19226 10852
rect 8156 10780 8220 10844
rect 20668 10840 20732 10844
rect 20668 10784 20718 10840
rect 20718 10784 20732 10840
rect 20668 10780 20732 10784
rect 10364 10508 10428 10572
rect 17172 10508 17236 10572
rect 22140 10508 22204 10572
rect 5444 10364 5508 10368
rect 5444 10308 5448 10364
rect 5448 10308 5504 10364
rect 5504 10308 5508 10364
rect 5444 10304 5508 10308
rect 5524 10364 5588 10368
rect 5524 10308 5528 10364
rect 5528 10308 5584 10364
rect 5584 10308 5588 10364
rect 5524 10304 5588 10308
rect 5604 10364 5668 10368
rect 5604 10308 5608 10364
rect 5608 10308 5664 10364
rect 5664 10308 5668 10364
rect 5604 10304 5668 10308
rect 5684 10364 5748 10368
rect 5684 10308 5688 10364
rect 5688 10308 5744 10364
rect 5744 10308 5748 10364
rect 5684 10304 5748 10308
rect 14430 10364 14494 10368
rect 14430 10308 14434 10364
rect 14434 10308 14490 10364
rect 14490 10308 14494 10364
rect 14430 10304 14494 10308
rect 14510 10364 14574 10368
rect 14510 10308 14514 10364
rect 14514 10308 14570 10364
rect 14570 10308 14574 10364
rect 14510 10304 14574 10308
rect 14590 10364 14654 10368
rect 14590 10308 14594 10364
rect 14594 10308 14650 10364
rect 14650 10308 14654 10364
rect 14590 10304 14654 10308
rect 14670 10364 14734 10368
rect 14670 10308 14674 10364
rect 14674 10308 14730 10364
rect 14730 10308 14734 10364
rect 14670 10304 14734 10308
rect 23415 10364 23479 10368
rect 23415 10308 23419 10364
rect 23419 10308 23475 10364
rect 23475 10308 23479 10364
rect 23415 10304 23479 10308
rect 23495 10364 23559 10368
rect 23495 10308 23499 10364
rect 23499 10308 23555 10364
rect 23555 10308 23559 10364
rect 23495 10304 23559 10308
rect 23575 10364 23639 10368
rect 23575 10308 23579 10364
rect 23579 10308 23635 10364
rect 23635 10308 23639 10364
rect 23575 10304 23639 10308
rect 23655 10364 23719 10368
rect 23655 10308 23659 10364
rect 23659 10308 23715 10364
rect 23715 10308 23719 10364
rect 23655 10304 23719 10308
rect 3740 10100 3804 10164
rect 9260 10100 9324 10164
rect 2820 9964 2884 10028
rect 6132 9964 6196 10028
rect 7052 9964 7116 10028
rect 5212 9828 5276 9892
rect 7972 9828 8036 9892
rect 10364 9888 10428 9892
rect 10364 9832 10378 9888
rect 10378 9832 10428 9888
rect 10364 9828 10428 9832
rect 14044 9828 14108 9892
rect 9937 9820 10001 9824
rect 9937 9764 9941 9820
rect 9941 9764 9997 9820
rect 9997 9764 10001 9820
rect 9937 9760 10001 9764
rect 10017 9820 10081 9824
rect 10017 9764 10021 9820
rect 10021 9764 10077 9820
rect 10077 9764 10081 9820
rect 10017 9760 10081 9764
rect 10097 9820 10161 9824
rect 10097 9764 10101 9820
rect 10101 9764 10157 9820
rect 10157 9764 10161 9820
rect 10097 9760 10161 9764
rect 10177 9820 10241 9824
rect 10177 9764 10181 9820
rect 10181 9764 10237 9820
rect 10237 9764 10241 9820
rect 10177 9760 10241 9764
rect 18922 9820 18986 9824
rect 18922 9764 18926 9820
rect 18926 9764 18982 9820
rect 18982 9764 18986 9820
rect 18922 9760 18986 9764
rect 19002 9820 19066 9824
rect 19002 9764 19006 9820
rect 19006 9764 19062 9820
rect 19062 9764 19066 9820
rect 19002 9760 19066 9764
rect 19082 9820 19146 9824
rect 19082 9764 19086 9820
rect 19086 9764 19142 9820
rect 19142 9764 19146 9820
rect 19082 9760 19146 9764
rect 19162 9820 19226 9824
rect 19162 9764 19166 9820
rect 19166 9764 19222 9820
rect 19222 9764 19226 9820
rect 19162 9760 19226 9764
rect 5028 9752 5092 9756
rect 5028 9696 5078 9752
rect 5078 9696 5092 9752
rect 5028 9692 5092 9696
rect 11100 9692 11164 9756
rect 18644 9556 18708 9620
rect 23980 9556 24044 9620
rect 21956 9420 22020 9484
rect 5444 9276 5508 9280
rect 5444 9220 5448 9276
rect 5448 9220 5504 9276
rect 5504 9220 5508 9276
rect 5444 9216 5508 9220
rect 5524 9276 5588 9280
rect 5524 9220 5528 9276
rect 5528 9220 5584 9276
rect 5584 9220 5588 9276
rect 5524 9216 5588 9220
rect 5604 9276 5668 9280
rect 5604 9220 5608 9276
rect 5608 9220 5664 9276
rect 5664 9220 5668 9276
rect 5604 9216 5668 9220
rect 5684 9276 5748 9280
rect 5684 9220 5688 9276
rect 5688 9220 5744 9276
rect 5744 9220 5748 9276
rect 5684 9216 5748 9220
rect 14430 9276 14494 9280
rect 14430 9220 14434 9276
rect 14434 9220 14490 9276
rect 14490 9220 14494 9276
rect 14430 9216 14494 9220
rect 14510 9276 14574 9280
rect 14510 9220 14514 9276
rect 14514 9220 14570 9276
rect 14570 9220 14574 9276
rect 14510 9216 14574 9220
rect 14590 9276 14654 9280
rect 14590 9220 14594 9276
rect 14594 9220 14650 9276
rect 14650 9220 14654 9276
rect 14590 9216 14654 9220
rect 14670 9276 14734 9280
rect 14670 9220 14674 9276
rect 14674 9220 14730 9276
rect 14730 9220 14734 9276
rect 14670 9216 14734 9220
rect 23415 9276 23479 9280
rect 23415 9220 23419 9276
rect 23419 9220 23475 9276
rect 23475 9220 23479 9276
rect 23415 9216 23479 9220
rect 23495 9276 23559 9280
rect 23495 9220 23499 9276
rect 23499 9220 23555 9276
rect 23555 9220 23559 9276
rect 23495 9216 23559 9220
rect 23575 9276 23639 9280
rect 23575 9220 23579 9276
rect 23579 9220 23635 9276
rect 23635 9220 23639 9276
rect 23575 9216 23639 9220
rect 23655 9276 23719 9280
rect 23655 9220 23659 9276
rect 23659 9220 23715 9276
rect 23715 9220 23719 9276
rect 23655 9216 23719 9220
rect 15700 9012 15764 9076
rect 16804 8876 16868 8940
rect 18460 8876 18524 8940
rect 9937 8732 10001 8736
rect 9937 8676 9941 8732
rect 9941 8676 9997 8732
rect 9997 8676 10001 8732
rect 9937 8672 10001 8676
rect 10017 8732 10081 8736
rect 10017 8676 10021 8732
rect 10021 8676 10077 8732
rect 10077 8676 10081 8732
rect 10017 8672 10081 8676
rect 10097 8732 10161 8736
rect 10097 8676 10101 8732
rect 10101 8676 10157 8732
rect 10157 8676 10161 8732
rect 10097 8672 10161 8676
rect 10177 8732 10241 8736
rect 10177 8676 10181 8732
rect 10181 8676 10237 8732
rect 10237 8676 10241 8732
rect 10177 8672 10241 8676
rect 18922 8732 18986 8736
rect 18922 8676 18926 8732
rect 18926 8676 18982 8732
rect 18982 8676 18986 8732
rect 18922 8672 18986 8676
rect 19002 8732 19066 8736
rect 19002 8676 19006 8732
rect 19006 8676 19062 8732
rect 19062 8676 19066 8732
rect 19002 8672 19066 8676
rect 19082 8732 19146 8736
rect 19082 8676 19086 8732
rect 19086 8676 19142 8732
rect 19142 8676 19146 8732
rect 19082 8672 19146 8676
rect 19162 8732 19226 8736
rect 19162 8676 19166 8732
rect 19166 8676 19222 8732
rect 19222 8676 19226 8732
rect 19162 8672 19226 8676
rect 2820 8468 2884 8532
rect 3740 8468 3804 8532
rect 9260 8468 9324 8532
rect 10364 8332 10428 8396
rect 11468 8332 11532 8396
rect 5444 8188 5508 8192
rect 5444 8132 5448 8188
rect 5448 8132 5504 8188
rect 5504 8132 5508 8188
rect 5444 8128 5508 8132
rect 5524 8188 5588 8192
rect 5524 8132 5528 8188
rect 5528 8132 5584 8188
rect 5584 8132 5588 8188
rect 5524 8128 5588 8132
rect 5604 8188 5668 8192
rect 5604 8132 5608 8188
rect 5608 8132 5664 8188
rect 5664 8132 5668 8188
rect 5604 8128 5668 8132
rect 5684 8188 5748 8192
rect 5684 8132 5688 8188
rect 5688 8132 5744 8188
rect 5744 8132 5748 8188
rect 5684 8128 5748 8132
rect 19564 8196 19628 8260
rect 20668 8196 20732 8260
rect 22324 8196 22388 8260
rect 14430 8188 14494 8192
rect 14430 8132 14434 8188
rect 14434 8132 14490 8188
rect 14490 8132 14494 8188
rect 14430 8128 14494 8132
rect 14510 8188 14574 8192
rect 14510 8132 14514 8188
rect 14514 8132 14570 8188
rect 14570 8132 14574 8188
rect 14510 8128 14574 8132
rect 14590 8188 14654 8192
rect 14590 8132 14594 8188
rect 14594 8132 14650 8188
rect 14650 8132 14654 8188
rect 14590 8128 14654 8132
rect 14670 8188 14734 8192
rect 14670 8132 14674 8188
rect 14674 8132 14730 8188
rect 14730 8132 14734 8188
rect 14670 8128 14734 8132
rect 23415 8188 23479 8192
rect 23415 8132 23419 8188
rect 23419 8132 23475 8188
rect 23475 8132 23479 8188
rect 23415 8128 23479 8132
rect 23495 8188 23559 8192
rect 23495 8132 23499 8188
rect 23499 8132 23555 8188
rect 23555 8132 23559 8188
rect 23495 8128 23559 8132
rect 23575 8188 23639 8192
rect 23575 8132 23579 8188
rect 23579 8132 23635 8188
rect 23635 8132 23639 8188
rect 23575 8128 23639 8132
rect 23655 8188 23719 8192
rect 23655 8132 23659 8188
rect 23659 8132 23715 8188
rect 23715 8132 23719 8188
rect 23655 8128 23719 8132
rect 14228 7924 14292 7988
rect 22876 7924 22940 7988
rect 9937 7644 10001 7648
rect 9937 7588 9941 7644
rect 9941 7588 9997 7644
rect 9997 7588 10001 7644
rect 9937 7584 10001 7588
rect 10017 7644 10081 7648
rect 10017 7588 10021 7644
rect 10021 7588 10077 7644
rect 10077 7588 10081 7644
rect 10017 7584 10081 7588
rect 10097 7644 10161 7648
rect 10097 7588 10101 7644
rect 10101 7588 10157 7644
rect 10157 7588 10161 7644
rect 10097 7584 10161 7588
rect 10177 7644 10241 7648
rect 10177 7588 10181 7644
rect 10181 7588 10237 7644
rect 10237 7588 10241 7644
rect 10177 7584 10241 7588
rect 18922 7644 18986 7648
rect 18922 7588 18926 7644
rect 18926 7588 18982 7644
rect 18982 7588 18986 7644
rect 18922 7584 18986 7588
rect 19002 7644 19066 7648
rect 19002 7588 19006 7644
rect 19006 7588 19062 7644
rect 19062 7588 19066 7644
rect 19002 7584 19066 7588
rect 19082 7644 19146 7648
rect 19082 7588 19086 7644
rect 19086 7588 19142 7644
rect 19142 7588 19146 7644
rect 19082 7584 19146 7588
rect 19162 7644 19226 7648
rect 19162 7588 19166 7644
rect 19166 7588 19222 7644
rect 19222 7588 19226 7644
rect 19162 7584 19226 7588
rect 6868 7380 6932 7444
rect 19932 7380 19996 7444
rect 7604 7244 7668 7308
rect 17908 7244 17972 7308
rect 25268 7380 25332 7444
rect 5444 7100 5508 7104
rect 5444 7044 5448 7100
rect 5448 7044 5504 7100
rect 5504 7044 5508 7100
rect 5444 7040 5508 7044
rect 5524 7100 5588 7104
rect 5524 7044 5528 7100
rect 5528 7044 5584 7100
rect 5584 7044 5588 7100
rect 5524 7040 5588 7044
rect 5604 7100 5668 7104
rect 5604 7044 5608 7100
rect 5608 7044 5664 7100
rect 5664 7044 5668 7100
rect 5604 7040 5668 7044
rect 5684 7100 5748 7104
rect 5684 7044 5688 7100
rect 5688 7044 5744 7100
rect 5744 7044 5748 7100
rect 5684 7040 5748 7044
rect 14430 7100 14494 7104
rect 14430 7044 14434 7100
rect 14434 7044 14490 7100
rect 14490 7044 14494 7100
rect 14430 7040 14494 7044
rect 14510 7100 14574 7104
rect 14510 7044 14514 7100
rect 14514 7044 14570 7100
rect 14570 7044 14574 7100
rect 14510 7040 14574 7044
rect 14590 7100 14654 7104
rect 14590 7044 14594 7100
rect 14594 7044 14650 7100
rect 14650 7044 14654 7100
rect 14590 7040 14654 7044
rect 14670 7100 14734 7104
rect 14670 7044 14674 7100
rect 14674 7044 14730 7100
rect 14730 7044 14734 7100
rect 14670 7040 14734 7044
rect 23415 7100 23479 7104
rect 23415 7044 23419 7100
rect 23419 7044 23475 7100
rect 23475 7044 23479 7100
rect 23415 7040 23479 7044
rect 23495 7100 23559 7104
rect 23495 7044 23499 7100
rect 23499 7044 23555 7100
rect 23555 7044 23559 7100
rect 23495 7040 23559 7044
rect 23575 7100 23639 7104
rect 23575 7044 23579 7100
rect 23579 7044 23635 7100
rect 23635 7044 23639 7100
rect 23575 7040 23639 7044
rect 23655 7100 23719 7104
rect 23655 7044 23659 7100
rect 23659 7044 23715 7100
rect 23715 7044 23719 7100
rect 23655 7040 23719 7044
rect 3372 6836 3436 6900
rect 3740 6836 3804 6900
rect 9937 6556 10001 6560
rect 9937 6500 9941 6556
rect 9941 6500 9997 6556
rect 9997 6500 10001 6556
rect 9937 6496 10001 6500
rect 10017 6556 10081 6560
rect 10017 6500 10021 6556
rect 10021 6500 10077 6556
rect 10077 6500 10081 6556
rect 10017 6496 10081 6500
rect 10097 6556 10161 6560
rect 10097 6500 10101 6556
rect 10101 6500 10157 6556
rect 10157 6500 10161 6556
rect 10097 6496 10161 6500
rect 10177 6556 10241 6560
rect 10177 6500 10181 6556
rect 10181 6500 10237 6556
rect 10237 6500 10241 6556
rect 10177 6496 10241 6500
rect 18922 6556 18986 6560
rect 18922 6500 18926 6556
rect 18926 6500 18982 6556
rect 18982 6500 18986 6556
rect 18922 6496 18986 6500
rect 19002 6556 19066 6560
rect 19002 6500 19006 6556
rect 19006 6500 19062 6556
rect 19062 6500 19066 6556
rect 19002 6496 19066 6500
rect 19082 6556 19146 6560
rect 19082 6500 19086 6556
rect 19086 6500 19142 6556
rect 19142 6500 19146 6556
rect 19082 6496 19146 6500
rect 19162 6556 19226 6560
rect 19162 6500 19166 6556
rect 19166 6500 19222 6556
rect 19222 6500 19226 6556
rect 19162 6496 19226 6500
rect 25084 6488 25148 6492
rect 25084 6432 25098 6488
rect 25098 6432 25148 6488
rect 25084 6428 25148 6432
rect 27476 6428 27540 6492
rect 23796 6156 23860 6220
rect 18092 6020 18156 6084
rect 20116 6020 20180 6084
rect 5444 6012 5508 6016
rect 5444 5956 5448 6012
rect 5448 5956 5504 6012
rect 5504 5956 5508 6012
rect 5444 5952 5508 5956
rect 5524 6012 5588 6016
rect 5524 5956 5528 6012
rect 5528 5956 5584 6012
rect 5584 5956 5588 6012
rect 5524 5952 5588 5956
rect 5604 6012 5668 6016
rect 5604 5956 5608 6012
rect 5608 5956 5664 6012
rect 5664 5956 5668 6012
rect 5604 5952 5668 5956
rect 5684 6012 5748 6016
rect 5684 5956 5688 6012
rect 5688 5956 5744 6012
rect 5744 5956 5748 6012
rect 5684 5952 5748 5956
rect 14430 6012 14494 6016
rect 14430 5956 14434 6012
rect 14434 5956 14490 6012
rect 14490 5956 14494 6012
rect 14430 5952 14494 5956
rect 14510 6012 14574 6016
rect 14510 5956 14514 6012
rect 14514 5956 14570 6012
rect 14570 5956 14574 6012
rect 14510 5952 14574 5956
rect 14590 6012 14654 6016
rect 14590 5956 14594 6012
rect 14594 5956 14650 6012
rect 14650 5956 14654 6012
rect 14590 5952 14654 5956
rect 14670 6012 14734 6016
rect 14670 5956 14674 6012
rect 14674 5956 14730 6012
rect 14730 5956 14734 6012
rect 14670 5952 14734 5956
rect 23415 6012 23479 6016
rect 23415 5956 23419 6012
rect 23419 5956 23475 6012
rect 23475 5956 23479 6012
rect 23415 5952 23479 5956
rect 23495 6012 23559 6016
rect 23495 5956 23499 6012
rect 23499 5956 23555 6012
rect 23555 5956 23559 6012
rect 23495 5952 23559 5956
rect 23575 6012 23639 6016
rect 23575 5956 23579 6012
rect 23579 5956 23635 6012
rect 23635 5956 23639 6012
rect 23575 5952 23639 5956
rect 23655 6012 23719 6016
rect 23655 5956 23659 6012
rect 23659 5956 23715 6012
rect 23715 5956 23719 6012
rect 23655 5952 23719 5956
rect 21036 5944 21100 5948
rect 21036 5888 21050 5944
rect 21050 5888 21100 5944
rect 21036 5884 21100 5888
rect 22508 5944 22572 5948
rect 22508 5888 22522 5944
rect 22522 5888 22572 5944
rect 22508 5884 22572 5888
rect 3004 5672 3068 5676
rect 3004 5616 3018 5672
rect 3018 5616 3068 5672
rect 3004 5612 3068 5616
rect 3556 5612 3620 5676
rect 9937 5468 10001 5472
rect 9937 5412 9941 5468
rect 9941 5412 9997 5468
rect 9997 5412 10001 5468
rect 9937 5408 10001 5412
rect 10017 5468 10081 5472
rect 10017 5412 10021 5468
rect 10021 5412 10077 5468
rect 10077 5412 10081 5468
rect 10017 5408 10081 5412
rect 10097 5468 10161 5472
rect 10097 5412 10101 5468
rect 10101 5412 10157 5468
rect 10157 5412 10161 5468
rect 10097 5408 10161 5412
rect 10177 5468 10241 5472
rect 10177 5412 10181 5468
rect 10181 5412 10237 5468
rect 10237 5412 10241 5468
rect 10177 5408 10241 5412
rect 18276 5612 18340 5676
rect 21956 5612 22020 5676
rect 17356 5476 17420 5540
rect 20668 5476 20732 5540
rect 18922 5468 18986 5472
rect 18922 5412 18926 5468
rect 18926 5412 18982 5468
rect 18982 5412 18986 5468
rect 18922 5408 18986 5412
rect 19002 5468 19066 5472
rect 19002 5412 19006 5468
rect 19006 5412 19062 5468
rect 19062 5412 19066 5468
rect 19002 5408 19066 5412
rect 19082 5468 19146 5472
rect 19082 5412 19086 5468
rect 19086 5412 19142 5468
rect 19142 5412 19146 5468
rect 19082 5408 19146 5412
rect 19162 5468 19226 5472
rect 19162 5412 19166 5468
rect 19166 5412 19222 5468
rect 19222 5412 19226 5468
rect 19162 5408 19226 5412
rect 20484 5340 20548 5404
rect 10548 5204 10612 5268
rect 7420 5068 7484 5132
rect 5444 4924 5508 4928
rect 5444 4868 5448 4924
rect 5448 4868 5504 4924
rect 5504 4868 5508 4924
rect 5444 4864 5508 4868
rect 5524 4924 5588 4928
rect 5524 4868 5528 4924
rect 5528 4868 5584 4924
rect 5584 4868 5588 4924
rect 5524 4864 5588 4868
rect 5604 4924 5668 4928
rect 5604 4868 5608 4924
rect 5608 4868 5664 4924
rect 5664 4868 5668 4924
rect 5604 4864 5668 4868
rect 5684 4924 5748 4928
rect 5684 4868 5688 4924
rect 5688 4868 5744 4924
rect 5744 4868 5748 4924
rect 5684 4864 5748 4868
rect 14430 4924 14494 4928
rect 14430 4868 14434 4924
rect 14434 4868 14490 4924
rect 14490 4868 14494 4924
rect 14430 4864 14494 4868
rect 14510 4924 14574 4928
rect 14510 4868 14514 4924
rect 14514 4868 14570 4924
rect 14570 4868 14574 4924
rect 14510 4864 14574 4868
rect 14590 4924 14654 4928
rect 14590 4868 14594 4924
rect 14594 4868 14650 4924
rect 14650 4868 14654 4924
rect 14590 4864 14654 4868
rect 14670 4924 14734 4928
rect 14670 4868 14674 4924
rect 14674 4868 14730 4924
rect 14730 4868 14734 4924
rect 14670 4864 14734 4868
rect 23415 4924 23479 4928
rect 23415 4868 23419 4924
rect 23419 4868 23475 4924
rect 23475 4868 23479 4924
rect 23415 4864 23479 4868
rect 23495 4924 23559 4928
rect 23495 4868 23499 4924
rect 23499 4868 23555 4924
rect 23555 4868 23559 4924
rect 23495 4864 23559 4868
rect 23575 4924 23639 4928
rect 23575 4868 23579 4924
rect 23579 4868 23635 4924
rect 23635 4868 23639 4924
rect 23575 4864 23639 4868
rect 23655 4924 23719 4928
rect 23655 4868 23659 4924
rect 23659 4868 23715 4924
rect 23715 4868 23719 4924
rect 23655 4864 23719 4868
rect 7972 4720 8036 4724
rect 7972 4664 8022 4720
rect 8022 4664 8036 4720
rect 7972 4660 8036 4664
rect 3188 4388 3252 4452
rect 9937 4380 10001 4384
rect 9937 4324 9941 4380
rect 9941 4324 9997 4380
rect 9997 4324 10001 4380
rect 9937 4320 10001 4324
rect 10017 4380 10081 4384
rect 10017 4324 10021 4380
rect 10021 4324 10077 4380
rect 10077 4324 10081 4380
rect 10017 4320 10081 4324
rect 10097 4380 10161 4384
rect 10097 4324 10101 4380
rect 10101 4324 10157 4380
rect 10157 4324 10161 4380
rect 10097 4320 10161 4324
rect 10177 4380 10241 4384
rect 10177 4324 10181 4380
rect 10181 4324 10237 4380
rect 10237 4324 10241 4380
rect 10177 4320 10241 4324
rect 18922 4380 18986 4384
rect 18922 4324 18926 4380
rect 18926 4324 18982 4380
rect 18982 4324 18986 4380
rect 18922 4320 18986 4324
rect 19002 4380 19066 4384
rect 19002 4324 19006 4380
rect 19006 4324 19062 4380
rect 19062 4324 19066 4380
rect 19002 4320 19066 4324
rect 19082 4380 19146 4384
rect 19082 4324 19086 4380
rect 19086 4324 19142 4380
rect 19142 4324 19146 4380
rect 19082 4320 19146 4324
rect 19162 4380 19226 4384
rect 19162 4324 19166 4380
rect 19166 4324 19222 4380
rect 19222 4324 19226 4380
rect 19162 4320 19226 4324
rect 20116 3980 20180 4044
rect 19932 3844 19996 3908
rect 5444 3836 5508 3840
rect 5444 3780 5448 3836
rect 5448 3780 5504 3836
rect 5504 3780 5508 3836
rect 5444 3776 5508 3780
rect 5524 3836 5588 3840
rect 5524 3780 5528 3836
rect 5528 3780 5584 3836
rect 5584 3780 5588 3836
rect 5524 3776 5588 3780
rect 5604 3836 5668 3840
rect 5604 3780 5608 3836
rect 5608 3780 5664 3836
rect 5664 3780 5668 3836
rect 5604 3776 5668 3780
rect 5684 3836 5748 3840
rect 5684 3780 5688 3836
rect 5688 3780 5744 3836
rect 5744 3780 5748 3836
rect 5684 3776 5748 3780
rect 14430 3836 14494 3840
rect 14430 3780 14434 3836
rect 14434 3780 14490 3836
rect 14490 3780 14494 3836
rect 14430 3776 14494 3780
rect 14510 3836 14574 3840
rect 14510 3780 14514 3836
rect 14514 3780 14570 3836
rect 14570 3780 14574 3836
rect 14510 3776 14574 3780
rect 14590 3836 14654 3840
rect 14590 3780 14594 3836
rect 14594 3780 14650 3836
rect 14650 3780 14654 3836
rect 14590 3776 14654 3780
rect 14670 3836 14734 3840
rect 14670 3780 14674 3836
rect 14674 3780 14730 3836
rect 14730 3780 14734 3836
rect 14670 3776 14734 3780
rect 23415 3836 23479 3840
rect 23415 3780 23419 3836
rect 23419 3780 23475 3836
rect 23475 3780 23479 3836
rect 23415 3776 23479 3780
rect 23495 3836 23559 3840
rect 23495 3780 23499 3836
rect 23499 3780 23555 3836
rect 23555 3780 23559 3836
rect 23495 3776 23559 3780
rect 23575 3836 23639 3840
rect 23575 3780 23579 3836
rect 23579 3780 23635 3836
rect 23635 3780 23639 3836
rect 23575 3776 23639 3780
rect 23655 3836 23719 3840
rect 23655 3780 23659 3836
rect 23659 3780 23715 3836
rect 23715 3780 23719 3836
rect 23655 3776 23719 3780
rect 16620 3436 16684 3500
rect 9937 3292 10001 3296
rect 9937 3236 9941 3292
rect 9941 3236 9997 3292
rect 9997 3236 10001 3292
rect 9937 3232 10001 3236
rect 10017 3292 10081 3296
rect 10017 3236 10021 3292
rect 10021 3236 10077 3292
rect 10077 3236 10081 3292
rect 10017 3232 10081 3236
rect 10097 3292 10161 3296
rect 10097 3236 10101 3292
rect 10101 3236 10157 3292
rect 10157 3236 10161 3292
rect 10097 3232 10161 3236
rect 10177 3292 10241 3296
rect 10177 3236 10181 3292
rect 10181 3236 10237 3292
rect 10237 3236 10241 3292
rect 10177 3232 10241 3236
rect 18922 3292 18986 3296
rect 18922 3236 18926 3292
rect 18926 3236 18982 3292
rect 18982 3236 18986 3292
rect 18922 3232 18986 3236
rect 19002 3292 19066 3296
rect 19002 3236 19006 3292
rect 19006 3236 19062 3292
rect 19062 3236 19066 3292
rect 19002 3232 19066 3236
rect 19082 3292 19146 3296
rect 19082 3236 19086 3292
rect 19086 3236 19142 3292
rect 19142 3236 19146 3292
rect 19082 3232 19146 3236
rect 19162 3292 19226 3296
rect 19162 3236 19166 3292
rect 19166 3236 19222 3292
rect 19222 3236 19226 3292
rect 19162 3232 19226 3236
rect 18644 3164 18708 3228
rect 4108 3028 4172 3092
rect 5444 2748 5508 2752
rect 5444 2692 5448 2748
rect 5448 2692 5504 2748
rect 5504 2692 5508 2748
rect 5444 2688 5508 2692
rect 5524 2748 5588 2752
rect 5524 2692 5528 2748
rect 5528 2692 5584 2748
rect 5584 2692 5588 2748
rect 5524 2688 5588 2692
rect 5604 2748 5668 2752
rect 5604 2692 5608 2748
rect 5608 2692 5664 2748
rect 5664 2692 5668 2748
rect 5604 2688 5668 2692
rect 5684 2748 5748 2752
rect 5684 2692 5688 2748
rect 5688 2692 5744 2748
rect 5744 2692 5748 2748
rect 5684 2688 5748 2692
rect 14430 2748 14494 2752
rect 14430 2692 14434 2748
rect 14434 2692 14490 2748
rect 14490 2692 14494 2748
rect 14430 2688 14494 2692
rect 14510 2748 14574 2752
rect 14510 2692 14514 2748
rect 14514 2692 14570 2748
rect 14570 2692 14574 2748
rect 14510 2688 14574 2692
rect 14590 2748 14654 2752
rect 14590 2692 14594 2748
rect 14594 2692 14650 2748
rect 14650 2692 14654 2748
rect 14590 2688 14654 2692
rect 14670 2748 14734 2752
rect 14670 2692 14674 2748
rect 14674 2692 14730 2748
rect 14730 2692 14734 2748
rect 14670 2688 14734 2692
rect 23415 2748 23479 2752
rect 23415 2692 23419 2748
rect 23419 2692 23475 2748
rect 23475 2692 23479 2748
rect 23415 2688 23479 2692
rect 23495 2748 23559 2752
rect 23495 2692 23499 2748
rect 23499 2692 23555 2748
rect 23555 2692 23559 2748
rect 23495 2688 23559 2692
rect 23575 2748 23639 2752
rect 23575 2692 23579 2748
rect 23579 2692 23635 2748
rect 23635 2692 23639 2748
rect 23575 2688 23639 2692
rect 23655 2748 23719 2752
rect 23655 2692 23659 2748
rect 23659 2692 23715 2748
rect 23715 2692 23719 2748
rect 23655 2688 23719 2692
rect 12204 2484 12268 2548
rect 9937 2204 10001 2208
rect 9937 2148 9941 2204
rect 9941 2148 9997 2204
rect 9997 2148 10001 2204
rect 9937 2144 10001 2148
rect 10017 2204 10081 2208
rect 10017 2148 10021 2204
rect 10021 2148 10077 2204
rect 10077 2148 10081 2204
rect 10017 2144 10081 2148
rect 10097 2204 10161 2208
rect 10097 2148 10101 2204
rect 10101 2148 10157 2204
rect 10157 2148 10161 2204
rect 10097 2144 10161 2148
rect 10177 2204 10241 2208
rect 10177 2148 10181 2204
rect 10181 2148 10237 2204
rect 10237 2148 10241 2204
rect 10177 2144 10241 2148
rect 18922 2204 18986 2208
rect 18922 2148 18926 2204
rect 18926 2148 18982 2204
rect 18982 2148 18986 2204
rect 18922 2144 18986 2148
rect 19002 2204 19066 2208
rect 19002 2148 19006 2204
rect 19006 2148 19062 2204
rect 19062 2148 19066 2204
rect 19002 2144 19066 2148
rect 19082 2204 19146 2208
rect 19082 2148 19086 2204
rect 19086 2148 19142 2204
rect 19142 2148 19146 2204
rect 19082 2144 19146 2148
rect 19162 2204 19226 2208
rect 19162 2148 19166 2204
rect 19166 2148 19222 2204
rect 19222 2148 19226 2204
rect 19162 2144 19226 2148
<< metal4 >>
rect 5436 28864 5756 28880
rect 5436 28800 5444 28864
rect 5508 28800 5524 28864
rect 5588 28800 5604 28864
rect 5668 28800 5684 28864
rect 5748 28800 5756 28864
rect 5436 27776 5756 28800
rect 5436 27712 5444 27776
rect 5508 27712 5524 27776
rect 5588 27712 5604 27776
rect 5668 27712 5684 27776
rect 5748 27712 5756 27776
rect 5436 26688 5756 27712
rect 9929 28320 10250 28880
rect 9929 28256 9937 28320
rect 10001 28256 10017 28320
rect 10081 28256 10097 28320
rect 10161 28256 10177 28320
rect 10241 28256 10250 28320
rect 9929 27232 10250 28256
rect 14422 28864 14742 28880
rect 14422 28800 14430 28864
rect 14494 28800 14510 28864
rect 14574 28800 14590 28864
rect 14654 28800 14670 28864
rect 14734 28800 14742 28864
rect 14227 27980 14293 27981
rect 14227 27916 14228 27980
rect 14292 27916 14293 27980
rect 14227 27915 14293 27916
rect 12203 27708 12269 27709
rect 12203 27644 12204 27708
rect 12268 27644 12269 27708
rect 12203 27643 12269 27644
rect 9929 27168 9937 27232
rect 10001 27168 10017 27232
rect 10081 27168 10097 27232
rect 10161 27168 10177 27232
rect 10241 27168 10250 27232
rect 6499 26892 6565 26893
rect 6499 26828 6500 26892
rect 6564 26828 6565 26892
rect 6499 26827 6565 26828
rect 5436 26624 5444 26688
rect 5508 26624 5524 26688
rect 5588 26624 5604 26688
rect 5668 26624 5684 26688
rect 5748 26624 5756 26688
rect 3371 26348 3437 26349
rect 3371 26284 3372 26348
rect 3436 26284 3437 26348
rect 3371 26283 3437 26284
rect 3003 19276 3069 19277
rect 3003 19212 3004 19276
rect 3068 19212 3069 19276
rect 3003 19211 3069 19212
rect 2635 18868 2701 18869
rect 2635 18804 2636 18868
rect 2700 18804 2701 18868
rect 2635 18803 2701 18804
rect 2638 9690 2698 18803
rect 2819 18732 2885 18733
rect 2819 18668 2820 18732
rect 2884 18668 2885 18732
rect 2819 18667 2885 18668
rect 2822 17781 2882 18667
rect 2819 17780 2885 17781
rect 2819 17716 2820 17780
rect 2884 17716 2885 17780
rect 2819 17715 2885 17716
rect 2819 16284 2885 16285
rect 2819 16220 2820 16284
rect 2884 16220 2885 16284
rect 2819 16219 2885 16220
rect 2822 10029 2882 16219
rect 3006 12477 3066 19211
rect 3187 18732 3253 18733
rect 3187 18668 3188 18732
rect 3252 18668 3253 18732
rect 3187 18667 3253 18668
rect 3190 13565 3250 18667
rect 3187 13564 3253 13565
rect 3187 13500 3188 13564
rect 3252 13500 3253 13564
rect 3187 13499 3253 13500
rect 3187 12884 3253 12885
rect 3187 12820 3188 12884
rect 3252 12820 3253 12884
rect 3187 12819 3253 12820
rect 3003 12476 3069 12477
rect 3003 12412 3004 12476
rect 3068 12412 3069 12476
rect 3003 12411 3069 12412
rect 3003 12068 3069 12069
rect 3003 12004 3004 12068
rect 3068 12004 3069 12068
rect 3003 12003 3069 12004
rect 2819 10028 2885 10029
rect 2819 9964 2820 10028
rect 2884 9964 2885 10028
rect 2819 9963 2885 9964
rect 2638 9630 2882 9690
rect 2822 8533 2882 9630
rect 2819 8532 2885 8533
rect 2819 8468 2820 8532
rect 2884 8468 2885 8532
rect 2819 8467 2885 8468
rect 3006 5677 3066 12003
rect 3003 5676 3069 5677
rect 3003 5612 3004 5676
rect 3068 5612 3069 5676
rect 3003 5611 3069 5612
rect 3190 4453 3250 12819
rect 3374 6901 3434 26283
rect 5436 25600 5756 26624
rect 5436 25536 5444 25600
rect 5508 25536 5524 25600
rect 5588 25536 5604 25600
rect 5668 25536 5684 25600
rect 5748 25536 5756 25600
rect 5436 24512 5756 25536
rect 5436 24448 5444 24512
rect 5508 24448 5524 24512
rect 5588 24448 5604 24512
rect 5668 24448 5684 24512
rect 5748 24448 5756 24512
rect 5436 23424 5756 24448
rect 5436 23360 5444 23424
rect 5508 23360 5524 23424
rect 5588 23360 5604 23424
rect 5668 23360 5684 23424
rect 5748 23360 5756 23424
rect 4475 22948 4541 22949
rect 4475 22884 4476 22948
rect 4540 22884 4541 22948
rect 4475 22883 4541 22884
rect 4107 22676 4173 22677
rect 4107 22612 4108 22676
rect 4172 22612 4173 22676
rect 4107 22611 4173 22612
rect 3555 20364 3621 20365
rect 3555 20300 3556 20364
rect 3620 20300 3621 20364
rect 3555 20299 3621 20300
rect 3558 13973 3618 20299
rect 3923 18596 3989 18597
rect 3923 18532 3924 18596
rect 3988 18532 3989 18596
rect 3923 18531 3989 18532
rect 3739 15740 3805 15741
rect 3739 15676 3740 15740
rect 3804 15676 3805 15740
rect 3739 15675 3805 15676
rect 3555 13972 3621 13973
rect 3555 13908 3556 13972
rect 3620 13908 3621 13972
rect 3555 13907 3621 13908
rect 3555 13020 3621 13021
rect 3555 12956 3556 13020
rect 3620 12956 3621 13020
rect 3555 12955 3621 12956
rect 3371 6900 3437 6901
rect 3371 6836 3372 6900
rect 3436 6836 3437 6900
rect 3371 6835 3437 6836
rect 3558 5677 3618 12955
rect 3742 10165 3802 15675
rect 3926 14381 3986 18531
rect 3923 14380 3989 14381
rect 3923 14316 3924 14380
rect 3988 14316 3989 14380
rect 3923 14315 3989 14316
rect 4110 14242 4170 22611
rect 4291 18324 4357 18325
rect 4291 18260 4292 18324
rect 4356 18260 4357 18324
rect 4291 18259 4357 18260
rect 3926 14182 4170 14242
rect 3926 11661 3986 14182
rect 4107 13700 4173 13701
rect 4107 13636 4108 13700
rect 4172 13636 4173 13700
rect 4107 13635 4173 13636
rect 3923 11660 3989 11661
rect 3923 11596 3924 11660
rect 3988 11596 3989 11660
rect 3923 11595 3989 11596
rect 3739 10164 3805 10165
rect 3739 10100 3740 10164
rect 3804 10100 3805 10164
rect 3739 10099 3805 10100
rect 3739 8532 3805 8533
rect 3739 8468 3740 8532
rect 3804 8468 3805 8532
rect 3739 8467 3805 8468
rect 3742 6901 3802 8467
rect 3739 6900 3805 6901
rect 3739 6836 3740 6900
rect 3804 6836 3805 6900
rect 3739 6835 3805 6836
rect 3555 5676 3621 5677
rect 3555 5612 3556 5676
rect 3620 5612 3621 5676
rect 3555 5611 3621 5612
rect 3187 4452 3253 4453
rect 3187 4388 3188 4452
rect 3252 4388 3253 4452
rect 3187 4387 3253 4388
rect 4110 3093 4170 13635
rect 4294 12069 4354 18259
rect 4478 12749 4538 22883
rect 4843 22540 4909 22541
rect 4843 22476 4844 22540
rect 4908 22476 4909 22540
rect 4843 22475 4909 22476
rect 5211 22540 5277 22541
rect 5211 22476 5212 22540
rect 5276 22476 5277 22540
rect 5211 22475 5277 22476
rect 4846 20637 4906 22475
rect 5214 21453 5274 22475
rect 5436 22336 5756 23360
rect 5436 22272 5444 22336
rect 5508 22272 5524 22336
rect 5588 22272 5604 22336
rect 5668 22272 5684 22336
rect 5748 22272 5756 22336
rect 5211 21452 5277 21453
rect 5211 21388 5212 21452
rect 5276 21388 5277 21452
rect 5211 21387 5277 21388
rect 5211 21316 5277 21317
rect 5211 21252 5212 21316
rect 5276 21252 5277 21316
rect 5211 21251 5277 21252
rect 4843 20636 4909 20637
rect 4843 20572 4844 20636
rect 4908 20572 4909 20636
rect 4843 20571 4909 20572
rect 4659 19004 4725 19005
rect 4659 18940 4660 19004
rect 4724 18940 4725 19004
rect 4659 18939 4725 18940
rect 4662 13021 4722 18939
rect 5214 18461 5274 21251
rect 5436 21248 5756 22272
rect 6315 21860 6381 21861
rect 6315 21796 6316 21860
rect 6380 21796 6381 21860
rect 6315 21795 6381 21796
rect 5436 21184 5444 21248
rect 5508 21184 5524 21248
rect 5588 21184 5604 21248
rect 5668 21184 5684 21248
rect 5748 21184 5756 21248
rect 5436 20160 5756 21184
rect 6131 21044 6197 21045
rect 6131 20980 6132 21044
rect 6196 20980 6197 21044
rect 6131 20979 6197 20980
rect 5436 20096 5444 20160
rect 5508 20096 5524 20160
rect 5588 20096 5604 20160
rect 5668 20096 5684 20160
rect 5748 20096 5756 20160
rect 5436 19072 5756 20096
rect 5947 19684 6013 19685
rect 5947 19620 5948 19684
rect 6012 19620 6013 19684
rect 5947 19619 6013 19620
rect 5436 19008 5444 19072
rect 5508 19008 5524 19072
rect 5588 19008 5604 19072
rect 5668 19008 5684 19072
rect 5748 19008 5756 19072
rect 5211 18460 5277 18461
rect 5211 18396 5212 18460
rect 5276 18396 5277 18460
rect 5211 18395 5277 18396
rect 5027 18188 5093 18189
rect 5027 18124 5028 18188
rect 5092 18124 5093 18188
rect 5027 18123 5093 18124
rect 5211 18188 5277 18189
rect 5211 18124 5212 18188
rect 5276 18124 5277 18188
rect 5211 18123 5277 18124
rect 4843 17644 4909 17645
rect 4843 17580 4844 17644
rect 4908 17580 4909 17644
rect 4843 17579 4909 17580
rect 4659 13020 4725 13021
rect 4659 12956 4660 13020
rect 4724 12956 4725 13020
rect 4659 12955 4725 12956
rect 4659 12884 4725 12885
rect 4659 12820 4660 12884
rect 4724 12820 4725 12884
rect 4659 12819 4725 12820
rect 4475 12748 4541 12749
rect 4475 12684 4476 12748
rect 4540 12684 4541 12748
rect 4475 12683 4541 12684
rect 4475 12612 4541 12613
rect 4475 12548 4476 12612
rect 4540 12548 4541 12612
rect 4475 12547 4541 12548
rect 4478 12341 4538 12547
rect 4475 12340 4541 12341
rect 4475 12276 4476 12340
rect 4540 12276 4541 12340
rect 4475 12275 4541 12276
rect 4662 12069 4722 12819
rect 4846 12477 4906 17579
rect 4843 12476 4909 12477
rect 4843 12412 4844 12476
rect 4908 12412 4909 12476
rect 4843 12411 4909 12412
rect 4291 12068 4357 12069
rect 4291 12004 4292 12068
rect 4356 12004 4357 12068
rect 4291 12003 4357 12004
rect 4659 12068 4725 12069
rect 4659 12004 4660 12068
rect 4724 12004 4725 12068
rect 4659 12003 4725 12004
rect 5030 9757 5090 18123
rect 5214 13293 5274 18123
rect 5436 17984 5756 19008
rect 5950 19005 6010 19619
rect 5947 19004 6013 19005
rect 5947 18940 5948 19004
rect 6012 18940 6013 19004
rect 5947 18939 6013 18940
rect 5947 18596 6013 18597
rect 5947 18532 5948 18596
rect 6012 18532 6013 18596
rect 5947 18531 6013 18532
rect 5436 17920 5444 17984
rect 5508 17920 5524 17984
rect 5588 17920 5604 17984
rect 5668 17920 5684 17984
rect 5748 17920 5756 17984
rect 5436 16896 5756 17920
rect 5436 16832 5444 16896
rect 5508 16832 5524 16896
rect 5588 16832 5604 16896
rect 5668 16832 5684 16896
rect 5748 16832 5756 16896
rect 5436 15808 5756 16832
rect 5436 15744 5444 15808
rect 5508 15744 5524 15808
rect 5588 15744 5604 15808
rect 5668 15744 5684 15808
rect 5748 15744 5756 15808
rect 5436 14720 5756 15744
rect 5436 14656 5444 14720
rect 5508 14656 5524 14720
rect 5588 14656 5604 14720
rect 5668 14656 5684 14720
rect 5748 14656 5756 14720
rect 5436 13632 5756 14656
rect 5436 13568 5444 13632
rect 5508 13568 5524 13632
rect 5588 13568 5604 13632
rect 5668 13568 5684 13632
rect 5748 13568 5756 13632
rect 5211 13292 5277 13293
rect 5211 13228 5212 13292
rect 5276 13228 5277 13292
rect 5211 13227 5277 13228
rect 5211 12612 5277 12613
rect 5211 12548 5212 12612
rect 5276 12548 5277 12612
rect 5211 12547 5277 12548
rect 5214 9893 5274 12547
rect 5436 12544 5756 13568
rect 5436 12480 5444 12544
rect 5508 12480 5524 12544
rect 5588 12480 5604 12544
rect 5668 12480 5684 12544
rect 5748 12480 5756 12544
rect 5436 11456 5756 12480
rect 5950 11933 6010 18531
rect 5947 11932 6013 11933
rect 5947 11868 5948 11932
rect 6012 11868 6013 11932
rect 5947 11867 6013 11868
rect 5436 11392 5444 11456
rect 5508 11392 5524 11456
rect 5588 11392 5604 11456
rect 5668 11392 5684 11456
rect 5748 11392 5756 11456
rect 5436 10368 5756 11392
rect 5436 10304 5444 10368
rect 5508 10304 5524 10368
rect 5588 10304 5604 10368
rect 5668 10304 5684 10368
rect 5748 10304 5756 10368
rect 5211 9892 5277 9893
rect 5211 9828 5212 9892
rect 5276 9828 5277 9892
rect 5211 9827 5277 9828
rect 5027 9756 5093 9757
rect 5027 9692 5028 9756
rect 5092 9692 5093 9756
rect 5027 9691 5093 9692
rect 5436 9280 5756 10304
rect 6134 10029 6194 20979
rect 6318 18597 6378 21795
rect 6315 18596 6381 18597
rect 6315 18532 6316 18596
rect 6380 18532 6381 18596
rect 6315 18531 6381 18532
rect 6502 18325 6562 26827
rect 9929 26144 10250 27168
rect 11467 26484 11533 26485
rect 11467 26420 11468 26484
rect 11532 26420 11533 26484
rect 11467 26419 11533 26420
rect 9929 26080 9937 26144
rect 10001 26080 10017 26144
rect 10081 26080 10097 26144
rect 10161 26080 10177 26144
rect 10241 26080 10250 26144
rect 9929 25056 10250 26080
rect 9929 24992 9937 25056
rect 10001 24992 10017 25056
rect 10081 24992 10097 25056
rect 10161 24992 10177 25056
rect 10241 24992 10250 25056
rect 9929 23968 10250 24992
rect 9929 23904 9937 23968
rect 10001 23904 10017 23968
rect 10081 23904 10097 23968
rect 10161 23904 10177 23968
rect 10241 23904 10250 23968
rect 9929 22880 10250 23904
rect 9929 22816 9937 22880
rect 10001 22816 10017 22880
rect 10081 22816 10097 22880
rect 10161 22816 10177 22880
rect 10241 22816 10250 22880
rect 9929 21792 10250 22816
rect 9929 21728 9937 21792
rect 10001 21728 10017 21792
rect 10081 21728 10097 21792
rect 10161 21728 10177 21792
rect 10241 21728 10250 21792
rect 7235 21452 7301 21453
rect 7235 21388 7236 21452
rect 7300 21388 7301 21452
rect 7235 21387 7301 21388
rect 6499 18324 6565 18325
rect 6499 18260 6500 18324
rect 6564 18260 6565 18324
rect 6499 18259 6565 18260
rect 7051 17372 7117 17373
rect 7051 17308 7052 17372
rect 7116 17308 7117 17372
rect 7051 17307 7117 17308
rect 6683 15604 6749 15605
rect 6683 15540 6684 15604
rect 6748 15540 6749 15604
rect 6683 15539 6749 15540
rect 6315 15332 6381 15333
rect 6315 15268 6316 15332
rect 6380 15268 6381 15332
rect 6315 15267 6381 15268
rect 6318 10981 6378 15267
rect 6499 12612 6565 12613
rect 6499 12548 6500 12612
rect 6564 12548 6565 12612
rect 6499 12547 6565 12548
rect 6502 12341 6562 12547
rect 6499 12340 6565 12341
rect 6499 12276 6500 12340
rect 6564 12276 6565 12340
rect 6499 12275 6565 12276
rect 6686 12069 6746 15539
rect 7054 12477 7114 17307
rect 7238 12477 7298 21387
rect 9627 20908 9693 20909
rect 9627 20844 9628 20908
rect 9692 20844 9693 20908
rect 9627 20843 9693 20844
rect 9259 20772 9325 20773
rect 9259 20708 9260 20772
rect 9324 20708 9325 20772
rect 9259 20707 9325 20708
rect 7971 20500 8037 20501
rect 7971 20436 7972 20500
rect 8036 20436 8037 20500
rect 7971 20435 8037 20436
rect 7787 19956 7853 19957
rect 7787 19892 7788 19956
rect 7852 19892 7853 19956
rect 7787 19891 7853 19892
rect 7790 18461 7850 19891
rect 7787 18460 7853 18461
rect 7787 18396 7788 18460
rect 7852 18396 7853 18460
rect 7787 18395 7853 18396
rect 7419 17100 7485 17101
rect 7419 17036 7420 17100
rect 7484 17036 7485 17100
rect 7419 17035 7485 17036
rect 7051 12476 7117 12477
rect 7051 12412 7052 12476
rect 7116 12412 7117 12476
rect 7051 12411 7117 12412
rect 7235 12476 7301 12477
rect 7235 12412 7236 12476
rect 7300 12412 7301 12476
rect 7422 12474 7482 17035
rect 7974 12749 8034 20435
rect 8155 19956 8221 19957
rect 8155 19892 8156 19956
rect 8220 19892 8221 19956
rect 8155 19891 8221 19892
rect 8158 19413 8218 19891
rect 8155 19412 8221 19413
rect 8155 19348 8156 19412
rect 8220 19348 8221 19412
rect 8155 19347 8221 19348
rect 8155 19140 8221 19141
rect 8155 19076 8156 19140
rect 8220 19076 8221 19140
rect 8155 19075 8221 19076
rect 7787 12748 7853 12749
rect 7787 12684 7788 12748
rect 7852 12684 7853 12748
rect 7787 12683 7853 12684
rect 7971 12748 8037 12749
rect 7971 12684 7972 12748
rect 8036 12684 8037 12748
rect 7971 12683 8037 12684
rect 7422 12414 7666 12474
rect 7235 12411 7301 12412
rect 6867 12340 6933 12341
rect 6867 12276 6868 12340
rect 6932 12276 6933 12340
rect 6867 12275 6933 12276
rect 7051 12340 7117 12341
rect 7051 12276 7052 12340
rect 7116 12276 7117 12340
rect 7051 12275 7117 12276
rect 7419 12340 7485 12341
rect 7419 12276 7420 12340
rect 7484 12276 7485 12340
rect 7419 12275 7485 12276
rect 6683 12068 6749 12069
rect 6683 12004 6684 12068
rect 6748 12004 6749 12068
rect 6683 12003 6749 12004
rect 6315 10980 6381 10981
rect 6315 10916 6316 10980
rect 6380 10916 6381 10980
rect 6315 10915 6381 10916
rect 6131 10028 6197 10029
rect 6131 9964 6132 10028
rect 6196 9964 6197 10028
rect 6131 9963 6197 9964
rect 5436 9216 5444 9280
rect 5508 9216 5524 9280
rect 5588 9216 5604 9280
rect 5668 9216 5684 9280
rect 5748 9216 5756 9280
rect 5436 8192 5756 9216
rect 5436 8128 5444 8192
rect 5508 8128 5524 8192
rect 5588 8128 5604 8192
rect 5668 8128 5684 8192
rect 5748 8128 5756 8192
rect 5436 7104 5756 8128
rect 6870 7445 6930 12275
rect 7054 10029 7114 12275
rect 7051 10028 7117 10029
rect 7051 9964 7052 10028
rect 7116 9964 7117 10028
rect 7051 9963 7117 9964
rect 6867 7444 6933 7445
rect 6867 7380 6868 7444
rect 6932 7380 6933 7444
rect 6867 7379 6933 7380
rect 5436 7040 5444 7104
rect 5508 7040 5524 7104
rect 5588 7040 5604 7104
rect 5668 7040 5684 7104
rect 5748 7040 5756 7104
rect 5436 6016 5756 7040
rect 5436 5952 5444 6016
rect 5508 5952 5524 6016
rect 5588 5952 5604 6016
rect 5668 5952 5684 6016
rect 5748 5952 5756 6016
rect 5436 4928 5756 5952
rect 7422 5133 7482 12275
rect 7606 12069 7666 12414
rect 7790 12341 7850 12683
rect 7787 12340 7853 12341
rect 7787 12276 7788 12340
rect 7852 12276 7853 12340
rect 7787 12275 7853 12276
rect 7603 12068 7669 12069
rect 7603 12004 7604 12068
rect 7668 12004 7669 12068
rect 7603 12003 7669 12004
rect 7603 11116 7669 11117
rect 7603 11052 7604 11116
rect 7668 11052 7669 11116
rect 7603 11051 7669 11052
rect 7606 7309 7666 11051
rect 8158 10845 8218 19075
rect 9075 14788 9141 14789
rect 9075 14724 9076 14788
rect 9140 14724 9141 14788
rect 9075 14723 9141 14724
rect 8707 13292 8773 13293
rect 8707 13228 8708 13292
rect 8772 13228 8773 13292
rect 8707 13227 8773 13228
rect 8523 12884 8589 12885
rect 8523 12820 8524 12884
rect 8588 12820 8589 12884
rect 8523 12819 8589 12820
rect 8526 12341 8586 12819
rect 8710 12613 8770 13227
rect 8707 12612 8773 12613
rect 8707 12548 8708 12612
rect 8772 12548 8773 12612
rect 8707 12547 8773 12548
rect 8523 12340 8589 12341
rect 8523 12276 8524 12340
rect 8588 12276 8589 12340
rect 8523 12275 8589 12276
rect 9078 11253 9138 14723
rect 9262 12477 9322 20707
rect 9630 19005 9690 20843
rect 9929 20704 10250 21728
rect 11283 20908 11349 20909
rect 11283 20844 11284 20908
rect 11348 20844 11349 20908
rect 11283 20843 11349 20844
rect 9929 20640 9937 20704
rect 10001 20640 10017 20704
rect 10081 20640 10097 20704
rect 10161 20640 10177 20704
rect 10241 20640 10250 20704
rect 9929 19616 10250 20640
rect 9929 19552 9937 19616
rect 10001 19552 10017 19616
rect 10081 19552 10097 19616
rect 10161 19552 10177 19616
rect 10241 19552 10250 19616
rect 9627 19004 9693 19005
rect 9627 18940 9628 19004
rect 9692 18940 9693 19004
rect 9627 18939 9693 18940
rect 9929 18528 10250 19552
rect 11099 19276 11165 19277
rect 11099 19212 11100 19276
rect 11164 19212 11165 19276
rect 11099 19211 11165 19212
rect 10731 18868 10797 18869
rect 10731 18804 10732 18868
rect 10796 18804 10797 18868
rect 10731 18803 10797 18804
rect 9929 18464 9937 18528
rect 10001 18464 10017 18528
rect 10081 18464 10097 18528
rect 10161 18464 10177 18528
rect 10241 18464 10250 18528
rect 9929 17440 10250 18464
rect 10363 18188 10429 18189
rect 10363 18124 10364 18188
rect 10428 18124 10429 18188
rect 10363 18123 10429 18124
rect 9929 17376 9937 17440
rect 10001 17376 10017 17440
rect 10081 17376 10097 17440
rect 10161 17376 10177 17440
rect 10241 17376 10250 17440
rect 9929 16352 10250 17376
rect 9929 16288 9937 16352
rect 10001 16288 10017 16352
rect 10081 16288 10097 16352
rect 10161 16288 10177 16352
rect 10241 16288 10250 16352
rect 9929 15264 10250 16288
rect 9929 15200 9937 15264
rect 10001 15200 10017 15264
rect 10081 15200 10097 15264
rect 10161 15200 10177 15264
rect 10241 15200 10250 15264
rect 9929 14176 10250 15200
rect 9929 14112 9937 14176
rect 10001 14112 10017 14176
rect 10081 14112 10097 14176
rect 10161 14112 10177 14176
rect 10241 14112 10250 14176
rect 9443 13156 9509 13157
rect 9443 13092 9444 13156
rect 9508 13092 9509 13156
rect 9443 13091 9509 13092
rect 9259 12476 9325 12477
rect 9259 12412 9260 12476
rect 9324 12412 9325 12476
rect 9259 12411 9325 12412
rect 9446 11797 9506 13091
rect 9929 13088 10250 14112
rect 9929 13024 9937 13088
rect 10001 13024 10017 13088
rect 10081 13024 10097 13088
rect 10161 13024 10177 13088
rect 10241 13024 10250 13088
rect 9929 12000 10250 13024
rect 9929 11936 9937 12000
rect 10001 11936 10017 12000
rect 10081 11936 10097 12000
rect 10161 11936 10177 12000
rect 10241 11936 10250 12000
rect 9443 11796 9509 11797
rect 9443 11732 9444 11796
rect 9508 11732 9509 11796
rect 9443 11731 9509 11732
rect 9075 11252 9141 11253
rect 9075 11188 9076 11252
rect 9140 11188 9141 11252
rect 9075 11187 9141 11188
rect 9929 10912 10250 11936
rect 9929 10848 9937 10912
rect 10001 10848 10017 10912
rect 10081 10848 10097 10912
rect 10161 10848 10177 10912
rect 10241 10848 10250 10912
rect 8155 10844 8221 10845
rect 8155 10780 8156 10844
rect 8220 10780 8221 10844
rect 8155 10779 8221 10780
rect 9259 10164 9325 10165
rect 9259 10100 9260 10164
rect 9324 10100 9325 10164
rect 9259 10099 9325 10100
rect 7971 9892 8037 9893
rect 7971 9828 7972 9892
rect 8036 9828 8037 9892
rect 7971 9827 8037 9828
rect 7603 7308 7669 7309
rect 7603 7244 7604 7308
rect 7668 7244 7669 7308
rect 7603 7243 7669 7244
rect 7419 5132 7485 5133
rect 7419 5068 7420 5132
rect 7484 5068 7485 5132
rect 7419 5067 7485 5068
rect 5436 4864 5444 4928
rect 5508 4864 5524 4928
rect 5588 4864 5604 4928
rect 5668 4864 5684 4928
rect 5748 4864 5756 4928
rect 5436 3840 5756 4864
rect 7974 4725 8034 9827
rect 9262 8533 9322 10099
rect 9929 9824 10250 10848
rect 10366 10573 10426 18123
rect 10547 17916 10613 17917
rect 10547 17852 10548 17916
rect 10612 17852 10613 17916
rect 10547 17851 10613 17852
rect 10363 10572 10429 10573
rect 10363 10508 10364 10572
rect 10428 10508 10429 10572
rect 10363 10507 10429 10508
rect 10363 9892 10429 9893
rect 10363 9828 10364 9892
rect 10428 9828 10429 9892
rect 10363 9827 10429 9828
rect 9929 9760 9937 9824
rect 10001 9760 10017 9824
rect 10081 9760 10097 9824
rect 10161 9760 10177 9824
rect 10241 9760 10250 9824
rect 9929 8736 10250 9760
rect 9929 8672 9937 8736
rect 10001 8672 10017 8736
rect 10081 8672 10097 8736
rect 10161 8672 10177 8736
rect 10241 8672 10250 8736
rect 9259 8532 9325 8533
rect 9259 8468 9260 8532
rect 9324 8468 9325 8532
rect 9259 8467 9325 8468
rect 9929 7648 10250 8672
rect 10366 8397 10426 9827
rect 10363 8396 10429 8397
rect 10363 8332 10364 8396
rect 10428 8332 10429 8396
rect 10363 8331 10429 8332
rect 9929 7584 9937 7648
rect 10001 7584 10017 7648
rect 10081 7584 10097 7648
rect 10161 7584 10177 7648
rect 10241 7584 10250 7648
rect 9929 6560 10250 7584
rect 9929 6496 9937 6560
rect 10001 6496 10017 6560
rect 10081 6496 10097 6560
rect 10161 6496 10177 6560
rect 10241 6496 10250 6560
rect 9929 5472 10250 6496
rect 9929 5408 9937 5472
rect 10001 5408 10017 5472
rect 10081 5408 10097 5472
rect 10161 5408 10177 5472
rect 10241 5408 10250 5472
rect 7971 4724 8037 4725
rect 7971 4660 7972 4724
rect 8036 4660 8037 4724
rect 7971 4659 8037 4660
rect 5436 3776 5444 3840
rect 5508 3776 5524 3840
rect 5588 3776 5604 3840
rect 5668 3776 5684 3840
rect 5748 3776 5756 3840
rect 4107 3092 4173 3093
rect 4107 3028 4108 3092
rect 4172 3028 4173 3092
rect 4107 3027 4173 3028
rect 5436 2752 5756 3776
rect 5436 2688 5444 2752
rect 5508 2688 5524 2752
rect 5588 2688 5604 2752
rect 5668 2688 5684 2752
rect 5748 2688 5756 2752
rect 5436 2128 5756 2688
rect 9929 4384 10250 5408
rect 10550 5269 10610 17851
rect 10734 12205 10794 18803
rect 10915 18460 10981 18461
rect 10915 18396 10916 18460
rect 10980 18396 10981 18460
rect 10915 18395 10981 18396
rect 10918 12341 10978 18395
rect 10915 12340 10981 12341
rect 10915 12276 10916 12340
rect 10980 12276 10981 12340
rect 10915 12275 10981 12276
rect 10731 12204 10797 12205
rect 10731 12140 10732 12204
rect 10796 12140 10797 12204
rect 10731 12139 10797 12140
rect 11102 9757 11162 19211
rect 11286 14245 11346 20843
rect 11470 18053 11530 26419
rect 12019 19004 12085 19005
rect 12019 18940 12020 19004
rect 12084 18940 12085 19004
rect 12019 18939 12085 18940
rect 11467 18052 11533 18053
rect 11467 17988 11468 18052
rect 11532 17988 11533 18052
rect 11467 17987 11533 17988
rect 11467 17508 11533 17509
rect 11467 17444 11468 17508
rect 11532 17444 11533 17508
rect 11467 17443 11533 17444
rect 11283 14244 11349 14245
rect 11283 14180 11284 14244
rect 11348 14180 11349 14244
rect 11283 14179 11349 14180
rect 11099 9756 11165 9757
rect 11099 9692 11100 9756
rect 11164 9692 11165 9756
rect 11099 9691 11165 9692
rect 11470 8397 11530 17443
rect 11835 17100 11901 17101
rect 11835 17036 11836 17100
rect 11900 17036 11901 17100
rect 11835 17035 11901 17036
rect 11651 14924 11717 14925
rect 11651 14860 11652 14924
rect 11716 14860 11717 14924
rect 11651 14859 11717 14860
rect 11654 13973 11714 14859
rect 11651 13972 11717 13973
rect 11651 13908 11652 13972
rect 11716 13908 11717 13972
rect 11651 13907 11717 13908
rect 11838 10981 11898 17035
rect 12022 11797 12082 18939
rect 12019 11796 12085 11797
rect 12019 11732 12020 11796
rect 12084 11732 12085 11796
rect 12019 11731 12085 11732
rect 11835 10980 11901 10981
rect 11835 10916 11836 10980
rect 11900 10916 11901 10980
rect 11835 10915 11901 10916
rect 11467 8396 11533 8397
rect 11467 8332 11468 8396
rect 11532 8332 11533 8396
rect 11467 8331 11533 8332
rect 10547 5268 10613 5269
rect 10547 5204 10548 5268
rect 10612 5204 10613 5268
rect 10547 5203 10613 5204
rect 9929 4320 9937 4384
rect 10001 4320 10017 4384
rect 10081 4320 10097 4384
rect 10161 4320 10177 4384
rect 10241 4320 10250 4384
rect 9929 3296 10250 4320
rect 9929 3232 9937 3296
rect 10001 3232 10017 3296
rect 10081 3232 10097 3296
rect 10161 3232 10177 3296
rect 10241 3232 10250 3296
rect 9929 2208 10250 3232
rect 12206 2549 12266 27643
rect 13675 21044 13741 21045
rect 13675 20980 13676 21044
rect 13740 20980 13741 21044
rect 13675 20979 13741 20980
rect 14043 21044 14109 21045
rect 14043 20980 14044 21044
rect 14108 20980 14109 21044
rect 14043 20979 14109 20980
rect 13491 20092 13557 20093
rect 13491 20028 13492 20092
rect 13556 20028 13557 20092
rect 13491 20027 13557 20028
rect 13494 19549 13554 20027
rect 13491 19548 13557 19549
rect 13491 19484 13492 19548
rect 13556 19484 13557 19548
rect 13491 19483 13557 19484
rect 13678 18189 13738 20979
rect 13675 18188 13741 18189
rect 13675 18124 13676 18188
rect 13740 18124 13741 18188
rect 13675 18123 13741 18124
rect 13491 17780 13557 17781
rect 13491 17716 13492 17780
rect 13556 17716 13557 17780
rect 13491 17715 13557 17716
rect 13494 14381 13554 17715
rect 14046 17237 14106 20979
rect 14043 17236 14109 17237
rect 14043 17172 14044 17236
rect 14108 17172 14109 17236
rect 14043 17171 14109 17172
rect 13491 14380 13557 14381
rect 13491 14316 13492 14380
rect 13556 14316 13557 14380
rect 13491 14315 13557 14316
rect 14043 12068 14109 12069
rect 14043 12004 14044 12068
rect 14108 12004 14109 12068
rect 14043 12003 14109 12004
rect 14046 9893 14106 12003
rect 14043 9892 14109 9893
rect 14043 9828 14044 9892
rect 14108 9828 14109 9892
rect 14043 9827 14109 9828
rect 14230 7989 14290 27915
rect 14422 27776 14742 28800
rect 14422 27712 14430 27776
rect 14494 27712 14510 27776
rect 14574 27712 14590 27776
rect 14654 27712 14670 27776
rect 14734 27712 14742 27776
rect 14422 26688 14742 27712
rect 14422 26624 14430 26688
rect 14494 26624 14510 26688
rect 14574 26624 14590 26688
rect 14654 26624 14670 26688
rect 14734 26624 14742 26688
rect 14422 25600 14742 26624
rect 18914 28320 19235 28880
rect 18914 28256 18922 28320
rect 18986 28256 19002 28320
rect 19066 28256 19082 28320
rect 19146 28256 19162 28320
rect 19226 28256 19235 28320
rect 18914 27232 19235 28256
rect 18914 27168 18922 27232
rect 18986 27168 19002 27232
rect 19066 27168 19082 27232
rect 19146 27168 19162 27232
rect 19226 27168 19235 27232
rect 15331 26348 15397 26349
rect 15331 26284 15332 26348
rect 15396 26284 15397 26348
rect 15331 26283 15397 26284
rect 18275 26348 18341 26349
rect 18275 26284 18276 26348
rect 18340 26284 18341 26348
rect 18275 26283 18341 26284
rect 14422 25536 14430 25600
rect 14494 25536 14510 25600
rect 14574 25536 14590 25600
rect 14654 25536 14670 25600
rect 14734 25536 14742 25600
rect 14422 24512 14742 25536
rect 14422 24448 14430 24512
rect 14494 24448 14510 24512
rect 14574 24448 14590 24512
rect 14654 24448 14670 24512
rect 14734 24448 14742 24512
rect 14422 23424 14742 24448
rect 14422 23360 14430 23424
rect 14494 23360 14510 23424
rect 14574 23360 14590 23424
rect 14654 23360 14670 23424
rect 14734 23360 14742 23424
rect 14422 22336 14742 23360
rect 14422 22272 14430 22336
rect 14494 22272 14510 22336
rect 14574 22272 14590 22336
rect 14654 22272 14670 22336
rect 14734 22272 14742 22336
rect 14422 21248 14742 22272
rect 14963 21452 15029 21453
rect 14963 21388 14964 21452
rect 15028 21388 15029 21452
rect 14963 21387 15029 21388
rect 14422 21184 14430 21248
rect 14494 21184 14510 21248
rect 14574 21184 14590 21248
rect 14654 21184 14670 21248
rect 14734 21184 14742 21248
rect 14422 20160 14742 21184
rect 14422 20096 14430 20160
rect 14494 20096 14510 20160
rect 14574 20096 14590 20160
rect 14654 20096 14670 20160
rect 14734 20096 14742 20160
rect 14422 19072 14742 20096
rect 14422 19008 14430 19072
rect 14494 19008 14510 19072
rect 14574 19008 14590 19072
rect 14654 19008 14670 19072
rect 14734 19008 14742 19072
rect 14422 17984 14742 19008
rect 14422 17920 14430 17984
rect 14494 17920 14510 17984
rect 14574 17920 14590 17984
rect 14654 17920 14670 17984
rect 14734 17920 14742 17984
rect 14422 16896 14742 17920
rect 14422 16832 14430 16896
rect 14494 16832 14510 16896
rect 14574 16832 14590 16896
rect 14654 16832 14670 16896
rect 14734 16832 14742 16896
rect 14422 15808 14742 16832
rect 14422 15744 14430 15808
rect 14494 15744 14510 15808
rect 14574 15744 14590 15808
rect 14654 15744 14670 15808
rect 14734 15744 14742 15808
rect 14422 14720 14742 15744
rect 14422 14656 14430 14720
rect 14494 14656 14510 14720
rect 14574 14656 14590 14720
rect 14654 14656 14670 14720
rect 14734 14656 14742 14720
rect 14422 13632 14742 14656
rect 14422 13568 14430 13632
rect 14494 13568 14510 13632
rect 14574 13568 14590 13632
rect 14654 13568 14670 13632
rect 14734 13568 14742 13632
rect 14422 12544 14742 13568
rect 14966 12885 15026 21387
rect 15147 19684 15213 19685
rect 15147 19620 15148 19684
rect 15212 19620 15213 19684
rect 15147 19619 15213 19620
rect 15150 17645 15210 19619
rect 15147 17644 15213 17645
rect 15147 17580 15148 17644
rect 15212 17580 15213 17644
rect 15147 17579 15213 17580
rect 15150 13021 15210 17579
rect 15147 13020 15213 13021
rect 15147 12956 15148 13020
rect 15212 12956 15213 13020
rect 15147 12955 15213 12956
rect 14963 12884 15029 12885
rect 14963 12820 14964 12884
rect 15028 12820 15029 12884
rect 14963 12819 15029 12820
rect 14422 12480 14430 12544
rect 14494 12480 14510 12544
rect 14574 12480 14590 12544
rect 14654 12480 14670 12544
rect 14734 12480 14742 12544
rect 14422 11456 14742 12480
rect 15334 11525 15394 26283
rect 15699 24852 15765 24853
rect 15699 24788 15700 24852
rect 15764 24788 15765 24852
rect 15699 24787 15765 24788
rect 15515 19140 15581 19141
rect 15515 19076 15516 19140
rect 15580 19076 15581 19140
rect 15515 19075 15581 19076
rect 15518 18733 15578 19075
rect 15515 18732 15581 18733
rect 15515 18668 15516 18732
rect 15580 18668 15581 18732
rect 15515 18667 15581 18668
rect 15515 16692 15581 16693
rect 15515 16628 15516 16692
rect 15580 16628 15581 16692
rect 15515 16627 15581 16628
rect 15518 13973 15578 16627
rect 15515 13972 15581 13973
rect 15515 13908 15516 13972
rect 15580 13908 15581 13972
rect 15515 13907 15581 13908
rect 15331 11524 15397 11525
rect 15331 11460 15332 11524
rect 15396 11460 15397 11524
rect 15331 11459 15397 11460
rect 14422 11392 14430 11456
rect 14494 11392 14510 11456
rect 14574 11392 14590 11456
rect 14654 11392 14670 11456
rect 14734 11392 14742 11456
rect 14422 10368 14742 11392
rect 14422 10304 14430 10368
rect 14494 10304 14510 10368
rect 14574 10304 14590 10368
rect 14654 10304 14670 10368
rect 14734 10304 14742 10368
rect 14422 9280 14742 10304
rect 14422 9216 14430 9280
rect 14494 9216 14510 9280
rect 14574 9216 14590 9280
rect 14654 9216 14670 9280
rect 14734 9216 14742 9280
rect 14422 8192 14742 9216
rect 15702 9077 15762 24787
rect 18278 21861 18338 26283
rect 18914 26144 19235 27168
rect 23407 28864 23727 28880
rect 23407 28800 23415 28864
rect 23479 28800 23495 28864
rect 23559 28800 23575 28864
rect 23639 28800 23655 28864
rect 23719 28800 23727 28864
rect 23407 27776 23727 28800
rect 23407 27712 23415 27776
rect 23479 27712 23495 27776
rect 23559 27712 23575 27776
rect 23639 27712 23655 27776
rect 23719 27712 23727 27776
rect 23407 26688 23727 27712
rect 23795 27708 23861 27709
rect 23795 27644 23796 27708
rect 23860 27644 23861 27708
rect 23795 27643 23861 27644
rect 23407 26624 23415 26688
rect 23479 26624 23495 26688
rect 23559 26624 23575 26688
rect 23639 26624 23655 26688
rect 23719 26624 23727 26688
rect 19563 26348 19629 26349
rect 19563 26284 19564 26348
rect 19628 26284 19629 26348
rect 19563 26283 19629 26284
rect 23243 26348 23309 26349
rect 23243 26284 23244 26348
rect 23308 26284 23309 26348
rect 23243 26283 23309 26284
rect 18914 26080 18922 26144
rect 18986 26080 19002 26144
rect 19066 26080 19082 26144
rect 19146 26080 19162 26144
rect 19226 26080 19235 26144
rect 18914 25056 19235 26080
rect 18914 24992 18922 25056
rect 18986 24992 19002 25056
rect 19066 24992 19082 25056
rect 19146 24992 19162 25056
rect 19226 24992 19235 25056
rect 18914 23968 19235 24992
rect 18914 23904 18922 23968
rect 18986 23904 19002 23968
rect 19066 23904 19082 23968
rect 19146 23904 19162 23968
rect 19226 23904 19235 23968
rect 18914 22880 19235 23904
rect 18914 22816 18922 22880
rect 18986 22816 19002 22880
rect 19066 22816 19082 22880
rect 19146 22816 19162 22880
rect 19226 22816 19235 22880
rect 18275 21860 18341 21861
rect 18275 21796 18276 21860
rect 18340 21796 18341 21860
rect 18275 21795 18341 21796
rect 18914 21792 19235 22816
rect 18914 21728 18922 21792
rect 18986 21728 19002 21792
rect 19066 21728 19082 21792
rect 19146 21728 19162 21792
rect 19226 21728 19235 21792
rect 18914 20704 19235 21728
rect 18914 20640 18922 20704
rect 18986 20640 19002 20704
rect 19066 20640 19082 20704
rect 19146 20640 19162 20704
rect 19226 20640 19235 20704
rect 15883 19956 15949 19957
rect 15883 19892 15884 19956
rect 15948 19892 15949 19956
rect 15883 19891 15949 19892
rect 18459 19956 18525 19957
rect 18459 19892 18460 19956
rect 18524 19892 18525 19956
rect 18459 19891 18525 19892
rect 15886 14653 15946 19891
rect 16435 19820 16501 19821
rect 16435 19756 16436 19820
rect 16500 19756 16501 19820
rect 16435 19755 16501 19756
rect 16251 19276 16317 19277
rect 16251 19212 16252 19276
rect 16316 19212 16317 19276
rect 16251 19211 16317 19212
rect 16067 18732 16133 18733
rect 16067 18668 16068 18732
rect 16132 18668 16133 18732
rect 16067 18667 16133 18668
rect 15883 14652 15949 14653
rect 15883 14588 15884 14652
rect 15948 14588 15949 14652
rect 15883 14587 15949 14588
rect 15886 11117 15946 14587
rect 16070 13837 16130 18667
rect 16254 16829 16314 19211
rect 16251 16828 16317 16829
rect 16251 16764 16252 16828
rect 16316 16764 16317 16828
rect 16251 16763 16317 16764
rect 16251 16148 16317 16149
rect 16251 16084 16252 16148
rect 16316 16084 16317 16148
rect 16251 16083 16317 16084
rect 16254 14245 16314 16083
rect 16251 14244 16317 14245
rect 16251 14180 16252 14244
rect 16316 14180 16317 14244
rect 16251 14179 16317 14180
rect 16067 13836 16133 13837
rect 16067 13772 16068 13836
rect 16132 13772 16133 13836
rect 16067 13771 16133 13772
rect 16438 12341 16498 19755
rect 16619 19276 16685 19277
rect 16619 19212 16620 19276
rect 16684 19212 16685 19276
rect 16619 19211 16685 19212
rect 16622 16421 16682 19211
rect 16803 19140 16869 19141
rect 16803 19076 16804 19140
rect 16868 19076 16869 19140
rect 16803 19075 16869 19076
rect 16806 18053 16866 19075
rect 17907 19004 17973 19005
rect 17907 18940 17908 19004
rect 17972 18940 17973 19004
rect 17907 18939 17973 18940
rect 16987 18188 17053 18189
rect 16987 18124 16988 18188
rect 17052 18124 17053 18188
rect 16987 18123 17053 18124
rect 16803 18052 16869 18053
rect 16803 17988 16804 18052
rect 16868 17988 16869 18052
rect 16803 17987 16869 17988
rect 16803 16964 16869 16965
rect 16803 16900 16804 16964
rect 16868 16900 16869 16964
rect 16803 16899 16869 16900
rect 16619 16420 16685 16421
rect 16619 16356 16620 16420
rect 16684 16356 16685 16420
rect 16619 16355 16685 16356
rect 16619 16012 16685 16013
rect 16619 15948 16620 16012
rect 16684 15948 16685 16012
rect 16619 15947 16685 15948
rect 16435 12340 16501 12341
rect 16435 12276 16436 12340
rect 16500 12276 16501 12340
rect 16435 12275 16501 12276
rect 15883 11116 15949 11117
rect 15883 11052 15884 11116
rect 15948 11052 15949 11116
rect 15883 11051 15949 11052
rect 15699 9076 15765 9077
rect 15699 9012 15700 9076
rect 15764 9012 15765 9076
rect 15699 9011 15765 9012
rect 14422 8128 14430 8192
rect 14494 8128 14510 8192
rect 14574 8128 14590 8192
rect 14654 8128 14670 8192
rect 14734 8128 14742 8192
rect 14227 7988 14293 7989
rect 14227 7924 14228 7988
rect 14292 7924 14293 7988
rect 14227 7923 14293 7924
rect 14422 7104 14742 8128
rect 14422 7040 14430 7104
rect 14494 7040 14510 7104
rect 14574 7040 14590 7104
rect 14654 7040 14670 7104
rect 14734 7040 14742 7104
rect 14422 6016 14742 7040
rect 14422 5952 14430 6016
rect 14494 5952 14510 6016
rect 14574 5952 14590 6016
rect 14654 5952 14670 6016
rect 14734 5952 14742 6016
rect 14422 4928 14742 5952
rect 14422 4864 14430 4928
rect 14494 4864 14510 4928
rect 14574 4864 14590 4928
rect 14654 4864 14670 4928
rect 14734 4864 14742 4928
rect 14422 3840 14742 4864
rect 14422 3776 14430 3840
rect 14494 3776 14510 3840
rect 14574 3776 14590 3840
rect 14654 3776 14670 3840
rect 14734 3776 14742 3840
rect 14422 2752 14742 3776
rect 16622 3501 16682 15947
rect 16806 8941 16866 16899
rect 16990 11933 17050 18123
rect 17355 17508 17421 17509
rect 17355 17444 17356 17508
rect 17420 17444 17421 17508
rect 17355 17443 17421 17444
rect 17171 17100 17237 17101
rect 17171 17036 17172 17100
rect 17236 17036 17237 17100
rect 17171 17035 17237 17036
rect 16987 11932 17053 11933
rect 16987 11868 16988 11932
rect 17052 11868 17053 11932
rect 16987 11867 17053 11868
rect 17174 10573 17234 17035
rect 17358 14925 17418 17443
rect 17355 14924 17421 14925
rect 17355 14860 17356 14924
rect 17420 14860 17421 14924
rect 17355 14859 17421 14860
rect 17358 12205 17418 14859
rect 17723 13836 17789 13837
rect 17723 13772 17724 13836
rect 17788 13772 17789 13836
rect 17723 13771 17789 13772
rect 17539 13700 17605 13701
rect 17539 13636 17540 13700
rect 17604 13636 17605 13700
rect 17539 13635 17605 13636
rect 17355 12204 17421 12205
rect 17355 12140 17356 12204
rect 17420 12140 17421 12204
rect 17355 12139 17421 12140
rect 17355 12068 17421 12069
rect 17355 12004 17356 12068
rect 17420 12004 17421 12068
rect 17355 12003 17421 12004
rect 17171 10572 17237 10573
rect 17171 10508 17172 10572
rect 17236 10508 17237 10572
rect 17171 10507 17237 10508
rect 16803 8940 16869 8941
rect 16803 8876 16804 8940
rect 16868 8876 16869 8940
rect 16803 8875 16869 8876
rect 17358 5541 17418 12003
rect 17542 11797 17602 13635
rect 17539 11796 17605 11797
rect 17539 11732 17540 11796
rect 17604 11732 17605 11796
rect 17539 11731 17605 11732
rect 17726 11661 17786 13771
rect 17910 13429 17970 18939
rect 18091 18868 18157 18869
rect 18091 18804 18092 18868
rect 18156 18804 18157 18868
rect 18091 18803 18157 18804
rect 17907 13428 17973 13429
rect 17907 13364 17908 13428
rect 17972 13364 17973 13428
rect 17907 13363 17973 13364
rect 17907 12204 17973 12205
rect 17907 12140 17908 12204
rect 17972 12140 17973 12204
rect 17907 12139 17973 12140
rect 17723 11660 17789 11661
rect 17723 11596 17724 11660
rect 17788 11596 17789 11660
rect 17723 11595 17789 11596
rect 17910 7309 17970 12139
rect 18094 11794 18154 18803
rect 18275 18460 18341 18461
rect 18275 18396 18276 18460
rect 18340 18396 18341 18460
rect 18275 18395 18341 18396
rect 18278 17101 18338 18395
rect 18275 17100 18341 17101
rect 18275 17036 18276 17100
rect 18340 17036 18341 17100
rect 18275 17035 18341 17036
rect 18462 16965 18522 19891
rect 18914 19616 19235 20640
rect 18914 19552 18922 19616
rect 18986 19552 19002 19616
rect 19066 19552 19082 19616
rect 19146 19552 19162 19616
rect 19226 19552 19235 19616
rect 18914 18528 19235 19552
rect 18914 18464 18922 18528
rect 18986 18464 19002 18528
rect 19066 18464 19082 18528
rect 19146 18464 19162 18528
rect 19226 18464 19235 18528
rect 18914 17440 19235 18464
rect 18914 17376 18922 17440
rect 18986 17376 19002 17440
rect 19066 17376 19082 17440
rect 19146 17376 19162 17440
rect 19226 17376 19235 17440
rect 18459 16964 18525 16965
rect 18459 16900 18460 16964
rect 18524 16900 18525 16964
rect 18459 16899 18525 16900
rect 18275 16828 18341 16829
rect 18275 16764 18276 16828
rect 18340 16764 18341 16828
rect 18275 16763 18341 16764
rect 18278 11933 18338 16763
rect 18914 16352 19235 17376
rect 18914 16288 18922 16352
rect 18986 16288 19002 16352
rect 19066 16288 19082 16352
rect 19146 16288 19162 16352
rect 19226 16288 19235 16352
rect 18643 16284 18709 16285
rect 18643 16220 18644 16284
rect 18708 16220 18709 16284
rect 18643 16219 18709 16220
rect 18646 14381 18706 16219
rect 18914 15264 19235 16288
rect 18914 15200 18922 15264
rect 18986 15200 19002 15264
rect 19066 15200 19082 15264
rect 19146 15200 19162 15264
rect 19226 15200 19235 15264
rect 18643 14380 18709 14381
rect 18643 14316 18644 14380
rect 18708 14316 18709 14380
rect 18643 14315 18709 14316
rect 18914 14176 19235 15200
rect 18914 14112 18922 14176
rect 18986 14112 19002 14176
rect 19066 14112 19082 14176
rect 19146 14112 19162 14176
rect 19226 14112 19235 14176
rect 18459 13156 18525 13157
rect 18459 13092 18460 13156
rect 18524 13092 18525 13156
rect 18459 13091 18525 13092
rect 18275 11932 18341 11933
rect 18275 11868 18276 11932
rect 18340 11868 18341 11932
rect 18275 11867 18341 11868
rect 18094 11734 18338 11794
rect 18091 11116 18157 11117
rect 18091 11052 18092 11116
rect 18156 11052 18157 11116
rect 18091 11051 18157 11052
rect 17907 7308 17973 7309
rect 17907 7244 17908 7308
rect 17972 7244 17973 7308
rect 17907 7243 17973 7244
rect 18094 6085 18154 11051
rect 18091 6084 18157 6085
rect 18091 6020 18092 6084
rect 18156 6020 18157 6084
rect 18091 6019 18157 6020
rect 18278 5677 18338 11734
rect 18462 11525 18522 13091
rect 18914 13088 19235 14112
rect 18914 13024 18922 13088
rect 18986 13024 19002 13088
rect 19066 13024 19082 13088
rect 19146 13024 19162 13088
rect 19226 13024 19235 13088
rect 18914 12000 19235 13024
rect 18914 11936 18922 12000
rect 18986 11936 19002 12000
rect 19066 11936 19082 12000
rect 19146 11936 19162 12000
rect 19226 11936 19235 12000
rect 18459 11524 18525 11525
rect 18459 11460 18460 11524
rect 18524 11460 18525 11524
rect 18459 11459 18525 11460
rect 18462 8941 18522 11459
rect 18914 10912 19235 11936
rect 18914 10848 18922 10912
rect 18986 10848 19002 10912
rect 19066 10848 19082 10912
rect 19146 10848 19162 10912
rect 19226 10848 19235 10912
rect 18914 9824 19235 10848
rect 18914 9760 18922 9824
rect 18986 9760 19002 9824
rect 19066 9760 19082 9824
rect 19146 9760 19162 9824
rect 19226 9760 19235 9824
rect 18643 9620 18709 9621
rect 18643 9556 18644 9620
rect 18708 9556 18709 9620
rect 18643 9555 18709 9556
rect 18459 8940 18525 8941
rect 18459 8876 18460 8940
rect 18524 8876 18525 8940
rect 18459 8875 18525 8876
rect 18275 5676 18341 5677
rect 18275 5612 18276 5676
rect 18340 5612 18341 5676
rect 18275 5611 18341 5612
rect 17355 5540 17421 5541
rect 17355 5476 17356 5540
rect 17420 5476 17421 5540
rect 17355 5475 17421 5476
rect 16619 3500 16685 3501
rect 16619 3436 16620 3500
rect 16684 3436 16685 3500
rect 16619 3435 16685 3436
rect 18646 3229 18706 9555
rect 18914 8736 19235 9760
rect 18914 8672 18922 8736
rect 18986 8672 19002 8736
rect 19066 8672 19082 8736
rect 19146 8672 19162 8736
rect 19226 8672 19235 8736
rect 18914 7648 19235 8672
rect 19566 8261 19626 26283
rect 22691 24036 22757 24037
rect 22691 23972 22692 24036
rect 22756 23972 22757 24036
rect 22691 23971 22757 23972
rect 21219 23492 21285 23493
rect 21219 23428 21220 23492
rect 21284 23428 21285 23492
rect 21219 23427 21285 23428
rect 22323 23492 22389 23493
rect 22323 23428 22324 23492
rect 22388 23428 22389 23492
rect 22323 23427 22389 23428
rect 20483 23084 20549 23085
rect 20483 23020 20484 23084
rect 20548 23020 20549 23084
rect 20483 23019 20549 23020
rect 19563 8260 19629 8261
rect 19563 8196 19564 8260
rect 19628 8196 19629 8260
rect 19563 8195 19629 8196
rect 18914 7584 18922 7648
rect 18986 7584 19002 7648
rect 19066 7584 19082 7648
rect 19146 7584 19162 7648
rect 19226 7584 19235 7648
rect 18914 6560 19235 7584
rect 19931 7444 19997 7445
rect 19931 7380 19932 7444
rect 19996 7380 19997 7444
rect 19931 7379 19997 7380
rect 18914 6496 18922 6560
rect 18986 6496 19002 6560
rect 19066 6496 19082 6560
rect 19146 6496 19162 6560
rect 19226 6496 19235 6560
rect 18914 5472 19235 6496
rect 18914 5408 18922 5472
rect 18986 5408 19002 5472
rect 19066 5408 19082 5472
rect 19146 5408 19162 5472
rect 19226 5408 19235 5472
rect 18914 4384 19235 5408
rect 18914 4320 18922 4384
rect 18986 4320 19002 4384
rect 19066 4320 19082 4384
rect 19146 4320 19162 4384
rect 19226 4320 19235 4384
rect 18914 3296 19235 4320
rect 19934 3909 19994 7379
rect 20115 6084 20181 6085
rect 20115 6020 20116 6084
rect 20180 6020 20181 6084
rect 20115 6019 20181 6020
rect 20118 4045 20178 6019
rect 20486 5405 20546 23019
rect 21035 17780 21101 17781
rect 21035 17716 21036 17780
rect 21100 17716 21101 17780
rect 21035 17715 21101 17716
rect 20667 14380 20733 14381
rect 20667 14316 20668 14380
rect 20732 14316 20733 14380
rect 20667 14315 20733 14316
rect 20670 10845 20730 14315
rect 20667 10844 20733 10845
rect 20667 10780 20668 10844
rect 20732 10780 20733 10844
rect 20667 10779 20733 10780
rect 20667 8260 20733 8261
rect 20667 8196 20668 8260
rect 20732 8196 20733 8260
rect 20667 8195 20733 8196
rect 20670 5541 20730 8195
rect 21038 5949 21098 17715
rect 21222 11933 21282 23427
rect 21955 20772 22021 20773
rect 21955 20708 21956 20772
rect 22020 20708 22021 20772
rect 21955 20707 22021 20708
rect 22139 20772 22205 20773
rect 22139 20708 22140 20772
rect 22204 20708 22205 20772
rect 22139 20707 22205 20708
rect 21771 15332 21837 15333
rect 21771 15268 21772 15332
rect 21836 15268 21837 15332
rect 21771 15267 21837 15268
rect 21403 12612 21469 12613
rect 21403 12548 21404 12612
rect 21468 12548 21469 12612
rect 21403 12547 21469 12548
rect 21406 12069 21466 12547
rect 21403 12068 21469 12069
rect 21403 12004 21404 12068
rect 21468 12004 21469 12068
rect 21403 12003 21469 12004
rect 21219 11932 21285 11933
rect 21219 11868 21220 11932
rect 21284 11868 21285 11932
rect 21219 11867 21285 11868
rect 21774 11661 21834 15267
rect 21771 11660 21837 11661
rect 21771 11596 21772 11660
rect 21836 11596 21837 11660
rect 21771 11595 21837 11596
rect 21958 11117 22018 20707
rect 21955 11116 22021 11117
rect 21955 11052 21956 11116
rect 22020 11052 22021 11116
rect 21955 11051 22021 11052
rect 22142 10573 22202 20707
rect 22139 10572 22205 10573
rect 22139 10508 22140 10572
rect 22204 10508 22205 10572
rect 22139 10507 22205 10508
rect 21955 9484 22021 9485
rect 21955 9420 21956 9484
rect 22020 9420 22021 9484
rect 21955 9419 22021 9420
rect 21035 5948 21101 5949
rect 21035 5884 21036 5948
rect 21100 5884 21101 5948
rect 21035 5883 21101 5884
rect 21958 5677 22018 9419
rect 22326 8261 22386 23427
rect 22507 22948 22573 22949
rect 22507 22884 22508 22948
rect 22572 22884 22573 22948
rect 22507 22883 22573 22884
rect 22323 8260 22389 8261
rect 22323 8196 22324 8260
rect 22388 8196 22389 8260
rect 22323 8195 22389 8196
rect 22510 5949 22570 22883
rect 22694 16693 22754 23971
rect 23246 23221 23306 26283
rect 23407 25600 23727 26624
rect 23407 25536 23415 25600
rect 23479 25536 23495 25600
rect 23559 25536 23575 25600
rect 23639 25536 23655 25600
rect 23719 25536 23727 25600
rect 23407 24512 23727 25536
rect 23407 24448 23415 24512
rect 23479 24448 23495 24512
rect 23559 24448 23575 24512
rect 23639 24448 23655 24512
rect 23719 24448 23727 24512
rect 23407 23424 23727 24448
rect 23407 23360 23415 23424
rect 23479 23360 23495 23424
rect 23559 23360 23575 23424
rect 23639 23360 23655 23424
rect 23719 23360 23727 23424
rect 23243 23220 23309 23221
rect 23243 23156 23244 23220
rect 23308 23156 23309 23220
rect 23243 23155 23309 23156
rect 23407 22336 23727 23360
rect 23407 22272 23415 22336
rect 23479 22272 23495 22336
rect 23559 22272 23575 22336
rect 23639 22272 23655 22336
rect 23719 22272 23727 22336
rect 23407 21248 23727 22272
rect 23407 21184 23415 21248
rect 23479 21184 23495 21248
rect 23559 21184 23575 21248
rect 23639 21184 23655 21248
rect 23719 21184 23727 21248
rect 23407 20160 23727 21184
rect 23407 20096 23415 20160
rect 23479 20096 23495 20160
rect 23559 20096 23575 20160
rect 23639 20096 23655 20160
rect 23719 20096 23727 20160
rect 22875 19412 22941 19413
rect 22875 19348 22876 19412
rect 22940 19348 22941 19412
rect 22875 19347 22941 19348
rect 22691 16692 22757 16693
rect 22691 16628 22692 16692
rect 22756 16628 22757 16692
rect 22691 16627 22757 16628
rect 22878 16421 22938 19347
rect 23407 19072 23727 20096
rect 23407 19008 23415 19072
rect 23479 19008 23495 19072
rect 23559 19008 23575 19072
rect 23639 19008 23655 19072
rect 23719 19008 23727 19072
rect 23407 17984 23727 19008
rect 23407 17920 23415 17984
rect 23479 17920 23495 17984
rect 23559 17920 23575 17984
rect 23639 17920 23655 17984
rect 23719 17920 23727 17984
rect 23407 16896 23727 17920
rect 23407 16832 23415 16896
rect 23479 16832 23495 16896
rect 23559 16832 23575 16896
rect 23639 16832 23655 16896
rect 23719 16832 23727 16896
rect 22875 16420 22941 16421
rect 22875 16356 22876 16420
rect 22940 16356 22941 16420
rect 22875 16355 22941 16356
rect 23407 15808 23727 16832
rect 23407 15744 23415 15808
rect 23479 15744 23495 15808
rect 23559 15744 23575 15808
rect 23639 15744 23655 15808
rect 23719 15744 23727 15808
rect 23243 15468 23309 15469
rect 23243 15404 23244 15468
rect 23308 15404 23309 15468
rect 23243 15403 23309 15404
rect 23246 13157 23306 15403
rect 23407 14720 23727 15744
rect 23407 14656 23415 14720
rect 23479 14656 23495 14720
rect 23559 14656 23575 14720
rect 23639 14656 23655 14720
rect 23719 14656 23727 14720
rect 23407 13632 23727 14656
rect 23407 13568 23415 13632
rect 23479 13568 23495 13632
rect 23559 13568 23575 13632
rect 23639 13568 23655 13632
rect 23719 13568 23727 13632
rect 23243 13156 23309 13157
rect 23243 13092 23244 13156
rect 23308 13092 23309 13156
rect 23243 13091 23309 13092
rect 22875 12748 22941 12749
rect 22875 12684 22876 12748
rect 22940 12684 22941 12748
rect 22875 12683 22941 12684
rect 22878 7989 22938 12683
rect 23407 12544 23727 13568
rect 23407 12480 23415 12544
rect 23479 12480 23495 12544
rect 23559 12480 23575 12544
rect 23639 12480 23655 12544
rect 23719 12480 23727 12544
rect 23407 11456 23727 12480
rect 23407 11392 23415 11456
rect 23479 11392 23495 11456
rect 23559 11392 23575 11456
rect 23639 11392 23655 11456
rect 23719 11392 23727 11456
rect 23407 10368 23727 11392
rect 23407 10304 23415 10368
rect 23479 10304 23495 10368
rect 23559 10304 23575 10368
rect 23639 10304 23655 10368
rect 23719 10304 23727 10368
rect 23407 9280 23727 10304
rect 23407 9216 23415 9280
rect 23479 9216 23495 9280
rect 23559 9216 23575 9280
rect 23639 9216 23655 9280
rect 23719 9216 23727 9280
rect 23407 8192 23727 9216
rect 23407 8128 23415 8192
rect 23479 8128 23495 8192
rect 23559 8128 23575 8192
rect 23639 8128 23655 8192
rect 23719 8128 23727 8192
rect 22875 7988 22941 7989
rect 22875 7924 22876 7988
rect 22940 7924 22941 7988
rect 22875 7923 22941 7924
rect 23407 7104 23727 8128
rect 23407 7040 23415 7104
rect 23479 7040 23495 7104
rect 23559 7040 23575 7104
rect 23639 7040 23655 7104
rect 23719 7040 23727 7104
rect 23407 6016 23727 7040
rect 23798 6221 23858 27643
rect 27475 25396 27541 25397
rect 27475 25332 27476 25396
rect 27540 25332 27541 25396
rect 27475 25331 27541 25332
rect 25083 25124 25149 25125
rect 25083 25060 25084 25124
rect 25148 25060 25149 25124
rect 25083 25059 25149 25060
rect 23979 23764 24045 23765
rect 23979 23700 23980 23764
rect 24044 23700 24045 23764
rect 23979 23699 24045 23700
rect 23982 9621 24042 23699
rect 24531 15060 24597 15061
rect 24531 14996 24532 15060
rect 24596 14996 24597 15060
rect 24531 14995 24597 14996
rect 24163 14516 24229 14517
rect 24163 14452 24164 14516
rect 24228 14452 24229 14516
rect 24163 14451 24229 14452
rect 24166 12477 24226 14451
rect 24163 12476 24229 12477
rect 24163 12412 24164 12476
rect 24228 12412 24229 12476
rect 24163 12411 24229 12412
rect 24534 11661 24594 14995
rect 24531 11660 24597 11661
rect 24531 11596 24532 11660
rect 24596 11596 24597 11660
rect 24531 11595 24597 11596
rect 23979 9620 24045 9621
rect 23979 9556 23980 9620
rect 24044 9556 24045 9620
rect 23979 9555 24045 9556
rect 25086 6493 25146 25059
rect 25267 24988 25333 24989
rect 25267 24924 25268 24988
rect 25332 24924 25333 24988
rect 25267 24923 25333 24924
rect 25270 7445 25330 24923
rect 25267 7444 25333 7445
rect 25267 7380 25268 7444
rect 25332 7380 25333 7444
rect 25267 7379 25333 7380
rect 27478 6493 27538 25331
rect 25083 6492 25149 6493
rect 25083 6428 25084 6492
rect 25148 6428 25149 6492
rect 25083 6427 25149 6428
rect 27475 6492 27541 6493
rect 27475 6428 27476 6492
rect 27540 6428 27541 6492
rect 27475 6427 27541 6428
rect 23795 6220 23861 6221
rect 23795 6156 23796 6220
rect 23860 6156 23861 6220
rect 23795 6155 23861 6156
rect 23407 5952 23415 6016
rect 23479 5952 23495 6016
rect 23559 5952 23575 6016
rect 23639 5952 23655 6016
rect 23719 5952 23727 6016
rect 22507 5948 22573 5949
rect 22507 5884 22508 5948
rect 22572 5884 22573 5948
rect 22507 5883 22573 5884
rect 21955 5676 22021 5677
rect 21955 5612 21956 5676
rect 22020 5612 22021 5676
rect 21955 5611 22021 5612
rect 20667 5540 20733 5541
rect 20667 5476 20668 5540
rect 20732 5476 20733 5540
rect 20667 5475 20733 5476
rect 20483 5404 20549 5405
rect 20483 5340 20484 5404
rect 20548 5340 20549 5404
rect 20483 5339 20549 5340
rect 23407 4928 23727 5952
rect 23407 4864 23415 4928
rect 23479 4864 23495 4928
rect 23559 4864 23575 4928
rect 23639 4864 23655 4928
rect 23719 4864 23727 4928
rect 20115 4044 20181 4045
rect 20115 3980 20116 4044
rect 20180 3980 20181 4044
rect 20115 3979 20181 3980
rect 19931 3908 19997 3909
rect 19931 3844 19932 3908
rect 19996 3844 19997 3908
rect 19931 3843 19997 3844
rect 18914 3232 18922 3296
rect 18986 3232 19002 3296
rect 19066 3232 19082 3296
rect 19146 3232 19162 3296
rect 19226 3232 19235 3296
rect 18643 3228 18709 3229
rect 18643 3164 18644 3228
rect 18708 3164 18709 3228
rect 18643 3163 18709 3164
rect 14422 2688 14430 2752
rect 14494 2688 14510 2752
rect 14574 2688 14590 2752
rect 14654 2688 14670 2752
rect 14734 2688 14742 2752
rect 12203 2548 12269 2549
rect 12203 2484 12204 2548
rect 12268 2484 12269 2548
rect 12203 2483 12269 2484
rect 9929 2144 9937 2208
rect 10001 2144 10017 2208
rect 10081 2144 10097 2208
rect 10161 2144 10177 2208
rect 10241 2144 10250 2208
rect 9929 2128 10250 2144
rect 14422 2128 14742 2688
rect 18914 2208 19235 3232
rect 18914 2144 18922 2208
rect 18986 2144 19002 2208
rect 19066 2144 19082 2208
rect 19146 2144 19162 2208
rect 19226 2144 19235 2208
rect 18914 2128 19235 2144
rect 23407 3840 23727 4864
rect 23407 3776 23415 3840
rect 23479 3776 23495 3840
rect 23559 3776 23575 3840
rect 23639 3776 23655 3840
rect 23719 3776 23727 3840
rect 23407 2752 23727 3776
rect 23407 2688 23415 2752
rect 23479 2688 23495 2752
rect 23559 2688 23575 2752
rect 23639 2688 23655 2752
rect 23719 2688 23727 2752
rect 23407 2128 23727 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 2484 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 3956 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform -1 0 2760 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform -1 0 4508 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 4232 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 5244 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform -1 0 2484 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1644511149
transform -1 0 2208 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1644511149
transform -1 0 3036 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1644511149
transform 1 0 11776 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1644511149
transform -1 0 3404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1644511149
transform -1 0 2668 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1644511149
transform -1 0 3036 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1644511149
transform -1 0 2116 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1644511149
transform -1 0 3404 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1644511149
transform -1 0 2392 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1644511149
transform -1 0 1748 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1644511149
transform -1 0 2852 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1644511149
transform -1 0 4140 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1644511149
transform -1 0 3220 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1644511149
transform 1 0 4232 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1644511149
transform 1 0 4600 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1644511149
transform 1 0 17112 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1644511149
transform -1 0 17020 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1644511149
transform 1 0 19688 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1644511149
transform -1 0 16560 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1644511149
transform 1 0 21160 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1644511149
transform 1 0 22080 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1644511149
transform -1 0 9936 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1644511149
transform 1 0 14812 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1644511149
transform 1 0 15456 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1644511149
transform 1 0 14444 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1644511149
transform 1 0 16928 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1644511149
transform 1 0 23552 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1644511149
transform -1 0 2760 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1644511149
transform -1 0 3128 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1644511149
transform -1 0 9568 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1644511149
transform 1 0 23276 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1644511149
transform -1 0 3496 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1644511149
transform -1 0 2208 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1644511149
transform -1 0 3036 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1644511149
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32
timestamp 1644511149
transform 1 0 4048 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38
timestamp 1644511149
transform 1 0 4600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5336 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68
timestamp 1644511149
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77
timestamp 1644511149
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1644511149
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88
timestamp 1644511149
transform 1 0 9200 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_96
timestamp 1644511149
transform 1 0 9936 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105
timestamp 1644511149
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_118
timestamp 1644511149
transform 1 0 11960 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_126
timestamp 1644511149
transform 1 0 12696 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132
timestamp 1644511149
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_149
timestamp 1644511149
transform 1 0 14812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_157
timestamp 1644511149
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1644511149
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp 1644511149
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1644511149
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1644511149
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_201
timestamp 1644511149
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1644511149
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1644511149
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_238
timestamp 1644511149
transform 1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_246
timestamp 1644511149
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257
timestamp 1644511149
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1644511149
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1644511149
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1644511149
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_20
timestamp 1644511149
transform 1 0 2944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_40
timestamp 1644511149
transform 1 0 4784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1644511149
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_73
timestamp 1644511149
transform 1 0 7820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_93
timestamp 1644511149
transform 1 0 9660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_104
timestamp 1644511149
transform 1 0 10672 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_129
timestamp 1644511149
transform 1 0 12972 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_138
timestamp 1644511149
transform 1 0 13800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1644511149
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_154
timestamp 1644511149
transform 1 0 15272 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1644511149
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_174
timestamp 1644511149
transform 1 0 17112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_183
timestamp 1644511149
transform 1 0 17940 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_192
timestamp 1644511149
transform 1 0 18768 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_200
timestamp 1644511149
transform 1 0 19504 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_208
timestamp 1644511149
transform 1 0 20240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1644511149
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_244
timestamp 1644511149
transform 1 0 23552 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_266
timestamp 1644511149
transform 1 0 25576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_275
timestamp 1644511149
transform 1 0 26404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_286
timestamp 1644511149
transform 1 0 27416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_10
timestamp 1644511149
transform 1 0 2024 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_17
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_35
timestamp 1644511149
transform 1 0 4324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_44
timestamp 1644511149
transform 1 0 5152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_60
timestamp 1644511149
transform 1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_70
timestamp 1644511149
transform 1 0 7544 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_79
timestamp 1644511149
transform 1 0 8372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_88
timestamp 1644511149
transform 1 0 9200 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_99
timestamp 1644511149
transform 1 0 10212 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_108
timestamp 1644511149
transform 1 0 11040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_119
timestamp 1644511149
transform 1 0 12052 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_128
timestamp 1644511149
transform 1 0 12880 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1644511149
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_157
timestamp 1644511149
transform 1 0 15548 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_168
timestamp 1644511149
transform 1 0 16560 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_185
timestamp 1644511149
transform 1 0 18124 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1644511149
transform 1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1644511149
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_211
timestamp 1644511149
transform 1 0 20516 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_220
timestamp 1644511149
transform 1 0 21344 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1644511149
transform 1 0 22632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_244
timestamp 1644511149
transform 1 0 23552 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_259
timestamp 1644511149
transform 1 0 24932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_266
timestamp 1644511149
transform 1 0 25576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_275
timestamp 1644511149
transform 1 0 26404 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_284
timestamp 1644511149
transform 1 0 27232 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_9
timestamp 1644511149
transform 1 0 1932 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_32
timestamp 1644511149
transform 1 0 4048 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_42
timestamp 1644511149
transform 1 0 4968 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_49
timestamp 1644511149
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_65
timestamp 1644511149
transform 1 0 7084 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_74
timestamp 1644511149
transform 1 0 7912 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_94
timestamp 1644511149
transform 1 0 9752 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1644511149
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_120
timestamp 1644511149
transform 1 0 12144 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_129
timestamp 1644511149
transform 1 0 12972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_145
timestamp 1644511149
transform 1 0 14444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_153
timestamp 1644511149
transform 1 0 15180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_157
timestamp 1644511149
transform 1 0 15548 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp 1644511149
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_173
timestamp 1644511149
transform 1 0 17020 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1644511149
transform 1 0 18308 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_197
timestamp 1644511149
transform 1 0 19228 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_205
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_212
timestamp 1644511149
transform 1 0 20608 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1644511149
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_228
timestamp 1644511149
transform 1 0 22080 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_248
timestamp 1644511149
transform 1 0 23920 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_252
timestamp 1644511149
transform 1 0 24288 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_259
timestamp 1644511149
transform 1 0 24932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_267
timestamp 1644511149
transform 1 0 25668 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_271
timestamp 1644511149
transform 1 0 26036 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1644511149
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_286
timestamp 1644511149
transform 1 0 27416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp 1644511149
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_36
timestamp 1644511149
transform 1 0 4416 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_42
timestamp 1644511149
transform 1 0 4968 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_59
timestamp 1644511149
transform 1 0 6532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_66
timestamp 1644511149
transform 1 0 7176 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_79
timestamp 1644511149
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_95
timestamp 1644511149
transform 1 0 9844 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_116
timestamp 1644511149
transform 1 0 11776 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1644511149
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_144
timestamp 1644511149
transform 1 0 14352 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_152
timestamp 1644511149
transform 1 0 15088 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_160
timestamp 1644511149
transform 1 0 15824 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_168
timestamp 1644511149
transform 1 0 16560 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_175
timestamp 1644511149
transform 1 0 17204 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_183
timestamp 1644511149
transform 1 0 17940 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_191
timestamp 1644511149
transform 1 0 18676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_213
timestamp 1644511149
transform 1 0 20700 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_243
timestamp 1644511149
transform 1 0 23460 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_271
timestamp 1644511149
transform 1 0 26036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_283
timestamp 1644511149
transform 1 0 27140 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1644511149
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_13
timestamp 1644511149
transform 1 0 2300 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_22
timestamp 1644511149
transform 1 0 3128 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_28
timestamp 1644511149
transform 1 0 3680 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_36
timestamp 1644511149
transform 1 0 4416 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1644511149
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_67
timestamp 1644511149
transform 1 0 7268 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_89
timestamp 1644511149
transform 1 0 9292 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_95
timestamp 1644511149
transform 1 0 9844 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_103
timestamp 1644511149
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_119
timestamp 1644511149
transform 1 0 12052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_128
timestamp 1644511149
transform 1 0 12880 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_139
timestamp 1644511149
transform 1 0 13892 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_160
timestamp 1644511149
transform 1 0 15824 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_186
timestamp 1644511149
transform 1 0 18216 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_199
timestamp 1644511149
transform 1 0 19412 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_204
timestamp 1644511149
transform 1 0 19872 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_213
timestamp 1644511149
transform 1 0 20700 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1644511149
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_231
timestamp 1644511149
transform 1 0 22356 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_235
timestamp 1644511149
transform 1 0 22724 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_240
timestamp 1644511149
transform 1 0 23184 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_258
timestamp 1644511149
transform 1 0 24840 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1644511149
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_286
timestamp 1644511149
transform 1 0 27416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_6
timestamp 1644511149
transform 1 0 1656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_13
timestamp 1644511149
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1644511149
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_39
timestamp 1644511149
transform 1 0 4692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_50
timestamp 1644511149
transform 1 0 5704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_58
timestamp 1644511149
transform 1 0 6440 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_78
timestamp 1644511149
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_92
timestamp 1644511149
transform 1 0 9568 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_100
timestamp 1644511149
transform 1 0 10304 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_118
timestamp 1644511149
transform 1 0 11960 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_125
timestamp 1644511149
transform 1 0 12604 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1644511149
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1644511149
transform 1 0 14812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_160
timestamp 1644511149
transform 1 0 15824 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_171
timestamp 1644511149
transform 1 0 16836 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_175
timestamp 1644511149
transform 1 0 17204 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1644511149
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_200
timestamp 1644511149
transform 1 0 19504 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_207
timestamp 1644511149
transform 1 0 20148 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_211
timestamp 1644511149
transform 1 0 20516 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_217
timestamp 1644511149
transform 1 0 21068 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_224
timestamp 1644511149
transform 1 0 21712 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_240
timestamp 1644511149
transform 1 0 23184 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp 1644511149
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_258
timestamp 1644511149
transform 1 0 24840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_266
timestamp 1644511149
transform 1 0 25576 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_286
timestamp 1644511149
transform 1 0 27416 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_20
timestamp 1644511149
transform 1 0 2944 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_31
timestamp 1644511149
transform 1 0 3956 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_48
timestamp 1644511149
transform 1 0 5520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_73
timestamp 1644511149
transform 1 0 7820 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_83
timestamp 1644511149
transform 1 0 8740 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_94
timestamp 1644511149
transform 1 0 9752 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_103
timestamp 1644511149
transform 1 0 10580 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_123
timestamp 1644511149
transform 1 0 12420 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_143
timestamp 1644511149
transform 1 0 14260 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_154
timestamp 1644511149
transform 1 0 15272 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_163
timestamp 1644511149
transform 1 0 16100 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_179
timestamp 1644511149
transform 1 0 17572 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_186
timestamp 1644511149
transform 1 0 18216 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_200
timestamp 1644511149
transform 1 0 19504 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1644511149
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_244
timestamp 1644511149
transform 1 0 23552 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_253
timestamp 1644511149
transform 1 0 24380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_286
timestamp 1644511149
transform 1 0 27416 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_14
timestamp 1644511149
transform 1 0 2392 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_20
timestamp 1644511149
transform 1 0 2944 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1644511149
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_39
timestamp 1644511149
transform 1 0 4692 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_48
timestamp 1644511149
transform 1 0 5520 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_55
timestamp 1644511149
transform 1 0 6164 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_63
timestamp 1644511149
transform 1 0 6900 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_69
timestamp 1644511149
transform 1 0 7452 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1644511149
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_95
timestamp 1644511149
transform 1 0 9844 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_117
timestamp 1644511149
transform 1 0 11868 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_128
timestamp 1644511149
transform 1 0 12880 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1644511149
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_147
timestamp 1644511149
transform 1 0 14628 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_168
timestamp 1644511149
transform 1 0 16560 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_174
timestamp 1644511149
transform 1 0 17112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1644511149
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_204
timestamp 1644511149
transform 1 0 19872 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_210
timestamp 1644511149
transform 1 0 20424 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_228
timestamp 1644511149
transform 1 0 22080 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_240
timestamp 1644511149
transform 1 0 23184 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1644511149
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_258
timestamp 1644511149
transform 1 0 24840 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_266
timestamp 1644511149
transform 1 0 25576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_286
timestamp 1644511149
transform 1 0 27416 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1644511149
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_13
timestamp 1644511149
transform 1 0 2300 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_19
timestamp 1644511149
transform 1 0 2852 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_33
timestamp 1644511149
transform 1 0 4140 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_38
timestamp 1644511149
transform 1 0 4600 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_44
timestamp 1644511149
transform 1 0 5152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1644511149
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1644511149
transform 1 0 6808 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_70
timestamp 1644511149
transform 1 0 7544 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_76
timestamp 1644511149
transform 1 0 8096 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_97
timestamp 1644511149
transform 1 0 10028 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_103
timestamp 1644511149
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_120
timestamp 1644511149
transform 1 0 12144 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_128
timestamp 1644511149
transform 1 0 12880 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_135
timestamp 1644511149
transform 1 0 13524 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_142
timestamp 1644511149
transform 1 0 14168 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_157
timestamp 1644511149
transform 1 0 15548 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1644511149
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_175
timestamp 1644511149
transform 1 0 17204 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_184
timestamp 1644511149
transform 1 0 18032 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_192
timestamp 1644511149
transform 1 0 18768 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_200
timestamp 1644511149
transform 1 0 19504 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_209
timestamp 1644511149
transform 1 0 20332 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_216
timestamp 1644511149
transform 1 0 20976 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_233
timestamp 1644511149
transform 1 0 22540 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_240
timestamp 1644511149
transform 1 0 23184 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_251
timestamp 1644511149
transform 1 0 24196 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_260
timestamp 1644511149
transform 1 0 25024 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_267
timestamp 1644511149
transform 1 0 25668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1644511149
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_286
timestamp 1644511149
transform 1 0 27416 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1644511149
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_45
timestamp 1644511149
transform 1 0 5244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_55
timestamp 1644511149
transform 1 0 6164 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_59
timestamp 1644511149
transform 1 0 6532 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_67
timestamp 1644511149
transform 1 0 7268 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp 1644511149
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_90
timestamp 1644511149
transform 1 0 9384 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_98
timestamp 1644511149
transform 1 0 10120 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_110
timestamp 1644511149
transform 1 0 11224 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_120
timestamp 1644511149
transform 1 0 12144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_128
timestamp 1644511149
transform 1 0 12880 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1644511149
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_148
timestamp 1644511149
transform 1 0 14720 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_155
timestamp 1644511149
transform 1 0 15364 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_159
timestamp 1644511149
transform 1 0 15732 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_167
timestamp 1644511149
transform 1 0 16468 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_175
timestamp 1644511149
transform 1 0 17204 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1644511149
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_202
timestamp 1644511149
transform 1 0 19688 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_206
timestamp 1644511149
transform 1 0 20056 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_223
timestamp 1644511149
transform 1 0 21620 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_231
timestamp 1644511149
transform 1 0 22356 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_248
timestamp 1644511149
transform 1 0 23920 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_270
timestamp 1644511149
transform 1 0 25944 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_274
timestamp 1644511149
transform 1 0 26312 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_281
timestamp 1644511149
transform 1 0 26956 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1644511149
transform 1 0 2116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_21
timestamp 1644511149
transform 1 0 3036 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_28
timestamp 1644511149
transform 1 0 3680 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_36
timestamp 1644511149
transform 1 0 4416 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_41
timestamp 1644511149
transform 1 0 4876 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1644511149
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_79
timestamp 1644511149
transform 1 0 8372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_86
timestamp 1644511149
transform 1 0 9016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_94
timestamp 1644511149
transform 1 0 9752 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1644511149
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_120
timestamp 1644511149
transform 1 0 12144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_124
timestamp 1644511149
transform 1 0 12512 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_132
timestamp 1644511149
transform 1 0 13248 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_139
timestamp 1644511149
transform 1 0 13892 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_148
timestamp 1644511149
transform 1 0 14720 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_154
timestamp 1644511149
transform 1 0 15272 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_162
timestamp 1644511149
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_174
timestamp 1644511149
transform 1 0 17112 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_182
timestamp 1644511149
transform 1 0 17848 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_189
timestamp 1644511149
transform 1 0 18492 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_196
timestamp 1644511149
transform 1 0 19136 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_211
timestamp 1644511149
transform 1 0 20516 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_215
timestamp 1644511149
transform 1 0 20884 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_229
timestamp 1644511149
transform 1 0 22172 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_234
timestamp 1644511149
transform 1 0 22632 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_242
timestamp 1644511149
transform 1 0 23368 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_256
timestamp 1644511149
transform 1 0 24656 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1644511149
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_285
timestamp 1644511149
transform 1 0 27324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_289
timestamp 1644511149
transform 1 0 27692 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_9
timestamp 1644511149
transform 1 0 1932 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1644511149
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_49
timestamp 1644511149
transform 1 0 5612 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_54
timestamp 1644511149
transform 1 0 6072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_68
timestamp 1644511149
transform 1 0 7360 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1644511149
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_93
timestamp 1644511149
transform 1 0 9660 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_99
timestamp 1644511149
transform 1 0 10212 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_105
timestamp 1644511149
transform 1 0 10764 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_125
timestamp 1644511149
transform 1 0 12604 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1644511149
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_164
timestamp 1644511149
transform 1 0 16192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_168
timestamp 1644511149
transform 1 0 16560 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_185
timestamp 1644511149
transform 1 0 18124 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1644511149
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_204
timestamp 1644511149
transform 1 0 19872 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_226
timestamp 1644511149
transform 1 0 21896 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_237
timestamp 1644511149
transform 1 0 22908 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1644511149
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_257
timestamp 1644511149
transform 1 0 24748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_274
timestamp 1644511149
transform 1 0 26312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_284
timestamp 1644511149
transform 1 0 27232 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_23
timestamp 1644511149
transform 1 0 3220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_29
timestamp 1644511149
transform 1 0 3772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_46
timestamp 1644511149
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1644511149
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_71
timestamp 1644511149
transform 1 0 7636 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_79
timestamp 1644511149
transform 1 0 8372 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_88
timestamp 1644511149
transform 1 0 9200 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_92
timestamp 1644511149
transform 1 0 9568 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_97
timestamp 1644511149
transform 1 0 10028 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1644511149
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_121
timestamp 1644511149
transform 1 0 12236 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_129
timestamp 1644511149
transform 1 0 12972 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_147
timestamp 1644511149
transform 1 0 14628 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_154
timestamp 1644511149
transform 1 0 15272 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_172
timestamp 1644511149
transform 1 0 16928 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_180
timestamp 1644511149
transform 1 0 17664 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_185
timestamp 1644511149
transform 1 0 18124 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_189
timestamp 1644511149
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_197
timestamp 1644511149
transform 1 0 19228 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_206
timestamp 1644511149
transform 1 0 20056 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_213
timestamp 1644511149
transform 1 0 20700 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1644511149
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_241
timestamp 1644511149
transform 1 0 23276 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_271
timestamp 1644511149
transform 1 0 26036 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_286
timestamp 1644511149
transform 1 0 27416 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_8
timestamp 1644511149
transform 1 0 1840 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1644511149
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_34
timestamp 1644511149
transform 1 0 4232 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_44
timestamp 1644511149
transform 1 0 5152 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_55
timestamp 1644511149
transform 1 0 6164 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_64
timestamp 1644511149
transform 1 0 6992 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_92
timestamp 1644511149
transform 1 0 9568 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_114
timestamp 1644511149
transform 1 0 11592 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_122
timestamp 1644511149
transform 1 0 12328 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_130
timestamp 1644511149
transform 1 0 13064 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1644511149
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_145
timestamp 1644511149
transform 1 0 14444 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_167
timestamp 1644511149
transform 1 0 16468 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_176
timestamp 1644511149
transform 1 0 17296 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_183
timestamp 1644511149
transform 1 0 17940 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_187
timestamp 1644511149
transform 1 0 18308 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1644511149
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_204
timestamp 1644511149
transform 1 0 19872 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_208
timestamp 1644511149
transform 1 0 20240 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_212
timestamp 1644511149
transform 1 0 20608 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_219
timestamp 1644511149
transform 1 0 21252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_227
timestamp 1644511149
transform 1 0 21988 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_238
timestamp 1644511149
transform 1 0 23000 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1644511149
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_257
timestamp 1644511149
transform 1 0 24748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_264
timestamp 1644511149
transform 1 0 25392 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_286
timestamp 1644511149
transform 1 0 27416 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1644511149
transform 1 0 1748 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_13
timestamp 1644511149
transform 1 0 2300 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_28
timestamp 1644511149
transform 1 0 3680 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_41
timestamp 1644511149
transform 1 0 4876 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1644511149
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_75
timestamp 1644511149
transform 1 0 8004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_84
timestamp 1644511149
transform 1 0 8832 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_92
timestamp 1644511149
transform 1 0 9568 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_99
timestamp 1644511149
transform 1 0 10212 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_107
timestamp 1644511149
transform 1 0 10948 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_121
timestamp 1644511149
transform 1 0 12236 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_129
timestamp 1644511149
transform 1 0 12972 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_133
timestamp 1644511149
transform 1 0 13340 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_150
timestamp 1644511149
transform 1 0 14904 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_162
timestamp 1644511149
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_185
timestamp 1644511149
transform 1 0 18124 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1644511149
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_219
timestamp 1644511149
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_230
timestamp 1644511149
transform 1 0 22264 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_255
timestamp 1644511149
transform 1 0 24564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_275
timestamp 1644511149
transform 1 0 26404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_284
timestamp 1644511149
transform 1 0 27232 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_22
timestamp 1644511149
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_46
timestamp 1644511149
transform 1 0 5336 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_55
timestamp 1644511149
transform 1 0 6164 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_62
timestamp 1644511149
transform 1 0 6808 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_76
timestamp 1644511149
transform 1 0 8096 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_90
timestamp 1644511149
transform 1 0 9384 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_98
timestamp 1644511149
transform 1 0 10120 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_106
timestamp 1644511149
transform 1 0 10856 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_110
timestamp 1644511149
transform 1 0 11224 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_118
timestamp 1644511149
transform 1 0 11960 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1644511149
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_148
timestamp 1644511149
transform 1 0 14720 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_156
timestamp 1644511149
transform 1 0 15456 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_164
timestamp 1644511149
transform 1 0 16192 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_172
timestamp 1644511149
transform 1 0 16928 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1644511149
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_204
timestamp 1644511149
transform 1 0 19872 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_224
timestamp 1644511149
transform 1 0 21712 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_244
timestamp 1644511149
transform 1 0 23552 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_270
timestamp 1644511149
transform 1 0 25944 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_280
timestamp 1644511149
transform 1 0 26864 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_288
timestamp 1644511149
transform 1 0 27600 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1644511149
transform 1 0 1748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_11
timestamp 1644511149
transform 1 0 2116 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_17
timestamp 1644511149
transform 1 0 2668 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_25
timestamp 1644511149
transform 1 0 3404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_36
timestamp 1644511149
transform 1 0 4416 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_42
timestamp 1644511149
transform 1 0 4968 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_50
timestamp 1644511149
transform 1 0 5704 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_62
timestamp 1644511149
transform 1 0 6808 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_70
timestamp 1644511149
transform 1 0 7544 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_88
timestamp 1644511149
transform 1 0 9200 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1644511149
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_122
timestamp 1644511149
transform 1 0 12328 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_131
timestamp 1644511149
transform 1 0 13156 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_139
timestamp 1644511149
transform 1 0 13892 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_148
timestamp 1644511149
transform 1 0 14720 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_156
timestamp 1644511149
transform 1 0 15456 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_162
timestamp 1644511149
transform 1 0 16008 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_182
timestamp 1644511149
transform 1 0 17848 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_191
timestamp 1644511149
transform 1 0 18676 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_203
timestamp 1644511149
transform 1 0 19780 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_211
timestamp 1644511149
transform 1 0 20516 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_216
timestamp 1644511149
transform 1 0 20976 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_233
timestamp 1644511149
transform 1 0 22540 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_245
timestamp 1644511149
transform 1 0 23644 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_255
timestamp 1644511149
transform 1 0 24564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_259
timestamp 1644511149
transform 1 0 24932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_276
timestamp 1644511149
transform 1 0 26496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_286
timestamp 1644511149
transform 1 0 27416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_11
timestamp 1644511149
transform 1 0 2116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_18
timestamp 1644511149
transform 1 0 2760 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1644511149
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_36
timestamp 1644511149
transform 1 0 4416 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_44
timestamp 1644511149
transform 1 0 5152 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_64
timestamp 1644511149
transform 1 0 6992 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_73
timestamp 1644511149
transform 1 0 7820 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1644511149
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_93
timestamp 1644511149
transform 1 0 9660 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_99
timestamp 1644511149
transform 1 0 10212 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_106
timestamp 1644511149
transform 1 0 10856 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_114
timestamp 1644511149
transform 1 0 11592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_131
timestamp 1644511149
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_159
timestamp 1644511149
transform 1 0 15732 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_163
timestamp 1644511149
transform 1 0 16100 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_180
timestamp 1644511149
transform 1 0 17664 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_203
timestamp 1644511149
transform 1 0 19780 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_223
timestamp 1644511149
transform 1 0 21620 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_237
timestamp 1644511149
transform 1 0 22908 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_247
timestamp 1644511149
transform 1 0 23828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_256
timestamp 1644511149
transform 1 0 24656 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_266
timestamp 1644511149
transform 1 0 25576 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_286
timestamp 1644511149
transform 1 0 27416 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_12
timestamp 1644511149
transform 1 0 2208 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_16
timestamp 1644511149
transform 1 0 2576 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_22
timestamp 1644511149
transform 1 0 3128 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_30
timestamp 1644511149
transform 1 0 3864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1644511149
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_63
timestamp 1644511149
transform 1 0 6900 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_70
timestamp 1644511149
transform 1 0 7544 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_79
timestamp 1644511149
transform 1 0 8372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_89
timestamp 1644511149
transform 1 0 9292 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_103
timestamp 1644511149
transform 1 0 10580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_117
timestamp 1644511149
transform 1 0 11868 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_124
timestamp 1644511149
transform 1 0 12512 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_145
timestamp 1644511149
transform 1 0 14444 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_153
timestamp 1644511149
transform 1 0 15180 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1644511149
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_175
timestamp 1644511149
transform 1 0 17204 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_183
timestamp 1644511149
transform 1 0 17940 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_203
timestamp 1644511149
transform 1 0 19780 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_211
timestamp 1644511149
transform 1 0 20516 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1644511149
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_228
timestamp 1644511149
transform 1 0 22080 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_241
timestamp 1644511149
transform 1 0 23276 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_269
timestamp 1644511149
transform 1 0 25852 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1644511149
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_286
timestamp 1644511149
transform 1 0 27416 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1644511149
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_39
timestamp 1644511149
transform 1 0 4692 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_48
timestamp 1644511149
transform 1 0 5520 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_56
timestamp 1644511149
transform 1 0 6256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_62
timestamp 1644511149
transform 1 0 6808 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_72
timestamp 1644511149
transform 1 0 7728 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_76
timestamp 1644511149
transform 1 0 8096 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1644511149
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_95
timestamp 1644511149
transform 1 0 9844 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_101
timestamp 1644511149
transform 1 0 10396 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_106
timestamp 1644511149
transform 1 0 10856 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_110
timestamp 1644511149
transform 1 0 11224 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_116
timestamp 1644511149
transform 1 0 11776 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_130
timestamp 1644511149
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1644511149
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_171
timestamp 1644511149
transform 1 0 16836 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_180
timestamp 1644511149
transform 1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1644511149
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_205
timestamp 1644511149
transform 1 0 19964 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_211
timestamp 1644511149
transform 1 0 20516 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_222
timestamp 1644511149
transform 1 0 21528 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_230
timestamp 1644511149
transform 1 0 22264 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_247
timestamp 1644511149
transform 1 0 23828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_266
timestamp 1644511149
transform 1 0 25576 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_286
timestamp 1644511149
transform 1 0 27416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_9
timestamp 1644511149
transform 1 0 1932 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_32
timestamp 1644511149
transform 1 0 4048 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1644511149
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_64
timestamp 1644511149
transform 1 0 6992 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_72
timestamp 1644511149
transform 1 0 7728 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_77
timestamp 1644511149
transform 1 0 8188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_90
timestamp 1644511149
transform 1 0 9384 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_98
timestamp 1644511149
transform 1 0 10120 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_106
timestamp 1644511149
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_116
timestamp 1644511149
transform 1 0 11776 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_129
timestamp 1644511149
transform 1 0 12972 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_146
timestamp 1644511149
transform 1 0 14536 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_155
timestamp 1644511149
transform 1 0 15364 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1644511149
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_185
timestamp 1644511149
transform 1 0 18124 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_197
timestamp 1644511149
transform 1 0 19228 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_201
timestamp 1644511149
transform 1 0 19596 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_207
timestamp 1644511149
transform 1 0 20148 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_211
timestamp 1644511149
transform 1 0 20516 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1644511149
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_229
timestamp 1644511149
transform 1 0 22172 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_242
timestamp 1644511149
transform 1 0 23368 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_255
timestamp 1644511149
transform 1 0 24564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_268
timestamp 1644511149
transform 1 0 25760 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_272
timestamp 1644511149
transform 1 0 26128 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1644511149
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_284
timestamp 1644511149
transform 1 0 27232 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_19
timestamp 1644511149
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_32
timestamp 1644511149
transform 1 0 4048 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_39
timestamp 1644511149
transform 1 0 4692 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_46
timestamp 1644511149
transform 1 0 5336 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_50
timestamp 1644511149
transform 1 0 5704 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_54
timestamp 1644511149
transform 1 0 6072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_74
timestamp 1644511149
transform 1 0 7912 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1644511149
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_92
timestamp 1644511149
transform 1 0 9568 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_102
timestamp 1644511149
transform 1 0 10488 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_119
timestamp 1644511149
transform 1 0 12052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_128
timestamp 1644511149
transform 1 0 12880 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_135
timestamp 1644511149
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_148
timestamp 1644511149
transform 1 0 14720 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_157
timestamp 1644511149
transform 1 0 15548 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_173
timestamp 1644511149
transform 1 0 17020 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_181
timestamp 1644511149
transform 1 0 17756 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_187
timestamp 1644511149
transform 1 0 18308 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_201
timestamp 1644511149
transform 1 0 19596 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_223
timestamp 1644511149
transform 1 0 21620 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_229
timestamp 1644511149
transform 1 0 22172 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_239
timestamp 1644511149
transform 1 0 23092 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_243
timestamp 1644511149
transform 1 0 23460 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1644511149
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_263
timestamp 1644511149
transform 1 0 25300 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_269
timestamp 1644511149
transform 1 0 25852 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_286
timestamp 1644511149
transform 1 0 27416 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_11
timestamp 1644511149
transform 1 0 2116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_18
timestamp 1644511149
transform 1 0 2760 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_38
timestamp 1644511149
transform 1 0 4600 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_47
timestamp 1644511149
transform 1 0 5428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_62
timestamp 1644511149
transform 1 0 6808 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_71
timestamp 1644511149
transform 1 0 7636 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_79
timestamp 1644511149
transform 1 0 8372 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_89
timestamp 1644511149
transform 1 0 9292 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_98
timestamp 1644511149
transform 1 0 10120 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_104
timestamp 1644511149
transform 1 0 10672 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1644511149
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_118
timestamp 1644511149
transform 1 0 11960 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_126
timestamp 1644511149
transform 1 0 12696 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_133
timestamp 1644511149
transform 1 0 13340 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_141
timestamp 1644511149
transform 1 0 14076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_147
timestamp 1644511149
transform 1 0 14628 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_154
timestamp 1644511149
transform 1 0 15272 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_163
timestamp 1644511149
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_175
timestamp 1644511149
transform 1 0 17204 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_183
timestamp 1644511149
transform 1 0 17940 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_201
timestamp 1644511149
transform 1 0 19596 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_213
timestamp 1644511149
transform 1 0 20700 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_220
timestamp 1644511149
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_231
timestamp 1644511149
transform 1 0 22356 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_244
timestamp 1644511149
transform 1 0 23552 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_250
timestamp 1644511149
transform 1 0 24104 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1644511149
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_284
timestamp 1644511149
transform 1 0 27232 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_19
timestamp 1644511149
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_36
timestamp 1644511149
transform 1 0 4416 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_45
timestamp 1644511149
transform 1 0 5244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_73
timestamp 1644511149
transform 1 0 7820 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_79
timestamp 1644511149
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_95
timestamp 1644511149
transform 1 0 9844 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_104
timestamp 1644511149
transform 1 0 10672 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_111
timestamp 1644511149
transform 1 0 11316 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_115
timestamp 1644511149
transform 1 0 11684 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_119
timestamp 1644511149
transform 1 0 12052 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_144
timestamp 1644511149
transform 1 0 14352 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_156
timestamp 1644511149
transform 1 0 15456 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_169
timestamp 1644511149
transform 1 0 16652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_186
timestamp 1644511149
transform 1 0 18216 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1644511149
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_201
timestamp 1644511149
transform 1 0 19596 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_208
timestamp 1644511149
transform 1 0 20240 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_223
timestamp 1644511149
transform 1 0 21620 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_236
timestamp 1644511149
transform 1 0 22816 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_246
timestamp 1644511149
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_263
timestamp 1644511149
transform 1 0 25300 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_269
timestamp 1644511149
transform 1 0 25852 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_286
timestamp 1644511149
transform 1 0 27416 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1644511149
transform 1 0 1748 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_11
timestamp 1644511149
transform 1 0 2116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_20
timestamp 1644511149
transform 1 0 2944 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_31
timestamp 1644511149
transform 1 0 3956 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_48
timestamp 1644511149
transform 1 0 5520 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_60
timestamp 1644511149
transform 1 0 6624 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_71
timestamp 1644511149
transform 1 0 7636 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_80
timestamp 1644511149
transform 1 0 8464 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_84
timestamp 1644511149
transform 1 0 8832 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_101
timestamp 1644511149
transform 1 0 10396 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1644511149
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_127
timestamp 1644511149
transform 1 0 12788 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_131
timestamp 1644511149
transform 1 0 13156 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_140
timestamp 1644511149
transform 1 0 13984 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1644511149
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_176
timestamp 1644511149
transform 1 0 17296 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1644511149
transform 1 0 17848 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_199
timestamp 1644511149
transform 1 0 19412 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1644511149
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_242
timestamp 1644511149
transform 1 0 23368 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_256
timestamp 1644511149
transform 1 0 24656 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_269
timestamp 1644511149
transform 1 0 25852 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1644511149
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_286
timestamp 1644511149
transform 1 0 27416 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_7
timestamp 1644511149
transform 1 0 1748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1644511149
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_36
timestamp 1644511149
transform 1 0 4416 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_43
timestamp 1644511149
transform 1 0 5060 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_50
timestamp 1644511149
transform 1 0 5704 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_59
timestamp 1644511149
transform 1 0 6532 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_63
timestamp 1644511149
transform 1 0 6900 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1644511149
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_88
timestamp 1644511149
transform 1 0 9200 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_99
timestamp 1644511149
transform 1 0 10212 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_119
timestamp 1644511149
transform 1 0 12052 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_126
timestamp 1644511149
transform 1 0 12696 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1644511149
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1644511149
transform 1 0 14812 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_161
timestamp 1644511149
transform 1 0 15916 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1644511149
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_178
timestamp 1644511149
transform 1 0 17480 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_188
timestamp 1644511149
transform 1 0 18400 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_205
timestamp 1644511149
transform 1 0 19964 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_212
timestamp 1644511149
transform 1 0 20608 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_227
timestamp 1644511149
transform 1 0 21988 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_235
timestamp 1644511149
transform 1 0 22724 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_246
timestamp 1644511149
transform 1 0 23736 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_262
timestamp 1644511149
transform 1 0 25208 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_286
timestamp 1644511149
transform 1 0 27416 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_25
timestamp 1644511149
transform 1 0 3404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_29
timestamp 1644511149
transform 1 0 3772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_33
timestamp 1644511149
transform 1 0 4140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_42
timestamp 1644511149
transform 1 0 4968 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_73
timestamp 1644511149
transform 1 0 7820 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_77
timestamp 1644511149
transform 1 0 8188 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_88
timestamp 1644511149
transform 1 0 9200 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_100
timestamp 1644511149
transform 1 0 10304 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_104
timestamp 1644511149
transform 1 0 10672 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1644511149
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_121
timestamp 1644511149
transform 1 0 12236 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_131
timestamp 1644511149
transform 1 0 13156 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_145
timestamp 1644511149
transform 1 0 14444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_155
timestamp 1644511149
transform 1 0 15364 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1644511149
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_174
timestamp 1644511149
transform 1 0 17112 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_178
timestamp 1644511149
transform 1 0 17480 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_185
timestamp 1644511149
transform 1 0 18124 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_206
timestamp 1644511149
transform 1 0 20056 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1644511149
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_234
timestamp 1644511149
transform 1 0 22632 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_247
timestamp 1644511149
transform 1 0 23828 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_257
timestamp 1644511149
transform 1 0 24748 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_265
timestamp 1644511149
transform 1 0 25484 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_285
timestamp 1644511149
transform 1 0 27324 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_289
timestamp 1644511149
transform 1 0 27692 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1644511149
transform 1 0 1748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_45
timestamp 1644511149
transform 1 0 5244 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_54
timestamp 1644511149
transform 1 0 6072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_66
timestamp 1644511149
transform 1 0 7176 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1644511149
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_107
timestamp 1644511149
transform 1 0 10948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_113
timestamp 1644511149
transform 1 0 11500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_130
timestamp 1644511149
transform 1 0 13064 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1644511149
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_157
timestamp 1644511149
transform 1 0 15548 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_166
timestamp 1644511149
transform 1 0 16376 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_174
timestamp 1644511149
transform 1 0 17112 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1644511149
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_222
timestamp 1644511149
transform 1 0 21528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_226
timestamp 1644511149
transform 1 0 21896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_243
timestamp 1644511149
transform 1 0 23460 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_269
timestamp 1644511149
transform 1 0 25852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_279
timestamp 1644511149
transform 1 0 26772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_286
timestamp 1644511149
transform 1 0 27416 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_25
timestamp 1644511149
transform 1 0 3404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_29
timestamp 1644511149
transform 1 0 3772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_33
timestamp 1644511149
transform 1 0 4140 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_42
timestamp 1644511149
transform 1 0 4968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_73
timestamp 1644511149
transform 1 0 7820 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_80
timestamp 1644511149
transform 1 0 8464 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_29_98
timestamp 1644511149
transform 1 0 10120 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1644511149
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_120
timestamp 1644511149
transform 1 0 12144 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_130
timestamp 1644511149
transform 1 0 13064 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_138
timestamp 1644511149
transform 1 0 13800 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_144
timestamp 1644511149
transform 1 0 14352 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_154
timestamp 1644511149
transform 1 0 15272 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1644511149
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_179
timestamp 1644511149
transform 1 0 17572 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_192
timestamp 1644511149
transform 1 0 18768 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_198
timestamp 1644511149
transform 1 0 19320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_205
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1644511149
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_234
timestamp 1644511149
transform 1 0 22632 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_254
timestamp 1644511149
transform 1 0 24472 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1644511149
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_284
timestamp 1644511149
transform 1 0 27232 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_8
timestamp 1644511149
transform 1 0 1840 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_12
timestamp 1644511149
transform 1 0 2208 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_17
timestamp 1644511149
transform 1 0 2668 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1644511149
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_35
timestamp 1644511149
transform 1 0 4324 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_43
timestamp 1644511149
transform 1 0 5060 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_63
timestamp 1644511149
transform 1 0 6900 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_90
timestamp 1644511149
transform 1 0 9384 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_102
timestamp 1644511149
transform 1 0 10488 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_114
timestamp 1644511149
transform 1 0 11592 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_125
timestamp 1644511149
transform 1 0 12604 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1644511149
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_151
timestamp 1644511149
transform 1 0 14996 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_162
timestamp 1644511149
transform 1 0 16008 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_166
timestamp 1644511149
transform 1 0 16376 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_190
timestamp 1644511149
transform 1 0 18584 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_213
timestamp 1644511149
transform 1 0 20700 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_220
timestamp 1644511149
transform 1 0 21344 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_235
timestamp 1644511149
transform 1 0 22724 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_273
timestamp 1644511149
transform 1 0 26220 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_281
timestamp 1644511149
transform 1 0 26956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_286
timestamp 1644511149
transform 1 0 27416 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_9
timestamp 1644511149
transform 1 0 1932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_16
timestamp 1644511149
transform 1 0 2576 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_23
timestamp 1644511149
transform 1 0 3220 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_43
timestamp 1644511149
transform 1 0 5060 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_65
timestamp 1644511149
transform 1 0 7084 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1644511149
transform 1 0 8372 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_99
timestamp 1644511149
transform 1 0 10212 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_107
timestamp 1644511149
transform 1 0 10948 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_121
timestamp 1644511149
transform 1 0 12236 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_130
timestamp 1644511149
transform 1 0 13064 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_134
timestamp 1644511149
transform 1 0 13432 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_143
timestamp 1644511149
transform 1 0 14260 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_147
timestamp 1644511149
transform 1 0 14628 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1644511149
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_172
timestamp 1644511149
transform 1 0 16928 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_176
timestamp 1644511149
transform 1 0 17296 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_186
timestamp 1644511149
transform 1 0 18216 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_192
timestamp 1644511149
transform 1 0 18768 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_202
timestamp 1644511149
transform 1 0 19688 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_210
timestamp 1644511149
transform 1 0 20424 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1644511149
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_229
timestamp 1644511149
transform 1 0 22172 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_244
timestamp 1644511149
transform 1 0 23552 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_255
timestamp 1644511149
transform 1 0 24564 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_268
timestamp 1644511149
transform 1 0 25760 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_272
timestamp 1644511149
transform 1 0 26128 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1644511149
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_286
timestamp 1644511149
transform 1 0 27416 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_9
timestamp 1644511149
transform 1 0 1932 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_16
timestamp 1644511149
transform 1 0 2576 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_20
timestamp 1644511149
transform 1 0 2944 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1644511149
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_37
timestamp 1644511149
transform 1 0 4508 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_50
timestamp 1644511149
transform 1 0 5704 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_57
timestamp 1644511149
transform 1 0 6348 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_71
timestamp 1644511149
transform 1 0 7636 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_79
timestamp 1644511149
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_93
timestamp 1644511149
transform 1 0 9660 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_99
timestamp 1644511149
transform 1 0 10212 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_116
timestamp 1644511149
transform 1 0 11776 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_120
timestamp 1644511149
transform 1 0 12144 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_126
timestamp 1644511149
transform 1 0 12696 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_134
timestamp 1644511149
transform 1 0 13432 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_148
timestamp 1644511149
transform 1 0 14720 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_152
timestamp 1644511149
transform 1 0 15088 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_161
timestamp 1644511149
transform 1 0 15916 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_181
timestamp 1644511149
transform 1 0 17756 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1644511149
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_200
timestamp 1644511149
transform 1 0 19504 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_212
timestamp 1644511149
transform 1 0 20608 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_223
timestamp 1644511149
transform 1 0 21620 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_237
timestamp 1644511149
transform 1 0 22908 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1644511149
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_266
timestamp 1644511149
transform 1 0 25576 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_286
timestamp 1644511149
transform 1 0 27416 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_8
timestamp 1644511149
transform 1 0 1840 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_12
timestamp 1644511149
transform 1 0 2208 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_17
timestamp 1644511149
transform 1 0 2668 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_28
timestamp 1644511149
transform 1 0 3680 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_32
timestamp 1644511149
transform 1 0 4048 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_36
timestamp 1644511149
transform 1 0 4416 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_49
timestamp 1644511149
transform 1 0 5612 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_64
timestamp 1644511149
transform 1 0 6992 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_70
timestamp 1644511149
transform 1 0 7544 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_89
timestamp 1644511149
transform 1 0 9292 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_97
timestamp 1644511149
transform 1 0 10028 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_103
timestamp 1644511149
transform 1 0 10580 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1644511149
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_129
timestamp 1644511149
transform 1 0 12972 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_135
timestamp 1644511149
transform 1 0 13524 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_155
timestamp 1644511149
transform 1 0 15364 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_162
timestamp 1644511149
transform 1 0 16008 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_177
timestamp 1644511149
transform 1 0 17388 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_197
timestamp 1644511149
transform 1 0 19228 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_211
timestamp 1644511149
transform 1 0 20516 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1644511149
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_232
timestamp 1644511149
transform 1 0 22448 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_241
timestamp 1644511149
transform 1 0 23276 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_254
timestamp 1644511149
transform 1 0 24472 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_262
timestamp 1644511149
transform 1 0 25208 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_270
timestamp 1644511149
transform 1 0 25944 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1644511149
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_286
timestamp 1644511149
transform 1 0 27416 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_10
timestamp 1644511149
transform 1 0 2024 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_17
timestamp 1644511149
transform 1 0 2668 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_21
timestamp 1644511149
transform 1 0 3036 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_32
timestamp 1644511149
transform 1 0 4048 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_39
timestamp 1644511149
transform 1 0 4692 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_43
timestamp 1644511149
transform 1 0 5060 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_51
timestamp 1644511149
transform 1 0 5796 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_75
timestamp 1644511149
transform 1 0 8004 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_88
timestamp 1644511149
transform 1 0 9200 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_99
timestamp 1644511149
transform 1 0 10212 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_108
timestamp 1644511149
transform 1 0 11040 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_115
timestamp 1644511149
transform 1 0 11684 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_135
timestamp 1644511149
transform 1 0 13524 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_145
timestamp 1644511149
transform 1 0 14444 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_152
timestamp 1644511149
transform 1 0 15088 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_173
timestamp 1644511149
transform 1 0 17020 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_179
timestamp 1644511149
transform 1 0 17572 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_184
timestamp 1644511149
transform 1 0 18032 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1644511149
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_208
timestamp 1644511149
transform 1 0 20240 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_219
timestamp 1644511149
transform 1 0 21252 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_226
timestamp 1644511149
transform 1 0 21896 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_236
timestamp 1644511149
transform 1 0 22816 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_247
timestamp 1644511149
transform 1 0 23828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_266
timestamp 1644511149
transform 1 0 25576 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_286
timestamp 1644511149
transform 1 0 27416 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_7
timestamp 1644511149
transform 1 0 1748 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_11
timestamp 1644511149
transform 1 0 2116 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_17
timestamp 1644511149
transform 1 0 2668 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_22
timestamp 1644511149
transform 1 0 3128 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_33
timestamp 1644511149
transform 1 0 4140 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_48
timestamp 1644511149
transform 1 0 5520 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_66
timestamp 1644511149
transform 1 0 7176 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_70
timestamp 1644511149
transform 1 0 7544 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_80
timestamp 1644511149
transform 1 0 8464 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_88
timestamp 1644511149
transform 1 0 9200 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_98
timestamp 1644511149
transform 1 0 10120 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_102
timestamp 1644511149
transform 1 0 10488 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1644511149
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_120
timestamp 1644511149
transform 1 0 12144 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_128
timestamp 1644511149
transform 1 0 12880 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_146
timestamp 1644511149
transform 1 0 14536 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_153
timestamp 1644511149
transform 1 0 15180 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1644511149
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_177
timestamp 1644511149
transform 1 0 17388 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_188
timestamp 1644511149
transform 1 0 18400 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_196
timestamp 1644511149
transform 1 0 19136 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_206
timestamp 1644511149
transform 1 0 20056 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1644511149
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_233
timestamp 1644511149
transform 1 0 22540 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_248
timestamp 1644511149
transform 1 0 23920 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_256
timestamp 1644511149
transform 1 0 24656 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_260
timestamp 1644511149
transform 1 0 25024 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_268
timestamp 1644511149
transform 1 0 25760 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1644511149
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_284
timestamp 1644511149
transform 1 0 27232 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_10
timestamp 1644511149
transform 1 0 2024 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_17
timestamp 1644511149
transform 1 0 2668 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_21
timestamp 1644511149
transform 1 0 3036 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_39
timestamp 1644511149
transform 1 0 4692 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_50
timestamp 1644511149
transform 1 0 5704 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_58
timestamp 1644511149
transform 1 0 6440 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_68
timestamp 1644511149
transform 1 0 7360 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1644511149
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_89
timestamp 1644511149
transform 1 0 9292 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_102
timestamp 1644511149
transform 1 0 10488 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_110
timestamp 1644511149
transform 1 0 11224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_122
timestamp 1644511149
transform 1 0 12328 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_129
timestamp 1644511149
transform 1 0 12972 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1644511149
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_145
timestamp 1644511149
transform 1 0 14444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_161
timestamp 1644511149
transform 1 0 15916 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_169
timestamp 1644511149
transform 1 0 16652 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_186
timestamp 1644511149
transform 1 0 18216 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1644511149
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_200
timestamp 1644511149
transform 1 0 19504 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_214
timestamp 1644511149
transform 1 0 20792 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_222
timestamp 1644511149
transform 1 0 21528 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_233
timestamp 1644511149
transform 1 0 22540 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1644511149
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_263
timestamp 1644511149
transform 1 0 25300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_274
timestamp 1644511149
transform 1 0 26312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_283
timestamp 1644511149
transform 1 0 27140 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_10
timestamp 1644511149
transform 1 0 2024 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_14
timestamp 1644511149
transform 1 0 2392 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_21
timestamp 1644511149
transform 1 0 3036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_28
timestamp 1644511149
transform 1 0 3680 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_37
timestamp 1644511149
transform 1 0 4508 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_48
timestamp 1644511149
transform 1 0 5520 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_61
timestamp 1644511149
transform 1 0 6716 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_68
timestamp 1644511149
transform 1 0 7360 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_75
timestamp 1644511149
transform 1 0 8004 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_88
timestamp 1644511149
transform 1 0 9200 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_99
timestamp 1644511149
transform 1 0 10212 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_106
timestamp 1644511149
transform 1 0 10856 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_117
timestamp 1644511149
transform 1 0 11868 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_135
timestamp 1644511149
transform 1 0 13524 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_139
timestamp 1644511149
transform 1 0 13892 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_145
timestamp 1644511149
transform 1 0 14444 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_155
timestamp 1644511149
transform 1 0 15364 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1644511149
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_176
timestamp 1644511149
transform 1 0 17296 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_184
timestamp 1644511149
transform 1 0 18032 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_188
timestamp 1644511149
transform 1 0 18400 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_197
timestamp 1644511149
transform 1 0 19228 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_206
timestamp 1644511149
transform 1 0 20056 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1644511149
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_239
timestamp 1644511149
transform 1 0 23092 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_37_255
timestamp 1644511149
transform 1 0 24564 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_270
timestamp 1644511149
transform 1 0 25944 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1644511149
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_286
timestamp 1644511149
transform 1 0 27416 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_7
timestamp 1644511149
transform 1 0 1748 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_11
timestamp 1644511149
transform 1 0 2116 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1644511149
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_38
timestamp 1644511149
transform 1 0 4600 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_46
timestamp 1644511149
transform 1 0 5336 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_54
timestamp 1644511149
transform 1 0 6072 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_60
timestamp 1644511149
transform 1 0 6624 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_64
timestamp 1644511149
transform 1 0 6992 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_68
timestamp 1644511149
transform 1 0 7360 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_94
timestamp 1644511149
transform 1 0 9752 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_102
timestamp 1644511149
transform 1 0 10488 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_116
timestamp 1644511149
transform 1 0 11776 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_127
timestamp 1644511149
transform 1 0 12788 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1644511149
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_148
timestamp 1644511149
transform 1 0 14720 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_152
timestamp 1644511149
transform 1 0 15088 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_159
timestamp 1644511149
transform 1 0 15732 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_180
timestamp 1644511149
transform 1 0 17664 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_186
timestamp 1644511149
transform 1 0 18216 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_190
timestamp 1644511149
transform 1 0 18584 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_203
timestamp 1644511149
transform 1 0 19780 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_211
timestamp 1644511149
transform 1 0 20516 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_219
timestamp 1644511149
transform 1 0 21252 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_226
timestamp 1644511149
transform 1 0 21896 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_236
timestamp 1644511149
transform 1 0 22816 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_246
timestamp 1644511149
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_262
timestamp 1644511149
transform 1 0 25208 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_286
timestamp 1644511149
transform 1 0 27416 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_7
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_12
timestamp 1644511149
transform 1 0 2208 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_19
timestamp 1644511149
transform 1 0 2852 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_30
timestamp 1644511149
transform 1 0 3864 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_38
timestamp 1644511149
transform 1 0 4600 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_46
timestamp 1644511149
transform 1 0 5336 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1644511149
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_66
timestamp 1644511149
transform 1 0 7176 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_78
timestamp 1644511149
transform 1 0 8280 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_88
timestamp 1644511149
transform 1 0 9200 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_101
timestamp 1644511149
transform 1 0 10396 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1644511149
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_117
timestamp 1644511149
transform 1 0 11868 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_151
timestamp 1644511149
transform 1 0 14996 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_155
timestamp 1644511149
transform 1 0 15364 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_195
timestamp 1644511149
transform 1 0 19044 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_199
timestamp 1644511149
transform 1 0 19412 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_204
timestamp 1644511149
transform 1 0 19872 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_218
timestamp 1644511149
transform 1 0 21160 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_231
timestamp 1644511149
transform 1 0 22356 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_241
timestamp 1644511149
transform 1 0 23276 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_245
timestamp 1644511149
transform 1 0 23644 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_256
timestamp 1644511149
transform 1 0 24656 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_269
timestamp 1644511149
transform 1 0 25852 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_286
timestamp 1644511149
transform 1 0 27416 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_19
timestamp 1644511149
transform 1 0 2852 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_35
timestamp 1644511149
transform 1 0 4324 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_48
timestamp 1644511149
transform 1 0 5520 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_61
timestamp 1644511149
transform 1 0 6716 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_69
timestamp 1644511149
transform 1 0 7452 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_78
timestamp 1644511149
transform 1 0 8280 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_88
timestamp 1644511149
transform 1 0 9200 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_94
timestamp 1644511149
transform 1 0 9752 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_102
timestamp 1644511149
transform 1 0 10488 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_116
timestamp 1644511149
transform 1 0 11776 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_122
timestamp 1644511149
transform 1 0 12328 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_127
timestamp 1644511149
transform 1 0 12788 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_134
timestamp 1644511149
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_151
timestamp 1644511149
transform 1 0 14996 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_159
timestamp 1644511149
transform 1 0 15732 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_166
timestamp 1644511149
transform 1 0 16376 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_178
timestamp 1644511149
transform 1 0 17480 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1644511149
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_206
timestamp 1644511149
transform 1 0 20056 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_213
timestamp 1644511149
transform 1 0 20700 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_226
timestamp 1644511149
transform 1 0 21896 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_237
timestamp 1644511149
transform 1 0 22908 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1644511149
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_256
timestamp 1644511149
transform 1 0 24656 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_260
timestamp 1644511149
transform 1 0 25024 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_266
timestamp 1644511149
transform 1 0 25576 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_286
timestamp 1644511149
transform 1 0 27416 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_8
timestamp 1644511149
transform 1 0 1840 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_19
timestamp 1644511149
transform 1 0 2852 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_30
timestamp 1644511149
transform 1 0 3864 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_41
timestamp 1644511149
transform 1 0 4876 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_47
timestamp 1644511149
transform 1 0 5428 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_52
timestamp 1644511149
transform 1 0 5888 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_63
timestamp 1644511149
transform 1 0 6900 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_73
timestamp 1644511149
transform 1 0 7820 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_85
timestamp 1644511149
transform 1 0 8924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_94
timestamp 1644511149
transform 1 0 9752 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_101
timestamp 1644511149
transform 1 0 10396 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1644511149
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_116
timestamp 1644511149
transform 1 0 11776 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_123
timestamp 1644511149
transform 1 0 12420 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_132
timestamp 1644511149
transform 1 0 13248 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_139
timestamp 1644511149
transform 1 0 13892 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_147
timestamp 1644511149
transform 1 0 14628 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_158
timestamp 1644511149
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1644511149
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_172
timestamp 1644511149
transform 1 0 16928 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_176
timestamp 1644511149
transform 1 0 17296 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_187
timestamp 1644511149
transform 1 0 18308 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_200
timestamp 1644511149
transform 1 0 19504 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_213
timestamp 1644511149
transform 1 0 20700 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1644511149
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_236
timestamp 1644511149
transform 1 0 22816 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_240
timestamp 1644511149
transform 1 0 23184 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_251
timestamp 1644511149
transform 1 0 24196 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_262
timestamp 1644511149
transform 1 0 25208 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_269
timestamp 1644511149
transform 1 0 25852 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1644511149
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_286
timestamp 1644511149
transform 1 0 27416 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_10
timestamp 1644511149
transform 1 0 2024 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_17
timestamp 1644511149
transform 1 0 2668 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_24
timestamp 1644511149
transform 1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_36
timestamp 1644511149
transform 1 0 4416 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_54
timestamp 1644511149
transform 1 0 6072 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_60
timestamp 1644511149
transform 1 0 6624 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_75
timestamp 1644511149
transform 1 0 8004 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_89
timestamp 1644511149
transform 1 0 9292 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_96
timestamp 1644511149
transform 1 0 9936 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_116
timestamp 1644511149
transform 1 0 11776 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_122
timestamp 1644511149
transform 1 0 12328 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_130
timestamp 1644511149
transform 1 0 13064 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1644511149
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_147
timestamp 1644511149
transform 1 0 14628 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_162
timestamp 1644511149
transform 1 0 16008 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_166
timestamp 1644511149
transform 1 0 16376 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_173
timestamp 1644511149
transform 1 0 17020 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_181
timestamp 1644511149
transform 1 0 17756 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1644511149
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_201
timestamp 1644511149
transform 1 0 19596 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1644511149
transform 1 0 20516 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_217
timestamp 1644511149
transform 1 0 21068 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_232
timestamp 1644511149
transform 1 0 22448 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_260
timestamp 1644511149
transform 1 0 25024 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_280
timestamp 1644511149
transform 1 0 26864 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_288
timestamp 1644511149
transform 1 0 27600 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_7
timestamp 1644511149
transform 1 0 1748 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_24
timestamp 1644511149
transform 1 0 3312 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_30
timestamp 1644511149
transform 1 0 3864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_40
timestamp 1644511149
transform 1 0 4784 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_50
timestamp 1644511149
transform 1 0 5704 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_64
timestamp 1644511149
transform 1 0 6992 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_72
timestamp 1644511149
transform 1 0 7728 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_78
timestamp 1644511149
transform 1 0 8280 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_88
timestamp 1644511149
transform 1 0 9200 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_97
timestamp 1644511149
transform 1 0 10028 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_117
timestamp 1644511149
transform 1 0 11868 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_133
timestamp 1644511149
transform 1 0 13340 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_142
timestamp 1644511149
transform 1 0 14168 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_155
timestamp 1644511149
transform 1 0 15364 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_163
timestamp 1644511149
transform 1 0 16100 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_172
timestamp 1644511149
transform 1 0 16928 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_176
timestamp 1644511149
transform 1 0 17296 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_186
timestamp 1644511149
transform 1 0 18216 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_195
timestamp 1644511149
transform 1 0 19044 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_206
timestamp 1644511149
transform 1 0 20056 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_213
timestamp 1644511149
transform 1 0 20700 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1644511149
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_232
timestamp 1644511149
transform 1 0 22448 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_247
timestamp 1644511149
transform 1 0 23828 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_256
timestamp 1644511149
transform 1 0 24656 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_265
timestamp 1644511149
transform 1 0 25484 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_271
timestamp 1644511149
transform 1 0 26036 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_275
timestamp 1644511149
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_284
timestamp 1644511149
transform 1 0 27232 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_7
timestamp 1644511149
transform 1 0 1748 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_11
timestamp 1644511149
transform 1 0 2116 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1644511149
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_44
timestamp 1644511149
transform 1 0 5152 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_49
timestamp 1644511149
transform 1 0 5612 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_56
timestamp 1644511149
transform 1 0 6256 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_64
timestamp 1644511149
transform 1 0 6992 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_75
timestamp 1644511149
transform 1 0 8004 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_92
timestamp 1644511149
transform 1 0 9568 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_104
timestamp 1644511149
transform 1 0 10672 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_115
timestamp 1644511149
transform 1 0 11684 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_123
timestamp 1644511149
transform 1 0 12420 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_135
timestamp 1644511149
transform 1 0 13524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_148
timestamp 1644511149
transform 1 0 14720 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_161
timestamp 1644511149
transform 1 0 15916 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_170
timestamp 1644511149
transform 1 0 16744 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_178
timestamp 1644511149
transform 1 0 17480 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_186
timestamp 1644511149
transform 1 0 18216 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1644511149
transform 1 0 18952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_204
timestamp 1644511149
transform 1 0 19872 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_213
timestamp 1644511149
transform 1 0 20700 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_222
timestamp 1644511149
transform 1 0 21528 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_242
timestamp 1644511149
transform 1 0 23368 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1644511149
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_269
timestamp 1644511149
transform 1 0 25852 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_276
timestamp 1644511149
transform 1 0 26496 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_283
timestamp 1644511149
transform 1 0 27140 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_6
timestamp 1644511149
transform 1 0 1656 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_10
timestamp 1644511149
transform 1 0 2024 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_14
timestamp 1644511149
transform 1 0 2392 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_18
timestamp 1644511149
transform 1 0 2760 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_22
timestamp 1644511149
transform 1 0 3128 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_26
timestamp 1644511149
transform 1 0 3496 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1644511149
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_65
timestamp 1644511149
transform 1 0 7084 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_73
timestamp 1644511149
transform 1 0 7820 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_84
timestamp 1644511149
transform 1 0 8832 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_97
timestamp 1644511149
transform 1 0 10028 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1644511149
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_118
timestamp 1644511149
transform 1 0 11960 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_131
timestamp 1644511149
transform 1 0 13156 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_141
timestamp 1644511149
transform 1 0 14076 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_185
timestamp 1644511149
transform 1 0 18124 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_196
timestamp 1644511149
transform 1 0 19136 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1644511149
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_228
timestamp 1644511149
transform 1 0 22080 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_235
timestamp 1644511149
transform 1 0 22724 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_242
timestamp 1644511149
transform 1 0 23368 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_256
timestamp 1644511149
transform 1 0 24656 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_264
timestamp 1644511149
transform 1 0 25392 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_269
timestamp 1644511149
transform 1 0 25852 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1644511149
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_286
timestamp 1644511149
transform 1 0 27416 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_10
timestamp 1644511149
transform 1 0 2024 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_17
timestamp 1644511149
transform 1 0 2668 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp 1644511149
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_33
timestamp 1644511149
transform 1 0 4140 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_40
timestamp 1644511149
transform 1 0 4784 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_44
timestamp 1644511149
transform 1 0 5152 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_47
timestamp 1644511149
transform 1 0 5428 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_52
timestamp 1644511149
transform 1 0 5888 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_74
timestamp 1644511149
transform 1 0 7912 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1644511149
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_101
timestamp 1644511149
transform 1 0 10396 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_107
timestamp 1644511149
transform 1 0 10948 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_124
timestamp 1644511149
transform 1 0 12512 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_151
timestamp 1644511149
transform 1 0 14996 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_156
timestamp 1644511149
transform 1 0 15456 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_164
timestamp 1644511149
transform 1 0 16192 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_168
timestamp 1644511149
transform 1 0 16560 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_173
timestamp 1644511149
transform 1 0 17020 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_178
timestamp 1644511149
transform 1 0 17480 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_186
timestamp 1644511149
transform 1 0 18216 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1644511149
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_213
timestamp 1644511149
transform 1 0 20700 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_219
timestamp 1644511149
transform 1 0 21252 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_244
timestamp 1644511149
transform 1 0 23552 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1644511149
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_256
timestamp 1644511149
transform 1 0 24656 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_263
timestamp 1644511149
transform 1 0 25300 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_267
timestamp 1644511149
transform 1 0 25668 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_271
timestamp 1644511149
transform 1 0 26036 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_278
timestamp 1644511149
transform 1 0 26680 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_286
timestamp 1644511149
transform 1 0 27416 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_18
timestamp 1644511149
transform 1 0 2760 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_23
timestamp 1644511149
transform 1 0 3220 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_31
timestamp 1644511149
transform 1 0 3956 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_52
timestamp 1644511149
transform 1 0 5888 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_65
timestamp 1644511149
transform 1 0 7084 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_82
timestamp 1644511149
transform 1 0 8648 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_90
timestamp 1644511149
transform 1 0 9384 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1644511149
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_134
timestamp 1644511149
transform 1 0 13432 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_142
timestamp 1644511149
transform 1 0 14168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_159
timestamp 1644511149
transform 1 0 15732 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_185
timestamp 1644511149
transform 1 0 18124 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_212
timestamp 1644511149
transform 1 0 20608 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_219
timestamp 1644511149
transform 1 0 21252 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_234
timestamp 1644511149
transform 1 0 22632 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_240
timestamp 1644511149
transform 1 0 23184 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_243
timestamp 1644511149
transform 1 0 23460 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_248
timestamp 1644511149
transform 1 0 23920 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_260
timestamp 1644511149
transform 1 0 25024 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_272
timestamp 1644511149
transform 1 0 26128 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1644511149
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_284
timestamp 1644511149
transform 1 0 27232 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_57
timestamp 1644511149
transform 1 0 6348 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_69
timestamp 1644511149
transform 1 0 7452 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_75
timestamp 1644511149
transform 1 0 8004 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_89
timestamp 1644511149
transform 1 0 9292 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_92
timestamp 1644511149
transform 1 0 9568 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_96
timestamp 1644511149
transform 1 0 9936 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_101
timestamp 1644511149
transform 1 0 10396 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_108
timestamp 1644511149
transform 1 0 11040 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_113
timestamp 1644511149
transform 1 0 11500 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_118
timestamp 1644511149
transform 1 0 11960 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_123
timestamp 1644511149
transform 1 0 12420 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_132
timestamp 1644511149
transform 1 0 13248 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_147
timestamp 1644511149
transform 1 0 14628 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_152
timestamp 1644511149
transform 1 0 15088 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_158
timestamp 1644511149
transform 1 0 15640 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_163
timestamp 1644511149
transform 1 0 16100 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_169
timestamp 1644511149
transform 1 0 16652 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_174
timestamp 1644511149
transform 1 0 17112 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_179
timestamp 1644511149
transform 1 0 17572 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_186
timestamp 1644511149
transform 1 0 18216 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_190
timestamp 1644511149
transform 1 0 18584 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_201
timestamp 1644511149
transform 1 0 19596 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_204
timestamp 1644511149
transform 1 0 19872 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_216
timestamp 1644511149
transform 1 0 20976 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_220
timestamp 1644511149
transform 1 0 21344 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_225
timestamp 1644511149
transform 1 0 21804 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_230
timestamp 1644511149
transform 1 0 22264 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_235
timestamp 1644511149
transform 1 0 22724 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_242
timestamp 1644511149
transform 1 0 23368 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_246
timestamp 1644511149
transform 1 0 23736 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_281
timestamp 1644511149
transform 1 0 26956 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_286
timestamp 1644511149
transform 1 0 27416 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 28060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 28060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 28060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 28060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 28060 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 28060 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 28060 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 28060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 28060 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 28060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 28060 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 28060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 28060 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 28060 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 28060 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 28060 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 28060 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 28060 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 28060 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 28060 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 28060 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 28060 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 28060 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 28060 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 28060 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 28060 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 28060 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 28060 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 28060 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 28060 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 28060 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 28060 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 28060 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 28060 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 28060 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 28060 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 28060 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 28060 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 28060 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 28060 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 28060 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 28060 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 28060 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 28060 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 28060 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 28060 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 28060 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 28060 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 28060 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 6256 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 11408 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 16560 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 21712 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 26864 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0787_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11040 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _0788_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5060 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0789_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6440 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0790_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4600 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0791_
timestamp 1644511149
transform 1 0 5612 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0792_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5244 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0793_
timestamp 1644511149
transform 1 0 9292 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0794_
timestamp 1644511149
transform 1 0 4416 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0795_
timestamp 1644511149
transform 1 0 6992 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0796_
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _0797_
timestamp 1644511149
transform 1 0 7728 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0798_
timestamp 1644511149
transform 1 0 8740 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2b_2  _0799_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11316 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0800_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9936 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0801_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9752 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _0802_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12420 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1644511149
transform 1 0 14996 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0804_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0805_
timestamp 1644511149
transform 1 0 14260 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0806_
timestamp 1644511149
transform 1 0 12420 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1644511149
transform 1 0 10120 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0808_
timestamp 1644511149
transform 1 0 4784 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0809_
timestamp 1644511149
transform 1 0 8188 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1644511149
transform 1 0 6072 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1644511149
transform 1 0 4140 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0812_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7452 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0813_
timestamp 1644511149
transform 1 0 6716 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0814_
timestamp 1644511149
transform 1 0 7268 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__nand3b_2  _0815_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4784 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _0816_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4048 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0817_
timestamp 1644511149
transform 1 0 5428 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_2  _0818_
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0819_
timestamp 1644511149
transform 1 0 6716 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_2  _0820_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5152 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0821_
timestamp 1644511149
transform 1 0 4876 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0822_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3496 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _0823_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5060 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0824_
timestamp 1644511149
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0825_
timestamp 1644511149
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0826_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0827_
timestamp 1644511149
transform 1 0 7912 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0828_
timestamp 1644511149
transform 1 0 8004 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _0829_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0830_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7084 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0831_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6624 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0832_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6532 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0833_
timestamp 1644511149
transform 1 0 10856 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _0834_
timestamp 1644511149
transform 1 0 9568 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0835_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10580 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0836_
timestamp 1644511149
transform 1 0 9568 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0837_
timestamp 1644511149
transform 1 0 8648 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0838_
timestamp 1644511149
transform 1 0 7636 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__a2111o_1  _0839_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7636 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0840_
timestamp 1644511149
transform 1 0 7912 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0841_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4048 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0842_
timestamp 1644511149
transform 1 0 4876 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0843_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0844_
timestamp 1644511149
transform 1 0 10120 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _0845_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9660 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_2  _0846_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9384 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_1  _0847_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10580 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0848_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0849_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14168 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0850_
timestamp 1644511149
transform 1 0 14812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _0851_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11592 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0852_
timestamp 1644511149
transform 1 0 11960 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0853_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12972 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0854_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27140 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1644511149
transform 1 0 13616 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0856_
timestamp 1644511149
transform 1 0 14904 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0857_
timestamp 1644511149
transform 1 0 15548 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0858_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15732 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0859_
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0860_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0861_
timestamp 1644511149
transform 1 0 21620 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _0862_
timestamp 1644511149
transform 1 0 14996 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0863_
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0864_
timestamp 1644511149
transform 1 0 18400 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0865_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22264 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _0866_
timestamp 1644511149
transform 1 0 18768 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0867_
timestamp 1644511149
transform 1 0 22448 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0868_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17572 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0869_
timestamp 1644511149
transform 1 0 20424 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0870_
timestamp 1644511149
transform 1 0 21896 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0871_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13984 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0872_
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0873_
timestamp 1644511149
transform 1 0 15364 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0874_
timestamp 1644511149
transform 1 0 16468 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0875_
timestamp 1644511149
transform 1 0 15824 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0876_
timestamp 1644511149
transform 1 0 17204 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0877_
timestamp 1644511149
transform 1 0 22172 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0878_
timestamp 1644511149
transform 1 0 22724 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0879_
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0880_
timestamp 1644511149
transform 1 0 19872 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0881_
timestamp 1644511149
transform 1 0 18124 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0882_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21160 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0883_
timestamp 1644511149
transform 1 0 22264 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _0884_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16468 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _0885_
timestamp 1644511149
transform 1 0 19504 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0886_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22172 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0887_
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0888_
timestamp 1644511149
transform 1 0 20792 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0889_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0890_
timestamp 1644511149
transform 1 0 18308 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0891_
timestamp 1644511149
transform 1 0 20516 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0892_
timestamp 1644511149
transform 1 0 19228 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0893_
timestamp 1644511149
transform 1 0 20884 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0894_
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0895_
timestamp 1644511149
transform 1 0 19596 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0896_
timestamp 1644511149
transform 1 0 19872 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _0897_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16744 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0898_
timestamp 1644511149
transform 1 0 20240 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _0899_
timestamp 1644511149
transform 1 0 20608 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0900_
timestamp 1644511149
transform 1 0 22816 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0901_
timestamp 1644511149
transform 1 0 27140 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0903_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11960 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0905_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7176 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0906_
timestamp 1644511149
transform 1 0 7912 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0907_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10304 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0908_
timestamp 1644511149
transform 1 0 9752 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0909_
timestamp 1644511149
transform 1 0 9752 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0911_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9844 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0912_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12696 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0913_
timestamp 1644511149
transform 1 0 15640 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0914_
timestamp 1644511149
transform 1 0 15916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0915_
timestamp 1644511149
transform 1 0 12144 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0916_
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0917_
timestamp 1644511149
transform 1 0 11868 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0918_
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0919_
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0920_
timestamp 1644511149
transform 1 0 11776 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0921_
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0922_
timestamp 1644511149
transform 1 0 14076 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _0923_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13248 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0924_
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0925_
timestamp 1644511149
transform 1 0 13340 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0926_
timestamp 1644511149
transform 1 0 14168 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0927_
timestamp 1644511149
transform 1 0 13064 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0928_
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0929_
timestamp 1644511149
transform 1 0 12880 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0930_
timestamp 1644511149
transform 1 0 12788 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0931_
timestamp 1644511149
transform 1 0 10764 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0932_
timestamp 1644511149
transform 1 0 14260 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0933_
timestamp 1644511149
transform 1 0 11316 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0934_
timestamp 1644511149
transform 1 0 20608 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0935_
timestamp 1644511149
transform 1 0 13248 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0936_
timestamp 1644511149
transform 1 0 15824 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0937_
timestamp 1644511149
transform 1 0 16928 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0938_
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0939_
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0940_
timestamp 1644511149
transform 1 0 21988 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0941_
timestamp 1644511149
transform 1 0 12420 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0942_
timestamp 1644511149
transform 1 0 12420 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0943_
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0944_
timestamp 1644511149
transform 1 0 15640 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0945_
timestamp 1644511149
transform 1 0 11500 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0946_
timestamp 1644511149
transform 1 0 14168 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0947_
timestamp 1644511149
transform 1 0 15548 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0948_
timestamp 1644511149
transform 1 0 14352 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0949_
timestamp 1644511149
transform 1 0 14352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0950_
timestamp 1644511149
transform 1 0 18584 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0951_
timestamp 1644511149
transform 1 0 12144 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0952_
timestamp 1644511149
transform 1 0 20608 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0953_
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0954_
timestamp 1644511149
transform 1 0 20332 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0955_
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0956_
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0957_
timestamp 1644511149
transform 1 0 14720 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0958_
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0959_
timestamp 1644511149
transform 1 0 16100 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0960_
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0961_
timestamp 1644511149
transform 1 0 15732 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0962_
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0963_
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0964_
timestamp 1644511149
transform 1 0 16928 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0965_
timestamp 1644511149
transform 1 0 17940 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0966_
timestamp 1644511149
transform 1 0 23276 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0967_
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_2  _0968_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23000 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0969_
timestamp 1644511149
transform 1 0 18584 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0970_
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0971_
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0972_
timestamp 1644511149
transform 1 0 20700 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0973_
timestamp 1644511149
transform 1 0 17480 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0974_
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_4  _0975_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__and2b_1  _0976_
timestamp 1644511149
transform 1 0 18676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0977_
timestamp 1644511149
transform 1 0 19228 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0978_
timestamp 1644511149
transform 1 0 15640 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0979_
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0980_
timestamp 1644511149
transform 1 0 18308 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0981_
timestamp 1644511149
transform 1 0 19872 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_4  _0982_
timestamp 1644511149
transform 1 0 23000 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_1  _0983_
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0984_
timestamp 1644511149
transform 1 0 19688 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0985_
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0986_
timestamp 1644511149
transform 1 0 21896 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0987_
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0988_
timestamp 1644511149
transform 1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0989_
timestamp 1644511149
transform 1 0 12880 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0990_
timestamp 1644511149
transform 1 0 18032 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0991_
timestamp 1644511149
transform 1 0 18216 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 1644511149
transform 1 0 20700 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0993_
timestamp 1644511149
transform 1 0 15088 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0994_
timestamp 1644511149
transform 1 0 18492 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0995_
timestamp 1644511149
transform 1 0 20056 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1644511149
transform 1 0 22908 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0997_
timestamp 1644511149
transform 1 0 15916 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1644511149
transform 1 0 20608 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0999_
timestamp 1644511149
transform 1 0 20608 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1000_
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1001_
timestamp 1644511149
transform 1 0 20884 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1003_
timestamp 1644511149
transform 1 0 20884 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1644511149
transform 1 0 23736 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1005_
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1006_
timestamp 1644511149
transform 1 0 22264 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1007_
timestamp 1644511149
transform 1 0 24380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1644511149
transform 1 0 25392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1009_
timestamp 1644511149
transform 1 0 23920 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1644511149
transform 1 0 25116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1011_
timestamp 1644511149
transform 1 0 23552 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1013_
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1644511149
transform 1 0 21988 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1015_
timestamp 1644511149
transform 1 0 24380 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1017_
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1644511149
transform 1 0 20976 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1019_
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1644511149
transform 1 0 20424 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1021_
timestamp 1644511149
transform 1 0 25944 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1023_
timestamp 1644511149
transform 1 0 25944 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1025_
timestamp 1644511149
transform 1 0 26772 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1027_
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1028_
timestamp 1644511149
transform 1 0 20700 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1029_
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1644511149
transform 1 0 18216 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1031_
timestamp 1644511149
transform 1 0 25576 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1032_
timestamp 1644511149
transform 1 0 26680 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1034_
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1644511149
transform 1 0 17848 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1036_
timestamp 1644511149
transform 1 0 8004 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1037_
timestamp 1644511149
transform 1 0 8004 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1038_
timestamp 1644511149
transform 1 0 10488 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1039_
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1040_
timestamp 1644511149
transform 1 0 8740 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1041_
timestamp 1644511149
transform 1 0 7544 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1042_
timestamp 1644511149
transform 1 0 7176 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1043_
timestamp 1644511149
transform 1 0 6256 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1044_
timestamp 1644511149
transform 1 0 7360 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1045_
timestamp 1644511149
transform 1 0 4140 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1046_
timestamp 1644511149
transform 1 0 4508 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1047_
timestamp 1644511149
transform 1 0 4784 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1048_
timestamp 1644511149
transform 1 0 8004 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1049_
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1050_
timestamp 1644511149
transform 1 0 4508 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1051_
timestamp 1644511149
transform 1 0 4048 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1052_
timestamp 1644511149
transform 1 0 16652 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1053_
timestamp 1644511149
transform 1 0 17112 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1054_
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1055_
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1056_
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1057_
timestamp 1644511149
transform 1 0 5612 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1058_
timestamp 1644511149
transform 1 0 3864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1059_
timestamp 1644511149
transform 1 0 4784 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1060_
timestamp 1644511149
transform 1 0 5428 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1061_
timestamp 1644511149
transform 1 0 5336 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1062_
timestamp 1644511149
transform 1 0 3864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1063_
timestamp 1644511149
transform 1 0 5336 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1064_
timestamp 1644511149
transform 1 0 4140 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1065_
timestamp 1644511149
transform 1 0 4968 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1066_
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1067_
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1068_
timestamp 1644511149
transform 1 0 1840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1069_
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1070_
timestamp 1644511149
transform 1 0 12236 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _1071_
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1072_
timestamp 1644511149
transform 1 0 9016 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1073_
timestamp 1644511149
transform 1 0 9292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1074_
timestamp 1644511149
transform 1 0 12512 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1075_
timestamp 1644511149
transform 1 0 8740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1076_
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1077_
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1078_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11868 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1079_
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1080_
timestamp 1644511149
transform 1 0 13064 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1081_
timestamp 1644511149
transform 1 0 10212 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1082_
timestamp 1644511149
transform 1 0 16468 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1083_
timestamp 1644511149
transform 1 0 13984 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1084_
timestamp 1644511149
transform 1 0 9752 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1085_
timestamp 1644511149
transform 1 0 8280 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1086_
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1087_
timestamp 1644511149
transform 1 0 9568 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1088_
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1089_
timestamp 1644511149
transform 1 0 13524 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1090_
timestamp 1644511149
transform 1 0 10580 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1091_
timestamp 1644511149
transform 1 0 11868 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1092_
timestamp 1644511149
transform 1 0 10120 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_2  _1093_
timestamp 1644511149
transform 1 0 9752 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1094_
timestamp 1644511149
transform 1 0 10304 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1095_
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1096_
timestamp 1644511149
transform 1 0 10304 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1097_
timestamp 1644511149
transform 1 0 13616 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1098_
timestamp 1644511149
transform 1 0 9384 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1099_
timestamp 1644511149
transform 1 0 11776 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1100_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8740 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1101_
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1102_
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1103_
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1104_
timestamp 1644511149
transform 1 0 12420 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1105_
timestamp 1644511149
transform 1 0 13248 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1106_
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1107_
timestamp 1644511149
transform 1 0 12972 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1108_
timestamp 1644511149
transform 1 0 15640 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1109_
timestamp 1644511149
transform 1 0 12972 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1110_
timestamp 1644511149
transform 1 0 13432 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1111_
timestamp 1644511149
transform 1 0 12328 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1112_
timestamp 1644511149
transform 1 0 7820 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1113_
timestamp 1644511149
transform 1 0 13892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1114_
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1115_
timestamp 1644511149
transform 1 0 14260 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1116_
timestamp 1644511149
transform 1 0 15088 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1117_
timestamp 1644511149
transform 1 0 14628 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1118_
timestamp 1644511149
transform 1 0 15640 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1119_
timestamp 1644511149
transform 1 0 14536 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1120_
timestamp 1644511149
transform 1 0 15364 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1121_
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1122_
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1123_
timestamp 1644511149
transform 1 0 15180 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1124_
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1125_
timestamp 1644511149
transform 1 0 14352 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1126_
timestamp 1644511149
transform 1 0 13248 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1127_
timestamp 1644511149
transform 1 0 15824 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1128_
timestamp 1644511149
transform 1 0 16744 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1129_
timestamp 1644511149
transform 1 0 17664 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1130_
timestamp 1644511149
transform 1 0 8096 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1131_
timestamp 1644511149
transform 1 0 16192 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1132_
timestamp 1644511149
transform 1 0 16744 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1133_
timestamp 1644511149
transform 1 0 16928 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1134_
timestamp 1644511149
transform 1 0 8004 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1135_
timestamp 1644511149
transform 1 0 5704 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1136_
timestamp 1644511149
transform 1 0 18584 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1137_
timestamp 1644511149
transform 1 0 19504 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1138_
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1139_
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1140_
timestamp 1644511149
transform 1 0 16928 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1141_
timestamp 1644511149
transform 1 0 17572 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1142_
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1143_
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1144_
timestamp 1644511149
transform 1 0 19596 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1145_
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1146_
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1147_
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1148_
timestamp 1644511149
transform 1 0 14996 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1149_
timestamp 1644511149
transform 1 0 9292 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1150_
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1151_
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1152_
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1153_
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1154_
timestamp 1644511149
transform 1 0 19872 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1155_
timestamp 1644511149
transform 1 0 5888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1156_
timestamp 1644511149
transform 1 0 10396 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1157_
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1158_
timestamp 1644511149
transform 1 0 7268 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1159_
timestamp 1644511149
transform 1 0 3956 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1160_
timestamp 1644511149
transform 1 0 2668 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1161_
timestamp 1644511149
transform 1 0 2576 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1162_
timestamp 1644511149
transform 1 0 2208 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1163_
timestamp 1644511149
transform 1 0 7544 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1164_
timestamp 1644511149
transform 1 0 8372 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1165_
timestamp 1644511149
transform 1 0 6532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1166_
timestamp 1644511149
transform 1 0 3404 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1167_
timestamp 1644511149
transform 1 0 2760 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1168_
timestamp 1644511149
transform 1 0 1656 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1169_
timestamp 1644511149
transform 1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1170_
timestamp 1644511149
transform 1 0 6716 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1171_
timestamp 1644511149
transform 1 0 6440 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1172_
timestamp 1644511149
transform 1 0 6348 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1173_
timestamp 1644511149
transform 1 0 7360 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1174_
timestamp 1644511149
transform 1 0 6716 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1175_
timestamp 1644511149
transform 1 0 3864 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1176_
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1177_
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1178_
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1179_
timestamp 1644511149
transform 1 0 5336 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1180_
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1181_
timestamp 1644511149
transform 1 0 5796 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1182_
timestamp 1644511149
transform 1 0 3772 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1183_
timestamp 1644511149
transform 1 0 2668 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1184_
timestamp 1644511149
transform 1 0 4416 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1185_
timestamp 1644511149
transform 1 0 7176 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1186_
timestamp 1644511149
transform 1 0 5060 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1187_
timestamp 1644511149
transform 1 0 5704 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1188_
timestamp 1644511149
transform 1 0 5060 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1189_
timestamp 1644511149
transform 1 0 3036 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1190_
timestamp 1644511149
transform 1 0 1840 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1191_
timestamp 1644511149
transform 1 0 1840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1192_
timestamp 1644511149
transform 1 0 5244 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1193_
timestamp 1644511149
transform 1 0 4416 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1194_
timestamp 1644511149
transform 1 0 3036 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1195_
timestamp 1644511149
transform 1 0 4232 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1196_
timestamp 1644511149
transform 1 0 2944 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1197_
timestamp 1644511149
transform 1 0 1840 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1198_
timestamp 1644511149
transform 1 0 1840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1199_
timestamp 1644511149
transform 1 0 5520 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1200_
timestamp 1644511149
transform 1 0 6532 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1201_
timestamp 1644511149
transform 1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1202_
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1203_
timestamp 1644511149
transform 1 0 2668 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1204_
timestamp 1644511149
transform 1 0 1932 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1205_
timestamp 1644511149
transform 1 0 3312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1206_
timestamp 1644511149
transform 1 0 7176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1207_
timestamp 1644511149
transform 1 0 6532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1208_
timestamp 1644511149
transform 1 0 5244 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1209_
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1210_
timestamp 1644511149
transform 1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1211_
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1212_
timestamp 1644511149
transform 1 0 5060 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1213_
timestamp 1644511149
transform 1 0 5060 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1214_
timestamp 1644511149
transform 1 0 6900 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1215_
timestamp 1644511149
transform 1 0 6624 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1216_
timestamp 1644511149
transform 1 0 7636 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1217_
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1218_
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1219_
timestamp 1644511149
transform 1 0 1840 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1220_
timestamp 1644511149
transform 1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1221_
timestamp 1644511149
transform 1 0 7544 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1222_
timestamp 1644511149
transform 1 0 5152 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1223_
timestamp 1644511149
transform 1 0 4692 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1224_
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1225_
timestamp 1644511149
transform 1 0 3772 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1226_
timestamp 1644511149
transform 1 0 2668 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1227_
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1228_
timestamp 1644511149
transform 1 0 4692 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1229_
timestamp 1644511149
transform 1 0 5520 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1230_
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1231_
timestamp 1644511149
transform 1 0 8372 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1232_
timestamp 1644511149
transform 1 0 6440 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1233_
timestamp 1644511149
transform 1 0 4968 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1234_
timestamp 1644511149
transform 1 0 5336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1235_
timestamp 1644511149
transform 1 0 6716 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1236_
timestamp 1644511149
transform 1 0 7728 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1237_
timestamp 1644511149
transform 1 0 6348 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1238_
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1239_
timestamp 1644511149
transform 1 0 6624 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1240_
timestamp 1644511149
transform 1 0 6624 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1241_
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1242_
timestamp 1644511149
transform 1 0 10212 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1243_
timestamp 1644511149
transform 1 0 10120 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1244_
timestamp 1644511149
transform 1 0 10028 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1245_
timestamp 1644511149
transform 1 0 7912 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1246_
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1247_
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1248_
timestamp 1644511149
transform 1 0 7820 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1249_
timestamp 1644511149
transform 1 0 2392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1250_
timestamp 1644511149
transform 1 0 9568 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1251_
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1252_
timestamp 1644511149
transform 1 0 1564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1253_
timestamp 1644511149
transform 1 0 9108 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1254_
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1255_
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1256_
timestamp 1644511149
transform 1 0 13248 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1257_
timestamp 1644511149
transform 1 0 10120 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1258_
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1259_
timestamp 1644511149
transform 1 0 3312 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1260_
timestamp 1644511149
transform 1 0 9936 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1261_
timestamp 1644511149
transform 1 0 10120 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1262_
timestamp 1644511149
transform 1 0 1840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1263_
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1264_
timestamp 1644511149
transform 1 0 12512 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1265_
timestamp 1644511149
transform 1 0 2392 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1266_
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1267_
timestamp 1644511149
transform 1 0 10120 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1268_
timestamp 1644511149
transform 1 0 12420 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1269_
timestamp 1644511149
transform 1 0 11408 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1270_
timestamp 1644511149
transform 1 0 12420 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1271_
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1272_
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1273_
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1274_
timestamp 1644511149
transform 1 0 9752 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1275_
timestamp 1644511149
transform 1 0 10856 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1276_
timestamp 1644511149
transform 1 0 9200 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1277_
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1278_
timestamp 1644511149
transform 1 0 19596 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1279_
timestamp 1644511149
transform 1 0 17664 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1280_
timestamp 1644511149
transform 1 0 11868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1281_
timestamp 1644511149
transform 1 0 9200 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1282_
timestamp 1644511149
transform 1 0 4416 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1283_
timestamp 1644511149
transform 1 0 9384 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1284_
timestamp 1644511149
transform 1 0 9568 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1285_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_2  _1286_
timestamp 1644511149
transform 1 0 9016 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1287_
timestamp 1644511149
transform 1 0 14168 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1288_
timestamp 1644511149
transform 1 0 14904 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _1289_
timestamp 1644511149
transform 1 0 14352 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1290_
timestamp 1644511149
transform 1 0 8832 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1291_
timestamp 1644511149
transform 1 0 10120 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1292_
timestamp 1644511149
transform 1 0 5520 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1293_
timestamp 1644511149
transform 1 0 8648 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1294_
timestamp 1644511149
transform 1 0 10396 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1295_
timestamp 1644511149
transform 1 0 11040 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1296_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9936 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1297_
timestamp 1644511149
transform 1 0 7912 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1298_
timestamp 1644511149
transform 1 0 6716 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1299_
timestamp 1644511149
transform 1 0 9568 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _1300_
timestamp 1644511149
transform 1 0 7544 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1301_
timestamp 1644511149
transform 1 0 14996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1302_
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1303_
timestamp 1644511149
transform 1 0 7636 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1304_
timestamp 1644511149
transform 1 0 9844 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1305_
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1306_
timestamp 1644511149
transform 1 0 9016 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1307_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7452 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _1308_
timestamp 1644511149
transform 1 0 7544 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1309_
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1310_
timestamp 1644511149
transform 1 0 6624 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1311_
timestamp 1644511149
transform 1 0 8188 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1312_
timestamp 1644511149
transform 1 0 5520 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1313_
timestamp 1644511149
transform 1 0 7728 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1314_
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1315_
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1316_
timestamp 1644511149
transform 1 0 4140 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1317_
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1318_
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1319_
timestamp 1644511149
transform 1 0 6716 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1320_
timestamp 1644511149
transform 1 0 5888 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _1321_
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1322_
timestamp 1644511149
transform 1 0 5704 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1323_
timestamp 1644511149
transform 1 0 5244 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1324_
timestamp 1644511149
transform 1 0 5244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1325_
timestamp 1644511149
transform 1 0 3404 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1326_
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1327_
timestamp 1644511149
transform 1 0 3036 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1328_
timestamp 1644511149
transform 1 0 4600 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1329_
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1330_
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1331_
timestamp 1644511149
transform 1 0 2760 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1332_
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _1333_
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1334_
timestamp 1644511149
transform 1 0 3220 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1335_
timestamp 1644511149
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _1336_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3404 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _1337_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5704 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1338_
timestamp 1644511149
transform 1 0 4692 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1339_
timestamp 1644511149
transform 1 0 4508 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1340_
timestamp 1644511149
transform 1 0 5152 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1341_
timestamp 1644511149
transform 1 0 3956 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1342_
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_1  _1343_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7360 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1344_
timestamp 1644511149
transform 1 0 9016 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1345_
timestamp 1644511149
transform 1 0 8096 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1346_
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _1347_
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1348_
timestamp 1644511149
transform 1 0 9384 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _1349_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _1350_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10856 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _1351_
timestamp 1644511149
transform 1 0 19596 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1352_
timestamp 1644511149
transform 1 0 19412 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _1353_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1354_
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1355_
timestamp 1644511149
transform 1 0 17940 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1356_
timestamp 1644511149
transform 1 0 17848 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1357_
timestamp 1644511149
transform 1 0 17756 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1358_
timestamp 1644511149
transform 1 0 17572 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1359_
timestamp 1644511149
transform 1 0 17388 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1360_
timestamp 1644511149
transform 1 0 18124 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1361_
timestamp 1644511149
transform 1 0 22816 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1362_
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1363_
timestamp 1644511149
transform 1 0 19412 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1364_
timestamp 1644511149
transform 1 0 20424 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1365_
timestamp 1644511149
transform 1 0 20700 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1366_
timestamp 1644511149
transform 1 0 19688 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1367_
timestamp 1644511149
transform 1 0 27048 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1368_
timestamp 1644511149
transform 1 0 23736 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1369_
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1370_
timestamp 1644511149
transform 1 0 23184 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1371_
timestamp 1644511149
transform 1 0 21160 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1372_
timestamp 1644511149
transform 1 0 23092 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1373_
timestamp 1644511149
transform 1 0 23000 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1374_
timestamp 1644511149
transform 1 0 24196 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1375_
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1376_
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1377_
timestamp 1644511149
transform 1 0 25668 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1378_
timestamp 1644511149
transform 1 0 24196 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1379_
timestamp 1644511149
transform 1 0 25024 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1380_
timestamp 1644511149
transform 1 0 26220 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1381_
timestamp 1644511149
transform 1 0 23552 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1382_
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1383_
timestamp 1644511149
transform 1 0 24932 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1384_
timestamp 1644511149
transform 1 0 25944 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1385_
timestamp 1644511149
transform 1 0 25484 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1386_
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1387_
timestamp 1644511149
transform 1 0 24748 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1388_
timestamp 1644511149
transform 1 0 25024 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1389_
timestamp 1644511149
transform 1 0 23736 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1390_
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1391_
timestamp 1644511149
transform 1 0 22540 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1392_
timestamp 1644511149
transform 1 0 26312 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1393_
timestamp 1644511149
transform 1 0 21988 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1394_
timestamp 1644511149
transform 1 0 23276 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1395_
timestamp 1644511149
transform 1 0 12696 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1396_
timestamp 1644511149
transform 1 0 14904 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1397_
timestamp 1644511149
transform 1 0 15732 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1398_
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1399_
timestamp 1644511149
transform 1 0 19412 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1400_
timestamp 1644511149
transform 1 0 11868 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1401_
timestamp 1644511149
transform 1 0 3036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1402_
timestamp 1644511149
transform 1 0 15732 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1403_
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1404_
timestamp 1644511149
transform 1 0 16928 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1405_
timestamp 1644511149
transform 1 0 18032 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1406_
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1407_
timestamp 1644511149
transform 1 0 14260 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1408_
timestamp 1644511149
transform 1 0 21068 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1409_
timestamp 1644511149
transform 1 0 19688 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1410_
timestamp 1644511149
transform 1 0 23276 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1411_
timestamp 1644511149
transform 1 0 1564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1412_
timestamp 1644511149
transform 1 0 22172 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1413_
timestamp 1644511149
transform 1 0 16836 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1414_
timestamp 1644511149
transform 1 0 21620 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1415_
timestamp 1644511149
transform 1 0 16744 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1416_
timestamp 1644511149
transform 1 0 27140 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1417_
timestamp 1644511149
transform 1 0 22632 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1418_
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1419_
timestamp 1644511149
transform 1 0 19320 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1420_
timestamp 1644511149
transform 1 0 26220 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1421_
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1422_
timestamp 1644511149
transform 1 0 17848 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1423_
timestamp 1644511149
transform 1 0 14812 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1424_
timestamp 1644511149
transform 1 0 21620 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1425_
timestamp 1644511149
transform 1 0 19412 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1426_
timestamp 1644511149
transform 1 0 20424 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1427_
timestamp 1644511149
transform 1 0 15548 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1428_
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1429_
timestamp 1644511149
transform 1 0 18216 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1430_
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1431_
timestamp 1644511149
transform 1 0 20240 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1432_
timestamp 1644511149
transform 1 0 22264 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1433_
timestamp 1644511149
transform 1 0 21712 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1434_
timestamp 1644511149
transform 1 0 22264 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1435_
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1436_
timestamp 1644511149
transform 1 0 20608 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1437_
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1438_
timestamp 1644511149
transform 1 0 23000 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1439_
timestamp 1644511149
transform 1 0 22080 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1440_
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1441_
timestamp 1644511149
transform 1 0 22908 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1442_
timestamp 1644511149
transform 1 0 27140 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1443_
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1444_
timestamp 1644511149
transform 1 0 23736 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1445_
timestamp 1644511149
transform 1 0 25576 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1446_
timestamp 1644511149
transform 1 0 24380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1447_
timestamp 1644511149
transform 1 0 24564 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1448_
timestamp 1644511149
transform 1 0 26128 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1449_
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1450_
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1451_
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1452_
timestamp 1644511149
transform 1 0 25484 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1453_
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1454_
timestamp 1644511149
transform 1 0 26220 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1455_
timestamp 1644511149
transform 1 0 26680 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1456_
timestamp 1644511149
transform 1 0 26036 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1457_
timestamp 1644511149
transform 1 0 21160 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1458_
timestamp 1644511149
transform 1 0 26404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1459_
timestamp 1644511149
transform 1 0 2944 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1460_
timestamp 1644511149
transform 1 0 15456 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1461_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15364 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1462_
timestamp 1644511149
transform 1 0 12696 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1463_
timestamp 1644511149
transform 1 0 14720 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1464_
timestamp 1644511149
transform 1 0 15916 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1465_
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1466_
timestamp 1644511149
transform 1 0 15640 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1467_
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1468_
timestamp 1644511149
transform 1 0 13156 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1469_
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1470_
timestamp 1644511149
transform 1 0 13524 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1471_
timestamp 1644511149
transform 1 0 10488 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1472_
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1473_
timestamp 1644511149
transform 1 0 11408 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1474_
timestamp 1644511149
transform 1 0 7636 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1475_
timestamp 1644511149
transform 1 0 10580 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1476_
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1477_
timestamp 1644511149
transform 1 0 2300 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1478_
timestamp 1644511149
transform 1 0 6440 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1479_
timestamp 1644511149
transform 1 0 10672 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1480_
timestamp 1644511149
transform 1 0 10672 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1481_
timestamp 1644511149
transform 1 0 13156 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _1482_
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1483_
timestamp 1644511149
transform 1 0 12512 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1484_
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1485_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1486_
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1487_
timestamp 1644511149
transform 1 0 12144 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1488_
timestamp 1644511149
transform 1 0 12604 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1489_
timestamp 1644511149
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1490_
timestamp 1644511149
transform 1 0 13248 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1491_
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1492_
timestamp 1644511149
transform 1 0 12972 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1493_
timestamp 1644511149
transform 1 0 12880 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1494_
timestamp 1644511149
transform 1 0 12788 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1495_
timestamp 1644511149
transform 1 0 12512 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1496_
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a311oi_1  _1497_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1498_
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1499_
timestamp 1644511149
transform 1 0 12972 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1500_
timestamp 1644511149
transform 1 0 12420 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1501_
timestamp 1644511149
transform 1 0 11960 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1502_
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1503_
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1504_
timestamp 1644511149
transform 1 0 11500 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1505_
timestamp 1644511149
transform 1 0 12144 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1506_
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1507_
timestamp 1644511149
transform 1 0 17848 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1508_
timestamp 1644511149
transform 1 0 23736 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1509_
timestamp 1644511149
transform 1 0 15456 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1510_
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1511_
timestamp 1644511149
transform 1 0 18492 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1512_
timestamp 1644511149
transform 1 0 18676 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1513_
timestamp 1644511149
transform 1 0 15732 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1514_
timestamp 1644511149
transform 1 0 17388 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1515_
timestamp 1644511149
transform 1 0 17572 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1516_
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1517_
timestamp 1644511149
transform 1 0 15640 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1518_
timestamp 1644511149
transform 1 0 20700 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1519_
timestamp 1644511149
transform 1 0 17848 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1520_
timestamp 1644511149
transform 1 0 17572 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1521_
timestamp 1644511149
transform 1 0 15456 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1522_
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1523_
timestamp 1644511149
transform 1 0 20424 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1524_
timestamp 1644511149
transform 1 0 27048 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1525_
timestamp 1644511149
transform 1 0 19596 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1526_
timestamp 1644511149
transform 1 0 18768 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1527_
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1528_
timestamp 1644511149
transform 1 0 18492 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1529_
timestamp 1644511149
transform 1 0 18308 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1530_
timestamp 1644511149
transform 1 0 17940 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1531_
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1532_
timestamp 1644511149
transform 1 0 19872 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1533_
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1534_
timestamp 1644511149
transform 1 0 18676 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1535_
timestamp 1644511149
transform 1 0 20332 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1536_
timestamp 1644511149
transform 1 0 19504 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1537_
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1538_
timestamp 1644511149
transform 1 0 19688 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1539_
timestamp 1644511149
transform 1 0 19412 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1540_
timestamp 1644511149
transform 1 0 20240 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1541_
timestamp 1644511149
transform 1 0 22448 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1542_
timestamp 1644511149
transform 1 0 23000 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1543_
timestamp 1644511149
transform 1 0 23092 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1544_
timestamp 1644511149
transform 1 0 22724 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1545_
timestamp 1644511149
transform 1 0 21988 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1546_
timestamp 1644511149
transform 1 0 23276 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1547_
timestamp 1644511149
transform 1 0 21804 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1548_
timestamp 1644511149
transform 1 0 21344 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1549_
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1550_
timestamp 1644511149
transform 1 0 18768 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1551_
timestamp 1644511149
transform 1 0 24380 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1552_
timestamp 1644511149
transform 1 0 21068 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1553_
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1554_
timestamp 1644511149
transform 1 0 21068 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1555_
timestamp 1644511149
transform 1 0 22356 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1556_
timestamp 1644511149
transform 1 0 23736 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1557_
timestamp 1644511149
transform 1 0 22264 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1558_
timestamp 1644511149
transform 1 0 23000 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1559_
timestamp 1644511149
transform 1 0 23184 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1560_
timestamp 1644511149
transform 1 0 24196 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1561_
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1562_
timestamp 1644511149
transform 1 0 25576 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1563_
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1564_
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1565_
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1566_
timestamp 1644511149
transform 1 0 25024 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1567_
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1568_
timestamp 1644511149
transform 1 0 23184 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1569_
timestamp 1644511149
transform 1 0 25024 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1570_
timestamp 1644511149
transform 1 0 24564 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1571_
timestamp 1644511149
transform 1 0 25116 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1572_
timestamp 1644511149
transform 1 0 26864 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1573_
timestamp 1644511149
transform 1 0 24288 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1574_
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1575_
timestamp 1644511149
transform 1 0 25116 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1576_
timestamp 1644511149
transform 1 0 23644 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1577_
timestamp 1644511149
transform 1 0 25668 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1578_
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1579_
timestamp 1644511149
transform 1 0 26404 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1580_
timestamp 1644511149
transform 1 0 21988 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1581_
timestamp 1644511149
transform 1 0 24472 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1582_
timestamp 1644511149
transform 1 0 25116 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1583_
timestamp 1644511149
transform 1 0 26680 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1584_
timestamp 1644511149
transform 1 0 25760 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1585_
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1586_
timestamp 1644511149
transform 1 0 24748 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1587_
timestamp 1644511149
transform 1 0 25300 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1588_
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1589_
timestamp 1644511149
transform 1 0 27140 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1590_
timestamp 1644511149
transform 1 0 22264 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1591_
timestamp 1644511149
transform 1 0 23644 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1592_
timestamp 1644511149
transform 1 0 23920 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1593_
timestamp 1644511149
transform 1 0 23460 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1594_
timestamp 1644511149
transform 1 0 25024 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1595_
timestamp 1644511149
transform 1 0 23276 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1596_
timestamp 1644511149
transform 1 0 24748 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1597_
timestamp 1644511149
transform 1 0 25116 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1598_
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1599_
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1600_
timestamp 1644511149
transform 1 0 20792 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1601_
timestamp 1644511149
transform 1 0 23092 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1602_
timestamp 1644511149
transform 1 0 23276 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1603_
timestamp 1644511149
transform 1 0 23368 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1604_
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1605_
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1606_
timestamp 1644511149
transform 1 0 13064 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1607_
timestamp 1644511149
transform 1 0 10856 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1608_
timestamp 1644511149
transform 1 0 14904 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1609_
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1610_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1611_
timestamp 1644511149
transform 1 0 1840 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1612_
timestamp 1644511149
transform 1 0 6992 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1613_
timestamp 1644511149
transform 1 0 1932 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1614_
timestamp 1644511149
transform 1 0 5612 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1615_
timestamp 1644511149
transform 1 0 1932 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1616_
timestamp 1644511149
transform 1 0 4048 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1617_
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1618_
timestamp 1644511149
transform 1 0 1840 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1619_
timestamp 1644511149
transform 1 0 3128 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1620_
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1621_
timestamp 1644511149
transform 1 0 10120 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1622_
timestamp 1644511149
transform 1 0 8740 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1623_
timestamp 1644511149
transform 1 0 9476 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1624_
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1625_
timestamp 1644511149
transform 1 0 12788 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1626_
timestamp 1644511149
transform 1 0 13156 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1627_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14260 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1628_
timestamp 1644511149
transform 1 0 14628 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1629_
timestamp 1644511149
transform 1 0 14996 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1630_
timestamp 1644511149
transform 1 0 16652 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1631_
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1632_
timestamp 1644511149
transform 1 0 17296 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1633_
timestamp 1644511149
transform 1 0 17296 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1634_
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1635_
timestamp 1644511149
transform 1 0 17204 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1636_
timestamp 1644511149
transform 1 0 20424 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1637_
timestamp 1644511149
transform 1 0 20148 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1638_
timestamp 1644511149
transform 1 0 19688 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1639_
timestamp 1644511149
transform 1 0 20516 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1640_
timestamp 1644511149
transform 1 0 7728 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1641_
timestamp 1644511149
transform 1 0 1748 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1642_
timestamp 1644511149
transform 1 0 6532 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1643_
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1644_
timestamp 1644511149
transform 1 0 6440 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1645_
timestamp 1644511149
transform 1 0 1564 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1646_
timestamp 1644511149
transform 1 0 4416 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1647_
timestamp 1644511149
transform 1 0 2576 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1648_
timestamp 1644511149
transform 1 0 3956 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1649_
timestamp 1644511149
transform 1 0 1656 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1650_
timestamp 1644511149
transform 1 0 3864 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1651_
timestamp 1644511149
transform 1 0 1564 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1652_
timestamp 1644511149
transform 1 0 3864 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1653_
timestamp 1644511149
transform 1 0 1472 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1654_
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1655_
timestamp 1644511149
transform 1 0 4048 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1656_
timestamp 1644511149
transform 1 0 6900 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1657_
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1658_
timestamp 1644511149
transform 1 0 1472 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1659_
timestamp 1644511149
transform 1 0 2576 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1660_
timestamp 1644511149
transform 1 0 3312 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1661_
timestamp 1644511149
transform 1 0 5060 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1662_
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1663_
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1664_
timestamp 1644511149
transform 1 0 8188 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1665_
timestamp 1644511149
transform 1 0 7820 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1666_
timestamp 1644511149
transform 1 0 8280 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1667_
timestamp 1644511149
transform 1 0 8188 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1668_
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1669_
timestamp 1644511149
transform 1 0 10488 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1670_
timestamp 1644511149
transform 1 0 12144 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1671_
timestamp 1644511149
transform 1 0 10396 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1672_
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1673_
timestamp 1644511149
transform 1 0 13432 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1674_
timestamp 1644511149
transform 1 0 10304 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1675_
timestamp 1644511149
transform 1 0 12052 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1676_
timestamp 1644511149
transform 1 0 9568 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1677_
timestamp 1644511149
transform 1 0 10304 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1678_
timestamp 1644511149
transform 1 0 7176 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1679_
timestamp 1644511149
transform 1 0 6440 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1680_
timestamp 1644511149
transform 1 0 4416 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1681_
timestamp 1644511149
transform 1 0 3772 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1682_
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1683_
timestamp 1644511149
transform 1 0 1840 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1684_
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1685_
timestamp 1644511149
transform 1 0 17940 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1686_
timestamp 1644511149
transform 1 0 17296 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1687_
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1688_
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1689_
timestamp 1644511149
transform 1 0 19780 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1690_
timestamp 1644511149
transform 1 0 21896 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1691_
timestamp 1644511149
transform 1 0 21988 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1692_
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1693_
timestamp 1644511149
transform 1 0 25944 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1694_
timestamp 1644511149
transform 1 0 25944 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1695_
timestamp 1644511149
transform 1 0 25944 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1696_
timestamp 1644511149
transform 1 0 25944 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1697_
timestamp 1644511149
transform 1 0 25024 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1698_
timestamp 1644511149
transform 1 0 23644 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1699_
timestamp 1644511149
transform 1 0 25944 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1700_
timestamp 1644511149
transform 1 0 22356 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1701_
timestamp 1644511149
transform 1 0 13064 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1702_
timestamp 1644511149
transform 1 0 11684 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1703_
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1704_
timestamp 1644511149
transform 1 0 18308 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1705_
timestamp 1644511149
transform 1 0 14260 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1706_
timestamp 1644511149
transform 1 0 20148 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1707_
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1708_
timestamp 1644511149
transform 1 0 16744 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1709_
timestamp 1644511149
transform 1 0 23644 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1710_
timestamp 1644511149
transform 1 0 20148 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1711_
timestamp 1644511149
transform 1 0 24932 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1712_
timestamp 1644511149
transform 1 0 18124 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1713_
timestamp 1644511149
transform 1 0 22080 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 1644511149
transform 1 0 20240 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 1644511149
transform 1 0 16192 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1716_
timestamp 1644511149
transform 1 0 17296 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1717_
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1718_
timestamp 1644511149
transform 1 0 21068 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1719_
timestamp 1644511149
transform 1 0 19872 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 1644511149
transform 1 0 22080 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1721_
timestamp 1644511149
transform 1 0 22080 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1722_
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1723_
timestamp 1644511149
transform 1 0 22448 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1724_
timestamp 1644511149
transform 1 0 24564 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1725_
timestamp 1644511149
transform 1 0 24472 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1726_
timestamp 1644511149
transform 1 0 24104 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1727_
timestamp 1644511149
transform 1 0 24748 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1728_
timestamp 1644511149
transform 1 0 24840 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1729_
timestamp 1644511149
transform 1 0 25944 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1730_
timestamp 1644511149
transform 1 0 25944 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1731_
timestamp 1644511149
transform 1 0 25944 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1732_
timestamp 1644511149
transform 1 0 25024 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1733_
timestamp 1644511149
transform 1 0 9568 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1734_
timestamp 1644511149
transform 1 0 14996 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1735_
timestamp 1644511149
transform 1 0 14720 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1736_
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1737_
timestamp 1644511149
transform 1 0 15456 0 1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1738_
timestamp 1644511149
transform 1 0 13892 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1739_
timestamp 1644511149
transform 1 0 8924 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1740_
timestamp 1644511149
transform 1 0 5428 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1741_
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1742_
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1743_
timestamp 1644511149
transform 1 0 11592 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1744_
timestamp 1644511149
transform 1 0 10580 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1745_
timestamp 1644511149
transform 1 0 14260 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1746_
timestamp 1644511149
transform 1 0 11868 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1747_
timestamp 1644511149
transform 1 0 14444 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1748_
timestamp 1644511149
transform 1 0 11040 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1749_
timestamp 1644511149
transform 1 0 12236 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1750_
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1751_
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1752_
timestamp 1644511149
transform 1 0 18492 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1753_
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1754_
timestamp 1644511149
transform 1 0 19872 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1755_
timestamp 1644511149
transform 1 0 21804 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1756_
timestamp 1644511149
transform 1 0 21896 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1757_
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1758_
timestamp 1644511149
transform 1 0 25392 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1759_
timestamp 1644511149
transform 1 0 25944 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1760_
timestamp 1644511149
transform 1 0 25944 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1761_
timestamp 1644511149
transform 1 0 25944 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1762_
timestamp 1644511149
transform 1 0 25944 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1763_
timestamp 1644511149
transform 1 0 24748 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1764_
timestamp 1644511149
transform 1 0 25024 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1765_
timestamp 1644511149
transform 1 0 23000 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1766_
timestamp 1644511149
transform 1 0 13064 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1767_
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1768__90 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2576 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1769__91
timestamp 1644511149
transform 1 0 4416 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CLK pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14352 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_CLK
timestamp 1644511149
transform 1 0 6532 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_CLK
timestamp 1644511149
transform 1 0 10488 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_CLK
timestamp 1644511149
transform 1 0 4140 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_CLK
timestamp 1644511149
transform 1 0 9016 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_CLK
timestamp 1644511149
transform 1 0 18400 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_CLK
timestamp 1644511149
transform 1 0 21620 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_CLK
timestamp 1644511149
transform 1 0 20056 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_CLK
timestamp 1644511149
transform 1 0 20976 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_CLK
timestamp 1644511149
transform 1 0 4508 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_CLK
timestamp 1644511149
transform 1 0 4324 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_CLK
timestamp 1644511149
transform 1 0 12512 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_CLK
timestamp 1644511149
transform 1 0 15088 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_CLK
timestamp 1644511149
transform 1 0 4692 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_CLK
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_CLK
timestamp 1644511149
transform 1 0 10580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_CLK
timestamp 1644511149
transform 1 0 10856 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_CLK
timestamp 1644511149
transform 1 0 17480 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_CLK
timestamp 1644511149
transform 1 0 17572 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_CLK
timestamp 1644511149
transform 1 0 23000 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_CLK
timestamp 1644511149
transform 1 0 23552 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_CLK
timestamp 1644511149
transform 1 0 18492 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_CLK
timestamp 1644511149
transform 1 0 17020 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_CLK
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_CLK
timestamp 1644511149
transform 1 0 26128 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 1656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1644511149
transform 1 0 1840 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform 1 0 3036 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1644511149
transform 1 0 2944 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1644511149
transform 1 0 2392 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform 1 0 1748 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1644511149
transform 1 0 5612 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform 1 0 2300 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform 1 0 3036 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1644511149
transform 1 0 3404 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform 1 0 3404 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform 1 0 3404 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1644511149
transform 1 0 1656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform 1 0 1840 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform 1 0 2392 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1644511149
transform 1 0 2392 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform 1 0 1564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform 1 0 12144 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform 1 0 1748 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 2852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 2116 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1644511149
transform 1 0 2392 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1644511149
transform 1 0 1472 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 1748 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 1748 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 1932 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 2208 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform 1 0 2392 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 1564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1644511149
transform 1 0 1748 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1644511149
transform 1 0 3036 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1644511149
transform 1 0 17204 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1644511149
transform 1 0 20056 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1644511149
transform 1 0 15916 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1644511149
transform 1 0 20700 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1644511149
transform 1 0 20976 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1644511149
transform 1 0 22448 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1644511149
transform 1 0 10764 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform 1 0 15824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1644511149
transform 1 0 14812 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1644511149
transform 1 0 17296 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1644511149
transform 1 0 23092 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1644511149
transform 1 0 2116 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1644511149
transform 1 0 10120 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform 1 0 23644 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1644511149
transform 1 0 27048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp 1644511149
transform 1 0 26128 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1644511149
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1644511149
transform 1 0 13248 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1644511149
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1644511149
transform 1 0 19964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1644511149
transform 1 0 19596 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1644511149
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1644511149
transform 1 0 23368 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1644511149
transform 1 0 25116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1644511149
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1644511149
transform 1 0 22816 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1644511149
transform 1 0 25300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1644511149
transform 1 0 23552 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1644511149
transform 1 0 25208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1644511149
transform 1 0 25208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1644511149
transform 1 0 20976 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1644511149
transform 1 0 23552 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1644511149
transform 1 0 27048 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1644511149
transform 1 0 13340 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1644511149
transform 1 0 22816 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1644511149
transform 1 0 19504 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1644511149
transform 1 0 14076 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1644511149
transform 1 0 14720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1644511149
transform 1 0 15456 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1644511149
transform 1 0 17572 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1644511149
transform 1 0 18308 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1644511149
transform 1 0 27048 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1644511149
transform 1 0 27048 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1644511149
transform 1 0 27048 0 1 27200
box -38 -48 406 592
<< labels >>
rlabel metal2 s 110 0 166 800 6 CLK
port 0 nsew signal input
rlabel metal2 s 294 0 350 800 6 RST_N
port 1 nsew signal input
rlabel metal4 s 9930 2128 10250 28880 6 VGND
port 2 nsew ground input
rlabel metal4 s 18915 2128 19235 28880 6 VGND
port 2 nsew ground input
rlabel metal4 s 5436 2128 5756 28880 6 VPWR
port 3 nsew power input
rlabel metal4 s 14422 2128 14742 28880 6 VPWR
port 3 nsew power input
rlabel metal4 s 23407 2128 23727 28880 6 VPWR
port 3 nsew power input
rlabel metal2 s 2226 0 2282 800 6 slave_ack_o
port 4 nsew signal tristate
rlabel metal2 s 3054 0 3110 800 6 slave_adr_i[0]
port 5 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 slave_adr_i[10]
port 6 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 slave_adr_i[11]
port 7 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 slave_adr_i[12]
port 8 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 slave_adr_i[13]
port 9 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 slave_adr_i[14]
port 10 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 slave_adr_i[15]
port 11 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 slave_adr_i[16]
port 12 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 slave_adr_i[17]
port 13 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 slave_adr_i[18]
port 14 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 slave_adr_i[19]
port 15 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 slave_adr_i[1]
port 16 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 slave_adr_i[20]
port 17 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 slave_adr_i[21]
port 18 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 slave_adr_i[22]
port 19 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 slave_adr_i[23]
port 20 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 slave_adr_i[24]
port 21 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 slave_adr_i[25]
port 22 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 slave_adr_i[26]
port 23 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 slave_adr_i[27]
port 24 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 slave_adr_i[28]
port 25 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 slave_adr_i[29]
port 26 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 slave_adr_i[2]
port 27 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 slave_adr_i[30]
port 28 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 slave_adr_i[31]
port 29 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 slave_adr_i[3]
port 30 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 slave_adr_i[4]
port 31 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 slave_adr_i[5]
port 32 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 slave_adr_i[6]
port 33 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 slave_adr_i[7]
port 34 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 slave_adr_i[8]
port 35 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 slave_adr_i[9]
port 36 nsew signal input
rlabel metal2 s 570 0 626 800 6 slave_cyc_i
port 37 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 slave_dat_i[0]
port 38 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 slave_dat_i[10]
port 39 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 slave_dat_i[11]
port 40 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 slave_dat_i[12]
port 41 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 slave_dat_i[13]
port 42 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 slave_dat_i[14]
port 43 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 slave_dat_i[15]
port 44 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 slave_dat_i[16]
port 45 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 slave_dat_i[17]
port 46 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 slave_dat_i[18]
port 47 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 slave_dat_i[19]
port 48 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 slave_dat_i[1]
port 49 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 slave_dat_i[20]
port 50 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 slave_dat_i[21]
port 51 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 slave_dat_i[22]
port 52 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 slave_dat_i[23]
port 53 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 slave_dat_i[24]
port 54 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 slave_dat_i[25]
port 55 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 slave_dat_i[26]
port 56 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 slave_dat_i[27]
port 57 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 slave_dat_i[28]
port 58 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 slave_dat_i[29]
port 59 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 slave_dat_i[2]
port 60 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 slave_dat_i[30]
port 61 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 slave_dat_i[31]
port 62 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 slave_dat_i[3]
port 63 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 slave_dat_i[4]
port 64 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 slave_dat_i[5]
port 65 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 slave_dat_i[6]
port 66 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 slave_dat_i[7]
port 67 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 slave_dat_i[8]
port 68 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 slave_dat_i[9]
port 69 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 slave_dat_o[0]
port 70 nsew signal tristate
rlabel metal2 s 17314 0 17370 800 6 slave_dat_o[10]
port 71 nsew signal tristate
rlabel metal2 s 17866 0 17922 800 6 slave_dat_o[11]
port 72 nsew signal tristate
rlabel metal2 s 18418 0 18474 800 6 slave_dat_o[12]
port 73 nsew signal tristate
rlabel metal2 s 18970 0 19026 800 6 slave_dat_o[13]
port 74 nsew signal tristate
rlabel metal2 s 19522 0 19578 800 6 slave_dat_o[14]
port 75 nsew signal tristate
rlabel metal2 s 20074 0 20130 800 6 slave_dat_o[15]
port 76 nsew signal tristate
rlabel metal2 s 20626 0 20682 800 6 slave_dat_o[16]
port 77 nsew signal tristate
rlabel metal2 s 21086 0 21142 800 6 slave_dat_o[17]
port 78 nsew signal tristate
rlabel metal2 s 21638 0 21694 800 6 slave_dat_o[18]
port 79 nsew signal tristate
rlabel metal2 s 22190 0 22246 800 6 slave_dat_o[19]
port 80 nsew signal tristate
rlabel metal2 s 12530 0 12586 800 6 slave_dat_o[1]
port 81 nsew signal tristate
rlabel metal2 s 22742 0 22798 800 6 slave_dat_o[20]
port 82 nsew signal tristate
rlabel metal2 s 23294 0 23350 800 6 slave_dat_o[21]
port 83 nsew signal tristate
rlabel metal2 s 23846 0 23902 800 6 slave_dat_o[22]
port 84 nsew signal tristate
rlabel metal2 s 24398 0 24454 800 6 slave_dat_o[23]
port 85 nsew signal tristate
rlabel metal2 s 24950 0 25006 800 6 slave_dat_o[24]
port 86 nsew signal tristate
rlabel metal2 s 25410 0 25466 800 6 slave_dat_o[25]
port 87 nsew signal tristate
rlabel metal2 s 25962 0 26018 800 6 slave_dat_o[26]
port 88 nsew signal tristate
rlabel metal2 s 26514 0 26570 800 6 slave_dat_o[27]
port 89 nsew signal tristate
rlabel metal2 s 27066 0 27122 800 6 slave_dat_o[28]
port 90 nsew signal tristate
rlabel metal2 s 27618 0 27674 800 6 slave_dat_o[29]
port 91 nsew signal tristate
rlabel metal2 s 12990 0 13046 800 6 slave_dat_o[2]
port 92 nsew signal tristate
rlabel metal2 s 28170 0 28226 800 6 slave_dat_o[30]
port 93 nsew signal tristate
rlabel metal2 s 28722 0 28778 800 6 slave_dat_o[31]
port 94 nsew signal tristate
rlabel metal2 s 13542 0 13598 800 6 slave_dat_o[3]
port 95 nsew signal tristate
rlabel metal2 s 14094 0 14150 800 6 slave_dat_o[4]
port 96 nsew signal tristate
rlabel metal2 s 14646 0 14702 800 6 slave_dat_o[5]
port 97 nsew signal tristate
rlabel metal2 s 15198 0 15254 800 6 slave_dat_o[6]
port 98 nsew signal tristate
rlabel metal2 s 15750 0 15806 800 6 slave_dat_o[7]
port 99 nsew signal tristate
rlabel metal2 s 16302 0 16358 800 6 slave_dat_o[8]
port 100 nsew signal tristate
rlabel metal2 s 16762 0 16818 800 6 slave_dat_o[9]
port 101 nsew signal tristate
rlabel metal2 s 2502 0 2558 800 6 slave_err_o
port 102 nsew signal tristate
rlabel metal2 s 2778 0 2834 800 6 slave_rty_o
port 103 nsew signal tristate
rlabel metal2 s 1122 0 1178 800 6 slave_sel_i[0]
port 104 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 slave_sel_i[1]
port 105 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 slave_sel_i[2]
port 106 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 slave_sel_i[3]
port 107 nsew signal input
rlabel metal2 s 846 0 902 800 6 slave_stb_i
port 108 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 slave_we_i
port 109 nsew signal input
rlabel metal3 s 28373 3816 29173 3936 6 spiMaster_miso
port 110 nsew signal input
rlabel metal3 s 28373 11568 29173 11688 6 spiMaster_mosi
port 111 nsew signal tristate
rlabel metal3 s 28373 19456 29173 19576 6 spiMaster_mosi_oe
port 112 nsew signal tristate
rlabel metal3 s 28373 27208 29173 27328 6 spiMaster_sclk
port 113 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 29173 31317
<< end >>
