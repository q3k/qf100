* NGSPICE file created from mkLanaiFrontend.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

.subckt mkLanaiFrontend CLK EN_core_dmem_request_put EN_core_dmem_response_get EN_core_imem_request_put
+ EN_core_imem_response_get EN_fmc_dmem_request_get EN_fmc_dmem_response_put EN_fmc_imem_request_get
+ EN_fmc_imem_response_put EN_ram_dmem_request_get EN_ram_dmem_response_put EN_ram_imem_request_get
+ EN_ram_imem_response_put RDY_core_dmem_request_put RDY_core_dmem_response_get RDY_core_imem_request_put
+ RDY_core_imem_response_get RDY_fmc_dmem_request_get RDY_fmc_dmem_response_put RDY_fmc_imem_request_get
+ RDY_fmc_imem_response_put RDY_ram_dmem_request_get RDY_ram_dmem_response_put RDY_ram_imem_request_get
+ RDY_ram_imem_response_put RST_N core_dmem_request_put[0] core_dmem_request_put[10]
+ core_dmem_request_put[11] core_dmem_request_put[12] core_dmem_request_put[13] core_dmem_request_put[14]
+ core_dmem_request_put[15] core_dmem_request_put[16] core_dmem_request_put[17] core_dmem_request_put[18]
+ core_dmem_request_put[19] core_dmem_request_put[1] core_dmem_request_put[20] core_dmem_request_put[21]
+ core_dmem_request_put[22] core_dmem_request_put[23] core_dmem_request_put[24] core_dmem_request_put[25]
+ core_dmem_request_put[26] core_dmem_request_put[27] core_dmem_request_put[28] core_dmem_request_put[29]
+ core_dmem_request_put[2] core_dmem_request_put[30] core_dmem_request_put[31] core_dmem_request_put[32]
+ core_dmem_request_put[33] core_dmem_request_put[34] core_dmem_request_put[35] core_dmem_request_put[36]
+ core_dmem_request_put[37] core_dmem_request_put[38] core_dmem_request_put[39] core_dmem_request_put[3]
+ core_dmem_request_put[40] core_dmem_request_put[41] core_dmem_request_put[42] core_dmem_request_put[43]
+ core_dmem_request_put[44] core_dmem_request_put[45] core_dmem_request_put[46] core_dmem_request_put[47]
+ core_dmem_request_put[48] core_dmem_request_put[49] core_dmem_request_put[4] core_dmem_request_put[50]
+ core_dmem_request_put[51] core_dmem_request_put[52] core_dmem_request_put[53] core_dmem_request_put[54]
+ core_dmem_request_put[55] core_dmem_request_put[56] core_dmem_request_put[57] core_dmem_request_put[58]
+ core_dmem_request_put[59] core_dmem_request_put[5] core_dmem_request_put[60] core_dmem_request_put[61]
+ core_dmem_request_put[62] core_dmem_request_put[63] core_dmem_request_put[64] core_dmem_request_put[65]
+ core_dmem_request_put[66] core_dmem_request_put[67] core_dmem_request_put[68] core_dmem_request_put[69]
+ core_dmem_request_put[6] core_dmem_request_put[70] core_dmem_request_put[71] core_dmem_request_put[72]
+ core_dmem_request_put[73] core_dmem_request_put[74] core_dmem_request_put[75] core_dmem_request_put[76]
+ core_dmem_request_put[77] core_dmem_request_put[78] core_dmem_request_put[79] core_dmem_request_put[7]
+ core_dmem_request_put[80] core_dmem_request_put[81] core_dmem_request_put[82] core_dmem_request_put[83]
+ core_dmem_request_put[84] core_dmem_request_put[85] core_dmem_request_put[86] core_dmem_request_put[87]
+ core_dmem_request_put[88] core_dmem_request_put[89] core_dmem_request_put[8] core_dmem_request_put[90]
+ core_dmem_request_put[91] core_dmem_request_put[92] core_dmem_request_put[93] core_dmem_request_put[94]
+ core_dmem_request_put[95] core_dmem_request_put[96] core_dmem_request_put[97] core_dmem_request_put[98]
+ core_dmem_request_put[99] core_dmem_request_put[9] core_dmem_response_get[0] core_dmem_response_get[10]
+ core_dmem_response_get[11] core_dmem_response_get[12] core_dmem_response_get[13]
+ core_dmem_response_get[14] core_dmem_response_get[15] core_dmem_response_get[16]
+ core_dmem_response_get[17] core_dmem_response_get[18] core_dmem_response_get[19]
+ core_dmem_response_get[1] core_dmem_response_get[20] core_dmem_response_get[21]
+ core_dmem_response_get[22] core_dmem_response_get[23] core_dmem_response_get[24]
+ core_dmem_response_get[25] core_dmem_response_get[26] core_dmem_response_get[27]
+ core_dmem_response_get[28] core_dmem_response_get[29] core_dmem_response_get[2]
+ core_dmem_response_get[30] core_dmem_response_get[31] core_dmem_response_get[3]
+ core_dmem_response_get[4] core_dmem_response_get[5] core_dmem_response_get[6] core_dmem_response_get[7]
+ core_dmem_response_get[8] core_dmem_response_get[9] core_imem_request_put[0] core_imem_request_put[10]
+ core_imem_request_put[11] core_imem_request_put[12] core_imem_request_put[13] core_imem_request_put[14]
+ core_imem_request_put[15] core_imem_request_put[16] core_imem_request_put[17] core_imem_request_put[18]
+ core_imem_request_put[19] core_imem_request_put[1] core_imem_request_put[20] core_imem_request_put[21]
+ core_imem_request_put[22] core_imem_request_put[23] core_imem_request_put[24] core_imem_request_put[25]
+ core_imem_request_put[26] core_imem_request_put[27] core_imem_request_put[28] core_imem_request_put[29]
+ core_imem_request_put[2] core_imem_request_put[30] core_imem_request_put[31] core_imem_request_put[3]
+ core_imem_request_put[4] core_imem_request_put[5] core_imem_request_put[6] core_imem_request_put[7]
+ core_imem_request_put[8] core_imem_request_put[9] core_imem_response_get[0] core_imem_response_get[10]
+ core_imem_response_get[11] core_imem_response_get[12] core_imem_response_get[13]
+ core_imem_response_get[14] core_imem_response_get[15] core_imem_response_get[16]
+ core_imem_response_get[17] core_imem_response_get[18] core_imem_response_get[19]
+ core_imem_response_get[1] core_imem_response_get[20] core_imem_response_get[21]
+ core_imem_response_get[22] core_imem_response_get[23] core_imem_response_get[24]
+ core_imem_response_get[25] core_imem_response_get[26] core_imem_response_get[27]
+ core_imem_response_get[28] core_imem_response_get[29] core_imem_response_get[2]
+ core_imem_response_get[30] core_imem_response_get[31] core_imem_response_get[3]
+ core_imem_response_get[4] core_imem_response_get[5] core_imem_response_get[6] core_imem_response_get[7]
+ core_imem_response_get[8] core_imem_response_get[9] fmc_dmem_request_get[0] fmc_dmem_request_get[10]
+ fmc_dmem_request_get[11] fmc_dmem_request_get[12] fmc_dmem_request_get[13] fmc_dmem_request_get[14]
+ fmc_dmem_request_get[15] fmc_dmem_request_get[16] fmc_dmem_request_get[17] fmc_dmem_request_get[18]
+ fmc_dmem_request_get[19] fmc_dmem_request_get[1] fmc_dmem_request_get[20] fmc_dmem_request_get[21]
+ fmc_dmem_request_get[22] fmc_dmem_request_get[23] fmc_dmem_request_get[24] fmc_dmem_request_get[25]
+ fmc_dmem_request_get[26] fmc_dmem_request_get[27] fmc_dmem_request_get[28] fmc_dmem_request_get[29]
+ fmc_dmem_request_get[2] fmc_dmem_request_get[30] fmc_dmem_request_get[31] fmc_dmem_request_get[32]
+ fmc_dmem_request_get[33] fmc_dmem_request_get[34] fmc_dmem_request_get[35] fmc_dmem_request_get[36]
+ fmc_dmem_request_get[37] fmc_dmem_request_get[38] fmc_dmem_request_get[39] fmc_dmem_request_get[3]
+ fmc_dmem_request_get[40] fmc_dmem_request_get[41] fmc_dmem_request_get[42] fmc_dmem_request_get[43]
+ fmc_dmem_request_get[44] fmc_dmem_request_get[45] fmc_dmem_request_get[46] fmc_dmem_request_get[47]
+ fmc_dmem_request_get[48] fmc_dmem_request_get[49] fmc_dmem_request_get[4] fmc_dmem_request_get[50]
+ fmc_dmem_request_get[51] fmc_dmem_request_get[52] fmc_dmem_request_get[53] fmc_dmem_request_get[54]
+ fmc_dmem_request_get[55] fmc_dmem_request_get[56] fmc_dmem_request_get[57] fmc_dmem_request_get[58]
+ fmc_dmem_request_get[59] fmc_dmem_request_get[5] fmc_dmem_request_get[60] fmc_dmem_request_get[61]
+ fmc_dmem_request_get[62] fmc_dmem_request_get[63] fmc_dmem_request_get[64] fmc_dmem_request_get[65]
+ fmc_dmem_request_get[66] fmc_dmem_request_get[67] fmc_dmem_request_get[68] fmc_dmem_request_get[69]
+ fmc_dmem_request_get[6] fmc_dmem_request_get[70] fmc_dmem_request_get[71] fmc_dmem_request_get[72]
+ fmc_dmem_request_get[73] fmc_dmem_request_get[74] fmc_dmem_request_get[75] fmc_dmem_request_get[76]
+ fmc_dmem_request_get[77] fmc_dmem_request_get[78] fmc_dmem_request_get[79] fmc_dmem_request_get[7]
+ fmc_dmem_request_get[80] fmc_dmem_request_get[81] fmc_dmem_request_get[82] fmc_dmem_request_get[83]
+ fmc_dmem_request_get[84] fmc_dmem_request_get[85] fmc_dmem_request_get[86] fmc_dmem_request_get[87]
+ fmc_dmem_request_get[88] fmc_dmem_request_get[89] fmc_dmem_request_get[8] fmc_dmem_request_get[90]
+ fmc_dmem_request_get[91] fmc_dmem_request_get[92] fmc_dmem_request_get[93] fmc_dmem_request_get[94]
+ fmc_dmem_request_get[95] fmc_dmem_request_get[96] fmc_dmem_request_get[97] fmc_dmem_request_get[98]
+ fmc_dmem_request_get[99] fmc_dmem_request_get[9] fmc_dmem_response_put[0] fmc_dmem_response_put[10]
+ fmc_dmem_response_put[11] fmc_dmem_response_put[12] fmc_dmem_response_put[13] fmc_dmem_response_put[14]
+ fmc_dmem_response_put[15] fmc_dmem_response_put[16] fmc_dmem_response_put[17] fmc_dmem_response_put[18]
+ fmc_dmem_response_put[19] fmc_dmem_response_put[1] fmc_dmem_response_put[20] fmc_dmem_response_put[21]
+ fmc_dmem_response_put[22] fmc_dmem_response_put[23] fmc_dmem_response_put[24] fmc_dmem_response_put[25]
+ fmc_dmem_response_put[26] fmc_dmem_response_put[27] fmc_dmem_response_put[28] fmc_dmem_response_put[29]
+ fmc_dmem_response_put[2] fmc_dmem_response_put[30] fmc_dmem_response_put[31] fmc_dmem_response_put[3]
+ fmc_dmem_response_put[4] fmc_dmem_response_put[5] fmc_dmem_response_put[6] fmc_dmem_response_put[7]
+ fmc_dmem_response_put[8] fmc_dmem_response_put[9] fmc_imem_request_get[0] fmc_imem_request_get[10]
+ fmc_imem_request_get[11] fmc_imem_request_get[12] fmc_imem_request_get[13] fmc_imem_request_get[14]
+ fmc_imem_request_get[15] fmc_imem_request_get[16] fmc_imem_request_get[17] fmc_imem_request_get[18]
+ fmc_imem_request_get[19] fmc_imem_request_get[1] fmc_imem_request_get[20] fmc_imem_request_get[21]
+ fmc_imem_request_get[22] fmc_imem_request_get[23] fmc_imem_request_get[24] fmc_imem_request_get[25]
+ fmc_imem_request_get[26] fmc_imem_request_get[27] fmc_imem_request_get[28] fmc_imem_request_get[29]
+ fmc_imem_request_get[2] fmc_imem_request_get[30] fmc_imem_request_get[31] fmc_imem_request_get[3]
+ fmc_imem_request_get[4] fmc_imem_request_get[5] fmc_imem_request_get[6] fmc_imem_request_get[7]
+ fmc_imem_request_get[8] fmc_imem_request_get[9] fmc_imem_response_put[0] fmc_imem_response_put[10]
+ fmc_imem_response_put[11] fmc_imem_response_put[12] fmc_imem_response_put[13] fmc_imem_response_put[14]
+ fmc_imem_response_put[15] fmc_imem_response_put[16] fmc_imem_response_put[17] fmc_imem_response_put[18]
+ fmc_imem_response_put[19] fmc_imem_response_put[1] fmc_imem_response_put[20] fmc_imem_response_put[21]
+ fmc_imem_response_put[22] fmc_imem_response_put[23] fmc_imem_response_put[24] fmc_imem_response_put[25]
+ fmc_imem_response_put[26] fmc_imem_response_put[27] fmc_imem_response_put[28] fmc_imem_response_put[29]
+ fmc_imem_response_put[2] fmc_imem_response_put[30] fmc_imem_response_put[31] fmc_imem_response_put[3]
+ fmc_imem_response_put[4] fmc_imem_response_put[5] fmc_imem_response_put[6] fmc_imem_response_put[7]
+ fmc_imem_response_put[8] fmc_imem_response_put[9] ram_dmem_request_get[0] ram_dmem_request_get[10]
+ ram_dmem_request_get[11] ram_dmem_request_get[12] ram_dmem_request_get[13] ram_dmem_request_get[14]
+ ram_dmem_request_get[15] ram_dmem_request_get[16] ram_dmem_request_get[17] ram_dmem_request_get[18]
+ ram_dmem_request_get[19] ram_dmem_request_get[1] ram_dmem_request_get[20] ram_dmem_request_get[21]
+ ram_dmem_request_get[22] ram_dmem_request_get[23] ram_dmem_request_get[24] ram_dmem_request_get[25]
+ ram_dmem_request_get[26] ram_dmem_request_get[27] ram_dmem_request_get[28] ram_dmem_request_get[29]
+ ram_dmem_request_get[2] ram_dmem_request_get[30] ram_dmem_request_get[31] ram_dmem_request_get[32]
+ ram_dmem_request_get[33] ram_dmem_request_get[34] ram_dmem_request_get[35] ram_dmem_request_get[36]
+ ram_dmem_request_get[37] ram_dmem_request_get[38] ram_dmem_request_get[39] ram_dmem_request_get[3]
+ ram_dmem_request_get[40] ram_dmem_request_get[41] ram_dmem_request_get[42] ram_dmem_request_get[43]
+ ram_dmem_request_get[44] ram_dmem_request_get[45] ram_dmem_request_get[46] ram_dmem_request_get[47]
+ ram_dmem_request_get[48] ram_dmem_request_get[49] ram_dmem_request_get[4] ram_dmem_request_get[50]
+ ram_dmem_request_get[51] ram_dmem_request_get[52] ram_dmem_request_get[53] ram_dmem_request_get[54]
+ ram_dmem_request_get[55] ram_dmem_request_get[56] ram_dmem_request_get[57] ram_dmem_request_get[58]
+ ram_dmem_request_get[59] ram_dmem_request_get[5] ram_dmem_request_get[60] ram_dmem_request_get[61]
+ ram_dmem_request_get[62] ram_dmem_request_get[63] ram_dmem_request_get[64] ram_dmem_request_get[65]
+ ram_dmem_request_get[66] ram_dmem_request_get[67] ram_dmem_request_get[68] ram_dmem_request_get[69]
+ ram_dmem_request_get[6] ram_dmem_request_get[70] ram_dmem_request_get[71] ram_dmem_request_get[72]
+ ram_dmem_request_get[73] ram_dmem_request_get[74] ram_dmem_request_get[75] ram_dmem_request_get[76]
+ ram_dmem_request_get[77] ram_dmem_request_get[78] ram_dmem_request_get[79] ram_dmem_request_get[7]
+ ram_dmem_request_get[80] ram_dmem_request_get[81] ram_dmem_request_get[82] ram_dmem_request_get[83]
+ ram_dmem_request_get[84] ram_dmem_request_get[85] ram_dmem_request_get[86] ram_dmem_request_get[87]
+ ram_dmem_request_get[88] ram_dmem_request_get[89] ram_dmem_request_get[8] ram_dmem_request_get[90]
+ ram_dmem_request_get[91] ram_dmem_request_get[92] ram_dmem_request_get[93] ram_dmem_request_get[94]
+ ram_dmem_request_get[95] ram_dmem_request_get[96] ram_dmem_request_get[97] ram_dmem_request_get[98]
+ ram_dmem_request_get[99] ram_dmem_request_get[9] ram_dmem_response_put[0] ram_dmem_response_put[10]
+ ram_dmem_response_put[11] ram_dmem_response_put[12] ram_dmem_response_put[13] ram_dmem_response_put[14]
+ ram_dmem_response_put[15] ram_dmem_response_put[16] ram_dmem_response_put[17] ram_dmem_response_put[18]
+ ram_dmem_response_put[19] ram_dmem_response_put[1] ram_dmem_response_put[20] ram_dmem_response_put[21]
+ ram_dmem_response_put[22] ram_dmem_response_put[23] ram_dmem_response_put[24] ram_dmem_response_put[25]
+ ram_dmem_response_put[26] ram_dmem_response_put[27] ram_dmem_response_put[28] ram_dmem_response_put[29]
+ ram_dmem_response_put[2] ram_dmem_response_put[30] ram_dmem_response_put[31] ram_dmem_response_put[3]
+ ram_dmem_response_put[4] ram_dmem_response_put[5] ram_dmem_response_put[6] ram_dmem_response_put[7]
+ ram_dmem_response_put[8] ram_dmem_response_put[9] ram_imem_request_get[0] ram_imem_request_get[10]
+ ram_imem_request_get[11] ram_imem_request_get[12] ram_imem_request_get[13] ram_imem_request_get[14]
+ ram_imem_request_get[15] ram_imem_request_get[16] ram_imem_request_get[17] ram_imem_request_get[18]
+ ram_imem_request_get[19] ram_imem_request_get[1] ram_imem_request_get[20] ram_imem_request_get[21]
+ ram_imem_request_get[22] ram_imem_request_get[23] ram_imem_request_get[24] ram_imem_request_get[25]
+ ram_imem_request_get[26] ram_imem_request_get[27] ram_imem_request_get[28] ram_imem_request_get[29]
+ ram_imem_request_get[2] ram_imem_request_get[30] ram_imem_request_get[31] ram_imem_request_get[3]
+ ram_imem_request_get[4] ram_imem_request_get[5] ram_imem_request_get[6] ram_imem_request_get[7]
+ ram_imem_request_get[8] ram_imem_request_get[9] ram_imem_response_put[0] ram_imem_response_put[10]
+ ram_imem_response_put[11] ram_imem_response_put[12] ram_imem_response_put[13] ram_imem_response_put[14]
+ ram_imem_response_put[15] ram_imem_response_put[16] ram_imem_response_put[17] ram_imem_response_put[18]
+ ram_imem_response_put[19] ram_imem_response_put[1] ram_imem_response_put[20] ram_imem_response_put[21]
+ ram_imem_response_put[22] ram_imem_response_put[23] ram_imem_response_put[24] ram_imem_response_put[25]
+ ram_imem_response_put[26] ram_imem_response_put[27] ram_imem_response_put[28] ram_imem_response_put[29]
+ ram_imem_response_put[2] ram_imem_response_put[30] ram_imem_response_put[31] ram_imem_response_put[3]
+ ram_imem_response_put[4] ram_imem_response_put[5] ram_imem_response_put[6] ram_imem_response_put[7]
+ ram_imem_response_put[8] ram_imem_response_put[9] vccd1 vssd1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3155_ _2462_/X _3155_/A2 _2587_/X _2588_/X _3130_/A vssd1 vssd1 vccd1 vccd1 _3489_/D
+ sky130_fd_sc_hd__a221o_1
X_3086_ _2077_/C _3077_/X _3081_/X _2399_/Y vssd1 vssd1 vccd1 vccd1 _3436_/D sky130_fd_sc_hd__o211ai_1
X_2106_ _2127_/A _2134_/B _2106_/C vssd1 vssd1 vccd1 vccd1 _2106_/Y sky130_fd_sc_hd__nand3_1
X_2037_ _3324_/Q _2020_/X _2036_/Y vssd1 vssd1 vccd1 vccd1 _2037_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1997__C _1997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2939_ _3341_/Q _2931_/X _2099_/Y vssd1 vssd1 vccd1 vccd1 _2940_/A sky130_fd_sc_hd__o21ai_1
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input127_A core_imem_request_put[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input92_A core_dmem_request_put[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_6_CLK clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3368_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_51_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2724_ _1541_/X _1534_/X _1562_/A _3223_/Q _2723_/X vssd1 vssd1 vccd1 vccd1 _3223_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_8_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput401 _2009_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[56] sky130_fd_sc_hd__buf_2
XFILLER_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2655_ _2655_/A _2655_/B vssd1 vssd1 vccd1 vccd1 _3178_/D sky130_fd_sc_hd__nand2_1
Xoutput434 _2118_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[86] sky130_fd_sc_hd__buf_2
Xoutput423 _2082_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[76] sky130_fd_sc_hd__buf_2
Xoutput412 _2045_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[66] sky130_fd_sc_hd__buf_2
X_1606_ _1606_/A vssd1 vssd1 vccd1 vccd1 _1606_/X sky130_fd_sc_hd__buf_4
Xoutput445 _2153_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[96] sky130_fd_sc_hd__buf_2
Xoutput467 _1517_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[25] sky130_fd_sc_hd__buf_2
X_2586_ _3154_/B vssd1 vssd1 vccd1 vccd1 _2586_/Y sky130_fd_sc_hd__inv_2
Xoutput478 _1448_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[6] sky130_fd_sc_hd__buf_2
Xoutput456 _1481_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[15] sky130_fd_sc_hd__buf_2
Xoutput489 _2229_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[16] sky130_fd_sc_hd__buf_2
XFILLER_59_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1537_ _1563_/A vssd1 vssd1 vccd1 vccd1 _1537_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1468_ _3172_/Q _1462_/X _1467_/Y vssd1 vssd1 vccd1 vccd1 _1468_/X sky130_fd_sc_hd__o21a_2
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3207_ _3225_/CLK _3207_/D vssd1 vssd1 vccd1 vccd1 _3207_/Q sky130_fd_sc_hd__dfxtp_1
X_3138_ _3127_/X _3138_/A2 _2530_/X _2531_/X _3128_/X vssd1 vssd1 vccd1 vccd1 _3475_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_27_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2872__B1 _2864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1801__B _1801_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3069_ _3423_/Q _3065_/X _2363_/Y _3061_/X vssd1 vssd1 vccd1 vccd1 _3423_/D sky130_fd_sc_hd__o211a_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1520__C _1520_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1529__A _1529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input244_A ram_imem_response_put[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2598__B_N _2473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output463_A _1504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2440_ _2156_/A _2159_/A _2162_/A _2131_/C _2434_/X vssd1 vssd1 vccd1 vccd1 _2440_/Y
+ sky130_fd_sc_hd__o311ai_4
XFILLER_5_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2371_ _2370_/X _2351_/X _3426_/Q vssd1 vssd1 vccd1 vccd1 _2371_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2707_ _2707_/A vssd1 vssd1 vccd1 vccd1 _2707_/X sky130_fd_sc_hd__clkbuf_2
X_2638_ _3170_/Q _2623_/X _1460_/Y vssd1 vssd1 vccd1 vccd1 _2640_/A sky130_fd_sc_hd__o21ai_1
Xoutput286 _2469_/Y vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[0] sky130_fd_sc_hd__buf_2
Xoutput275 _2616_/B vssd1 vssd1 vccd1 vccd1 RDY_core_dmem_response_get sky130_fd_sc_hd__buf_2
X_2569_ _2569_/A _2534_/X vssd1 vssd1 vccd1 vccd1 _2569_/X sky130_fd_sc_hd__or2b_1
Xoutput297 _2480_/X vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[1] sky130_fd_sc_hd__buf_2
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input194_A fmc_imem_response_put[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1584__B1 _1470_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2128__A2 _2111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input55_A core_dmem_request_put[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1940_ _2049_/A vssd1 vssd1 vccd1 vccd1 _1971_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_9_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1871_ _1871_/A vssd1 vssd1 vccd1 vccd1 _1871_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3472_ _3472_/CLK _3472_/D vssd1 vssd1 vccd1 vccd1 _3472_/Q sky130_fd_sc_hd__dfxtp_1
X_2423_ _2412_/X _2413_/X _2414_/X _2109_/C _2405_/X vssd1 vssd1 vccd1 vccd1 _2423_/Y
+ sky130_fd_sc_hd__o311ai_4
XFILLER_69_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2354_ _2973_/A vssd1 vssd1 vccd1 vccd1 _2459_/B sky130_fd_sc_hd__buf_2
XFILLER_69_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2285_ _2284_/X _2265_/X _3396_/Q vssd1 vssd1 vccd1 vccd1 _2285_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__1632__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2463__A _2605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input207_A fmc_imem_response_put[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output426_A _2092_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1452__A _1480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2070_ _3333_/Q _2056_/X _2069_/Y vssd1 vssd1 vccd1 vccd1 _2070_/X sky130_fd_sc_hd__o21a_2
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_11_CLK_A clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2283__A _2397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2972_ _3360_/Q _2145_/X _2797_/B vssd1 vssd1 vccd1 vccd1 _3360_/D sky130_fd_sc_hd__o21a_1
XFILLER_91_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1923_ _1923_/A vssd1 vssd1 vccd1 vccd1 _1924_/C sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_26_CLK_A clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1854_ _1869_/A _1877_/B _1854_/C vssd1 vssd1 vccd1 vccd1 _1854_/Y sky130_fd_sc_hd__nand3_1
X_1785_ input1/X vssd1 vssd1 vccd1 vccd1 _2163_/A sky130_fd_sc_hd__buf_4
X_3455_ _3457_/CLK _3455_/D vssd1 vssd1 vccd1 vccd1 _3455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2406_ _2384_/X _2385_/X _2386_/X _2088_/C _2405_/X vssd1 vssd1 vccd1 vccd1 _2406_/Y
+ sky130_fd_sc_hd__o311ai_4
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3386_ _3388_/CLK _3386_/D vssd1 vssd1 vccd1 vccd1 _3386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2337_ _1997_/C _2311_/X _2336_/Y vssd1 vssd1 vccd1 vccd1 _2337_/Y sky130_fd_sc_hd__o21ai_2
X_2268_ _2326_/A vssd1 vssd1 vccd1 vccd1 _2268_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2199_ _2176_/X _2178_/X _2180_/X _1821_/C _2152_/A vssd1 vssd1 vccd1 vccd1 _2199_/Y
+ sky130_fd_sc_hd__o311ai_4
XFILLER_25_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2736__C1 _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2751__A2 _2751_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input157_A fmc_dmem_response_put[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2503__A2 _2503_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2267__A1 _1909_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input18_A core_dmem_request_put[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output376_A _1925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1570_ _1563_/X _1569_/X _3201_/Q vssd1 vssd1 vccd1 vccd1 _1570_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2742__A2 _2742_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output543_A _2372_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _3258_/CLK _3240_/D vssd1 vssd1 vccd1 vccd1 _3240_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ _3482_/CLK _3171_/D vssd1 vssd1 vccd1 vccd1 _3171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2122_ _2206_/A vssd1 vssd1 vccd1 vccd1 _2152_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2053_ _2053_/A vssd1 vssd1 vccd1 vccd1 _2054_/C sky130_fd_sc_hd__inv_2
XFILLER_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2955_ _2955_/A _2965_/B vssd1 vssd1 vccd1 vccd1 _3349_/D sky130_fd_sc_hd__nand2_1
X_1906_ _1927_/A _1935_/B _1906_/C vssd1 vssd1 vccd1 vccd1 _1906_/Y sky130_fd_sc_hd__nand3_1
X_2886_ _3313_/Q _2873_/X _1997_/Y vssd1 vssd1 vccd1 vccd1 _2887_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__2981__A2 _2451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1837_ _3270_/Q _1834_/X _1836_/Y vssd1 vssd1 vccd1 vccd1 _1837_/X sky130_fd_sc_hd__o21a_1
X_1768_ _1637_/X _3257_/Q _1712_/A vssd1 vssd1 vccd1 vccd1 _1768_/X sky130_fd_sc_hd__o21ba_1
X_1699_ _2750_/B vssd1 vssd1 vccd1 vccd1 _1699_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3438_ _3440_/CLK _3438_/D vssd1 vssd1 vccd1 vccd1 _3438_/Q sky130_fd_sc_hd__dfxtp_1
X_3369_ _3461_/CLK _3369_/D vssd1 vssd1 vccd1 vccd1 _3369_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1523__C _1523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2972__A2 _2145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput120 core_imem_request_put[15] vssd1 vssd1 vccd1 vccd1 _1479_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_88_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput131 core_imem_request_put[25] vssd1 vssd1 vccd1 vccd1 _1515_/A sky130_fd_sc_hd__clkbuf_1
Xinput142 core_imem_request_put[6] vssd1 vssd1 vccd1 vccd1 _1446_/A sky130_fd_sc_hd__clkbuf_1
Xinput153 fmc_dmem_response_put[16] vssd1 vssd1 vccd1 vccd1 _2546_/A2 sky130_fd_sc_hd__buf_2
XFILLER_76_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput164 fmc_dmem_response_put[26] vssd1 vssd1 vccd1 vccd1 _2585_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput175 fmc_dmem_response_put[7] vssd1 vssd1 vccd1 vccd1 _3132_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput186 fmc_imem_response_put[17] vssd1 vssd1 vccd1 vccd1 _2755_/A2 sky130_fd_sc_hd__buf_2
Xinput197 fmc_imem_response_put[27] vssd1 vssd1 vccd1 vccd1 _2768_/A2 sky130_fd_sc_hd__buf_2
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2826__A _2864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2740_ _1772_/X _2740_/A2 _1665_/X _1666_/X _2771_/A vssd1 vssd1 vccd1 vccd1 _3232_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2963__A2 _2779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2671_ _3187_/Q _2660_/X _2661_/X _1520_/Y vssd1 vssd1 vccd1 vccd1 _3187_/D sky130_fd_sc_hd__o211a_1
X_1622_ _3220_/Q _1604_/X _1621_/Y vssd1 vssd1 vccd1 vccd1 _1622_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput605 _1628_/X vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[30] sky130_fd_sc_hd__buf_2
X_1553_ _1562_/A vssd1 vssd1 vccd1 vccd1 _1553_/X sky130_fd_sc_hd__clkbuf_2
X_1484_ _1512_/A _1484_/B _1484_/C vssd1 vssd1 vccd1 vccd1 _1484_/Y sky130_fd_sc_hd__nand3_1
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3223_ _3225_/CLK _3223_/D vssd1 vssd1 vccd1 vccd1 _3223_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3125__C1 _3154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3154_ _3154_/A _3154_/B vssd1 vssd1 vccd1 vccd1 _3488_/D sky130_fd_sc_hd__nor2_1
XFILLER_27_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3085_ _3435_/Q _3079_/X _2395_/Y _3075_/X vssd1 vssd1 vccd1 vccd1 _3435_/D sky130_fd_sc_hd__o211a_1
XFILLER_54_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2105_ _2105_/A vssd1 vssd1 vccd1 vccd1 _2106_/C sky130_fd_sc_hd__clkinv_2
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2036_ _2036_/A _2044_/B _2036_/C vssd1 vssd1 vccd1 vccd1 _2036_/Y sky130_fd_sc_hd__nand3_1
XFILLER_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2938_ _3340_/Q _2926_/X _2922_/X _2095_/Y vssd1 vssd1 vccd1 vccd1 _3340_/D sky130_fd_sc_hd__o211a_1
XFILLER_50_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2471__A _2520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2954__A2 _2950_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2869_ _3304_/Q _2868_/X _2864_/X _1963_/Y vssd1 vssd1 vccd1 vccd1 _3304_/D sky130_fd_sc_hd__o211a_1
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input85_A core_dmem_request_put[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output339_A _1767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output506_A _2275_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1460__A _1480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2723_ _2723_/A _2682_/B vssd1 vssd1 vccd1 vccd1 _2723_/X sky130_fd_sc_hd__or2b_1
Xoutput402 _2012_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[57] sky130_fd_sc_hd__buf_2
X_2654_ _3178_/Q _2644_/X _1488_/Y vssd1 vssd1 vccd1 vccd1 _2655_/A sky130_fd_sc_hd__o21ai_1
Xoutput435 _2121_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[87] sky130_fd_sc_hd__buf_2
Xoutput413 _2048_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[67] sky130_fd_sc_hd__buf_2
Xoutput424 _2085_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[77] sky130_fd_sc_hd__buf_2
X_1605_ _1605_/A vssd1 vssd1 vccd1 vccd1 _1605_/X sky130_fd_sc_hd__buf_4
X_2585_ _2520_/A _2585_/A2 _2583_/X _2584_/X vssd1 vssd1 vccd1 vccd1 _3154_/B sky130_fd_sc_hd__a22oi_4
Xoutput446 _2166_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[97] sky130_fd_sc_hd__buf_2
Xoutput468 _1521_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[26] sky130_fd_sc_hd__buf_2
X_1536_ _1591_/A vssd1 vssd1 vccd1 vccd1 _1563_/A sky130_fd_sc_hd__clkbuf_2
Xoutput457 _1485_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[16] sky130_fd_sc_hd__buf_2
Xoutput479 _1453_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[7] sky130_fd_sc_hd__buf_2
X_1467_ _1480_/A _1488_/B _1467_/C vssd1 vssd1 vccd1 vccd1 _1467_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__3113__A2 _2174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3206_ _3225_/CLK _3206_/D vssd1 vssd1 vccd1 vccd1 _3206_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2466__A _2605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3137_ _3139_/A _3137_/B vssd1 vssd1 vccd1 vccd1 _3474_/D sky130_fd_sc_hd__nor2_1
XFILLER_82_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1801__C _1801_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3068_ _2026_/C _3063_/X _3067_/X _2361_/Y vssd1 vssd1 vccd1 vccd1 _3422_/D sky130_fd_sc_hd__o211ai_1
XFILLER_23_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2019_ _3319_/Q _2002_/X _2018_/Y vssd1 vssd1 vccd1 vccd1 _2019_/X sky130_fd_sc_hd__o21a_2
XFILLER_23_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1545__A _1630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input237_A ram_dmem_response_put[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2615__A1 _2601_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_1_0_CLK_A clkbuf_2_1_0_CLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3040__A1 _1953_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output456_A _1481_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2370_ _2370_/A vssd1 vssd1 vccd1 vccd1 _2370_/X sky130_fd_sc_hd__buf_2
XFILLER_68_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2082__A2 _2075_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2706_ _3210_/Q _2695_/X _1595_/Y _2696_/X vssd1 vssd1 vccd1 vccd1 _3210_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1593__A1 _1480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2637_ _3169_/Q _2619_/X _2621_/X _1456_/Y vssd1 vssd1 vccd1 vccd1 _3169_/D sky130_fd_sc_hd__o211a_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput276 _1411_/Y vssd1 vssd1 vccd1 vccd1 RDY_core_imem_request_put sky130_fd_sc_hd__buf_2
X_2568_ _2542_/X _3484_/Q _2543_/X vssd1 vssd1 vccd1 vccd1 _2568_/X sky130_fd_sc_hd__o21ba_1
X_1519_ _1519_/A vssd1 vssd1 vccd1 vccd1 _1520_/C sky130_fd_sc_hd__inv_2
Xoutput287 _2519_/Y vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[10] sky130_fd_sc_hd__buf_2
Xoutput298 _2562_/Y vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[20] sky130_fd_sc_hd__buf_2
X_2499_ _2542_/A vssd1 vssd1 vccd1 vccd1 _2499_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_74_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2196__A _2225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2073__A2 _2056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3022__A1 _1909_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input187_A fmc_imem_response_put[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input48_A core_dmem_request_put[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3490__A _3490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1639__A2 _1639_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1870_ _3279_/Q _1852_/X _1869_/Y vssd1 vssd1 vccd1 vccd1 _1870_/X sky130_fd_sc_hd__o21a_2
XANTENNA_output573_A _2445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3013__A1 _1885_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1575__A1 _1460_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3471_ _3473_/CLK _3471_/D vssd1 vssd1 vccd1 vccd1 _3471_/Q sky130_fd_sc_hd__dfxtp_1
X_2422_ _2106_/C _2397_/X _2421_/Y vssd1 vssd1 vccd1 vccd1 _2422_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2353_ _2018_/C _2340_/X _2352_/Y vssd1 vssd1 vccd1 vccd1 _2353_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2284_ _2370_/A vssd1 vssd1 vccd1 vccd1 _2284_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2055__A2 _2038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1999_ _1999_/A vssd1 vssd1 vccd1 vccd1 _2000_/C sky130_fd_sc_hd__inv_2
XFILLER_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input102_A core_dmem_request_put[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1452__B _1452_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2971_ _2969_/A _3359_/Q _2959_/X vssd1 vssd1 vccd1 vccd1 _3359_/D sky130_fd_sc_hd__a21bo_1
XANTENNA__2037__A2 _2020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1922_ _2031_/A vssd1 vssd1 vccd1 vccd1 _1953_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_42_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1853_ _1853_/A vssd1 vssd1 vccd1 vccd1 _1854_/C sky130_fd_sc_hd__clkinv_4
X_1784_ _1871_/A vssd1 vssd1 vccd1 vccd1 _1784_/X sky130_fd_sc_hd__clkbuf_2
X_3454_ _3454_/CLK _3454_/D vssd1 vssd1 vccd1 vccd1 _3454_/Q sky130_fd_sc_hd__dfxtp_1
X_2405_ _2434_/A vssd1 vssd1 vccd1 vccd1 _2405_/X sky130_fd_sc_hd__buf_4
X_3385_ _3397_/CLK _3385_/D vssd1 vssd1 vccd1 vccd1 _3385_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1643__A _1776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2336_ _2312_/X _2323_/X _3414_/Q vssd1 vssd1 vccd1 vccd1 _2336_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_29_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2267_ _1909_/C _2253_/X _2266_/Y vssd1 vssd1 vccd1 vccd1 _2267_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2198_ _1815_/C _2195_/X _2197_/Y vssd1 vssd1 vccd1 vccd1 _2198_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2474__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2603__B_N _2464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2019__A2 _2002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1728__A _1728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output369_A _1902_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _3477_/CLK _3170_/D vssd1 vssd1 vccd1 vccd1 _3170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2121_ _3347_/Q _2111_/X _2120_/Y vssd1 vssd1 vccd1 vccd1 _2121_/X sky130_fd_sc_hd__o21a_2
X_2052_ _3328_/Q _2038_/X _2051_/Y vssd1 vssd1 vccd1 vccd1 _2052_/X sky130_fd_sc_hd__o21a_1
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2294__A _2351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2966__B1 _2959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2954_ _3349_/Q _2950_/X _2127_/Y vssd1 vssd1 vccd1 vccd1 _2955_/A sky130_fd_sc_hd__o21ai_1
X_2885_ _3312_/Q _2868_/X _2884_/X _1993_/Y vssd1 vssd1 vccd1 vccd1 _3312_/D sky130_fd_sc_hd__o211a_1
X_1905_ _1905_/A vssd1 vssd1 vccd1 vccd1 _1906_/C sky130_fd_sc_hd__clkinv_4
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1638__A _1638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1836_ _1850_/A _1859_/B _1836_/C vssd1 vssd1 vccd1 vccd1 _1836_/Y sky130_fd_sc_hd__nand3_2
X_1767_ _1734_/X _2770_/A2 _1765_/X _1766_/X vssd1 vssd1 vccd1 vccd1 _1767_/X sky130_fd_sc_hd__a22o_2
X_1698_ _1669_/X _1698_/A2 _1696_/X _1697_/X vssd1 vssd1 vccd1 vccd1 _2750_/B sky130_fd_sc_hd__a22oi_4
X_3437_ _3447_/CLK _3437_/D vssd1 vssd1 vccd1 vccd1 _3437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3368_ _3368_/CLK _3368_/D vssd1 vssd1 vccd1 vccd1 _3368_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1804__C _1804_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2319_ _2319_/A vssd1 vssd1 vccd1 vccd1 _2434_/A sky130_fd_sc_hd__clkbuf_2
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3299_ _3304_/CLK _3299_/D vssd1 vssd1 vccd1 vccd1 _3299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input267_A ram_imem_response_put[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_10_CLK_A clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput110 core_dmem_request_put[97] vssd1 vssd1 vccd1 vccd1 _1789_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__2488__A2 _3125_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput121 core_imem_request_put[16] vssd1 vssd1 vccd1 vccd1 _1483_/A sky130_fd_sc_hd__clkbuf_1
Xinput132 core_imem_request_put[26] vssd1 vssd1 vccd1 vccd1 _1519_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput143 core_imem_request_put[7] vssd1 vssd1 vccd1 vccd1 _1451_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input30_A core_dmem_request_put[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput154 fmc_dmem_response_put[17] vssd1 vssd1 vccd1 vccd1 _3145_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput165 fmc_dmem_response_put[27] vssd1 vssd1 vccd1 vccd1 _3155_/A2 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_25_CLK_A clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput176 fmc_dmem_response_put[8] vssd1 vssd1 vccd1 vccd1 _2510_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput187 fmc_imem_response_put[18] vssd1 vssd1 vccd1 vccd1 _1724_/A2 sky130_fd_sc_hd__buf_2
Xinput198 fmc_imem_response_put[28] vssd1 vssd1 vccd1 vccd1 _1763_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_91_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3003__A _3003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2670_ _2670_/A _2673_/B vssd1 vssd1 vccd1 vccd1 _3186_/D sky130_fd_sc_hd__nand2_1
X_1621_ _1605_/X _1606_/X _1607_/X _1520_/C _1443_/A vssd1 vssd1 vccd1 vccd1 _1621_/Y
+ sky130_fd_sc_hd__o311ai_4
Xoutput606 _1629_/X vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[31] sky130_fd_sc_hd__buf_2
X_1552_ _2707_/A vssd1 vssd1 vccd1 vccd1 _1562_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1483_ _1483_/A vssd1 vssd1 vccd1 vccd1 _1484_/C sky130_fd_sc_hd__inv_2
X_3222_ _3222_/CLK _3222_/D vssd1 vssd1 vccd1 vccd1 _3222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3153_ _2462_/X _3153_/A2 _2580_/X _2581_/X _3130_/A vssd1 vssd1 vccd1 vccd1 _3487_/D
+ sky130_fd_sc_hd__a221o_1
X_2104_ _2104_/A vssd1 vssd1 vccd1 vccd1 _2134_/B sky130_fd_sc_hd__clkbuf_2
X_3084_ _2069_/C _3077_/X _3081_/X _2393_/Y vssd1 vssd1 vccd1 vccd1 _3434_/D sky130_fd_sc_hd__o211ai_1
X_2035_ _2035_/A vssd1 vssd1 vccd1 vccd1 _2036_/C sky130_fd_sc_hd__clkinv_2
XFILLER_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2937_ _2937_/A _2952_/B vssd1 vssd1 vccd1 vccd1 _3339_/D sky130_fd_sc_hd__nand2_1
X_2868_ _2868_/A vssd1 vssd1 vccd1 vccd1 _2868_/X sky130_fd_sc_hd__buf_2
X_2799_ _3269_/Q _2795_/X _1832_/Y vssd1 vssd1 vccd1 vccd1 _2802_/A sky130_fd_sc_hd__o21ai_1
X_1819_ _2169_/A vssd1 vssd1 vccd1 vccd1 _1850_/A sky130_fd_sc_hd__buf_2
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input78_A core_dmem_request_put[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2722_ _3222_/Q _1630_/B _1625_/Y _2686_/X vssd1 vssd1 vccd1 vccd1 _3222_/D sky130_fd_sc_hd__o211a_1
X_2653_ _3177_/Q _2641_/X _2642_/X _1484_/Y vssd1 vssd1 vccd1 vccd1 _3177_/D sky130_fd_sc_hd__o211a_1
Xoutput425 _2089_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[78] sky130_fd_sc_hd__buf_2
Xoutput414 _2052_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[68] sky130_fd_sc_hd__buf_2
Xoutput403 _2016_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[58] sky130_fd_sc_hd__buf_2
X_1604_ _1630_/B vssd1 vssd1 vccd1 vccd1 _1604_/X sky130_fd_sc_hd__clkbuf_2
X_2584_ _2584_/A _2473_/A vssd1 vssd1 vccd1 vccd1 _2584_/X sky130_fd_sc_hd__or2b_1
Xoutput436 _2125_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[88] sky130_fd_sc_hd__buf_2
Xoutput447 _2167_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[98] sky130_fd_sc_hd__buf_2
Xoutput469 _1524_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[27] sky130_fd_sc_hd__buf_2
X_1535_ input3/X vssd1 vssd1 vccd1 vccd1 _1591_/A sky130_fd_sc_hd__inv_2
Xoutput458 _1489_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[17] sky130_fd_sc_hd__buf_2
X_1466_ _1466_/A vssd1 vssd1 vccd1 vccd1 _1467_/C sky130_fd_sc_hd__inv_2
XFILLER_79_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3205_ _3225_/CLK _3205_/D vssd1 vssd1 vccd1 vccd1 _3205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3136_ _3127_/X _3136_/A2 _2522_/X _2523_/X _3128_/X vssd1 vssd1 vccd1 vccd1 _3473_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2872__A2 _2868_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3067_ _3067_/A vssd1 vssd1 vccd1 vccd1 _3067_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2018_ _2018_/A _2026_/B _2018_/C vssd1 vssd1 vccd1 vccd1 _2018_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__2482__A _2482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input132_A core_imem_request_put[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2615__A2 _2615_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2705_ _1480_/C _2693_/X _2698_/X _1592_/Y vssd1 vssd1 vccd1 vccd1 _3209_/D sky130_fd_sc_hd__o211ai_1
XFILLER_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2636_ _2636_/A _2636_/B vssd1 vssd1 vccd1 vccd1 _3168_/D sky130_fd_sc_hd__nand2_1
X_2567_ _2563_/X _3149_/A2 _2565_/X _2566_/X vssd1 vssd1 vccd1 vccd1 _2567_/X sky130_fd_sc_hd__a22o_1
Xoutput277 _2773_/B vssd1 vssd1 vccd1 vccd1 RDY_core_imem_response_get sky130_fd_sc_hd__buf_2
XFILLER_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1518_ _2675_/A vssd1 vssd1 vccd1 vccd1 _1527_/A sky130_fd_sc_hd__clkbuf_4
Xoutput288 _2524_/X vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[11] sky130_fd_sc_hd__buf_2
Xoutput299 _2567_/X vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[21] sky130_fd_sc_hd__buf_2
X_2498_ _2541_/A vssd1 vssd1 vccd1 vccd1 _2498_/X sky130_fd_sc_hd__buf_4
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1449_ _1486_/A vssd1 vssd1 vccd1 vccd1 _2675_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2477__A _2605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3119_ _3116_/Y _3118_/Y _3114_/X vssd1 vssd1 vccd1 vccd1 _3459_/D sky130_fd_sc_hd__a21oi_1
XFILLER_70_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3470_ _3472_/CLK _3470_/D vssd1 vssd1 vccd1 vccd1 _3470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2421_ _2398_/X _2408_/X _3444_/Q vssd1 vssd1 vccd1 vccd1 _2421_/Y sky130_fd_sc_hd__o21ai_2
X_2352_ _2341_/X _2351_/X _3420_/Q vssd1 vssd1 vccd1 vccd1 _2352_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2283_ _2397_/A vssd1 vssd1 vccd1 vccd1 _2283_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2760__A _2760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1998_ _3313_/Q _1984_/X _1997_/Y vssd1 vssd1 vccd1 vccd1 _1998_/X sky130_fd_sc_hd__o21a_2
XFILLER_20_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2619_ _2660_/A vssd1 vssd1 vccd1 vccd1 _2619_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input60_A core_dmem_request_put[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1452__C _1452_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2845__A _2864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2970_ _2970_/A vssd1 vssd1 vccd1 vccd1 _3358_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1921_ _3292_/Q _1911_/X _1920_/Y vssd1 vssd1 vccd1 vccd1 _1921_/X sky130_fd_sc_hd__o21a_2
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_47_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3473_/CLK sky130_fd_sc_hd__clkbuf_16
X_1852_ _1871_/A vssd1 vssd1 vccd1 vccd1 _1852_/X sky130_fd_sc_hd__clkbuf_2
X_1783_ _2950_/A vssd1 vssd1 vccd1 vccd1 _1871_/A sky130_fd_sc_hd__clkbuf_2
X_3453_ _3457_/CLK _3453_/D vssd1 vssd1 vccd1 vccd1 _3453_/Q sky130_fd_sc_hd__dfxtp_1
X_2404_ _2084_/C _2397_/X _2403_/Y vssd1 vssd1 vccd1 vccd1 _2404_/Y sky130_fd_sc_hd__o21ai_4
X_3384_ _3384_/CLK _3384_/D vssd1 vssd1 vccd1 vccd1 _3384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2335_ _3413_/Q _2326_/X _2334_/Y vssd1 vssd1 vccd1 vccd1 _2335_/X sky130_fd_sc_hd__o21a_1
X_2266_ _2255_/X _2265_/X _3390_/Q vssd1 vssd1 vccd1 vccd1 _2266_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_29_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2197_ _2196_/X _2186_/X _3366_/Q vssd1 vssd1 vccd1 vccd1 _2197_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_80_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_38_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3489_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1711__A2 _2753_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input212_A ram_dmem_response_put[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3304_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1447__C _1447_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output431_A _2107_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2120_ _2127_/A _2134_/B _2120_/C vssd1 vssd1 vccd1 vccd1 _2120_/Y sky130_fd_sc_hd__nand3_1
XFILLER_94_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2051_ _2072_/A _2081_/B _2051_/C vssd1 vssd1 vccd1 vccd1 _2051_/Y sky130_fd_sc_hd__nand3_1
XFILLER_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2953_ _3348_/Q _2945_/X _2941_/X _2124_/Y vssd1 vssd1 vccd1 vccd1 _3348_/D sky130_fd_sc_hd__o211a_1
XFILLER_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1904_ _2049_/A vssd1 vssd1 vccd1 vccd1 _1935_/B sky130_fd_sc_hd__clkbuf_2
X_2884_ _2969_/B vssd1 vssd1 vccd1 vccd1 _2884_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1835_ _1835_/A vssd1 vssd1 vccd1 vccd1 _1836_/C sky130_fd_sc_hd__inv_4
X_1766_ _1766_/A _1635_/X vssd1 vssd1 vccd1 vccd1 _1766_/X sky130_fd_sc_hd__or2b_1
XFILLER_89_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1697_ _1697_/A _1661_/X vssd1 vssd1 vccd1 vccd1 _1697_/X sky130_fd_sc_hd__or2b_1
X_3436_ _3436_/CLK _3436_/D vssd1 vssd1 vccd1 vccd1 _3436_/Q sky130_fd_sc_hd__dfxtp_1
X_3367_ _3461_/CLK _3367_/D vssd1 vssd1 vccd1 vccd1 _3367_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ _1974_/C _2311_/X _2317_/Y vssd1 vssd1 vccd1 vccd1 _2318_/Y sky130_fd_sc_hd__o21ai_4
X_3298_ _3304_/CLK _3298_/D vssd1 vssd1 vccd1 vccd1 _3298_/Q sky130_fd_sc_hd__dfxtp_1
X_2249_ _2225_/X _2236_/X _3384_/Q vssd1 vssd1 vccd1 vccd1 _2249_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input162_A fmc_dmem_response_put[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput111 core_dmem_request_put[98] vssd1 vssd1 vccd1 vccd1 _1789_/B sky130_fd_sc_hd__clkbuf_2
Xinput100 core_dmem_request_put[88] vssd1 vssd1 vccd1 vccd1 _2123_/A sky130_fd_sc_hd__buf_2
XFILLER_76_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput144 core_imem_request_put[8] vssd1 vssd1 vccd1 vccd1 _1455_/A sky130_fd_sc_hd__clkbuf_1
Xinput133 core_imem_request_put[27] vssd1 vssd1 vccd1 vccd1 _1522_/A sky130_fd_sc_hd__clkbuf_1
Xinput122 core_imem_request_put[17] vssd1 vssd1 vccd1 vccd1 _1487_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput166 fmc_dmem_response_put[28] vssd1 vssd1 vccd1 vccd1 _2592_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput177 fmc_dmem_response_put[9] vssd1 vssd1 vccd1 vccd1 _3134_/A2 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input23_A core_dmem_request_put[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput155 fmc_dmem_response_put[18] vssd1 vssd1 vccd1 vccd1 _2553_/A2 sky130_fd_sc_hd__buf_2
XFILLER_91_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput199 fmc_imem_response_put[29] vssd1 vssd1 vccd1 vccd1 _2770_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput188 fmc_imem_response_put[19] vssd1 vssd1 vccd1 vccd1 _2759_/A2 sky130_fd_sc_hd__buf_2
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output381_A _1943_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1620__A1 _1516_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1620_ _1516_/C _1618_/X _1619_/Y vssd1 vssd1 vccd1 vccd1 _1620_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA_output479_A _1453_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput607 _1559_/Y vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[3] sky130_fd_sc_hd__buf_2
X_1551_ _1605_/A _1606_/A _1607_/A _1486_/A vssd1 vssd1 vccd1 vccd1 _2707_/A sky130_fd_sc_hd__o31ai_4
X_1482_ _1541_/A vssd1 vssd1 vccd1 vccd1 _1512_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_79_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3221_ _3221_/CLK _3221_/D vssd1 vssd1 vccd1 vccd1 _3221_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3125__A1 _2601_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_CLK clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3397_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3152_ _3152_/A _3152_/B vssd1 vssd1 vccd1 vccd1 _3486_/D sky130_fd_sc_hd__nor2_1
XFILLER_39_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2103_ _3342_/Q _2093_/X _2102_/Y vssd1 vssd1 vccd1 vccd1 _2103_/X sky130_fd_sc_hd__o21a_1
XFILLER_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3083_ _3433_/Q _3079_/X _2391_/Y _3075_/X vssd1 vssd1 vccd1 vccd1 _3433_/D sky130_fd_sc_hd__o211a_1
X_2034_ _3323_/Q _2020_/X _2033_/Y vssd1 vssd1 vccd1 vccd1 _2034_/X sky130_fd_sc_hd__o21a_2
XANTENNA__2100__A2 _2093_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2936_ _2936_/A vssd1 vssd1 vccd1 vccd1 _2952_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__1611__A1 _1503_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2867_ _2867_/A _2875_/B vssd1 vssd1 vccd1 vccd1 _3303_/D sky130_fd_sc_hd__nand2_1
X_1818_ _2097_/A vssd1 vssd1 vccd1 vccd1 _2169_/A sky130_fd_sc_hd__clkbuf_4
X_2798_ _3268_/Q _2789_/X _2784_/X _1829_/Y vssd1 vssd1 vccd1 vccd1 _3268_/D sky130_fd_sc_hd__o211a_1
X_1749_ _1712_/X _1749_/A2 _1747_/X _1748_/X vssd1 vssd1 vccd1 vccd1 _2765_/B sky130_fd_sc_hd__a22oi_4
XANTENNA__1815__C _1815_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3419_ _3431_/CLK _3419_/D vssd1 vssd1 vccd1 vccd1 _3419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1460__C _1460_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2721_ _1523_/C _1562_/A _2712_/X _1623_/Y vssd1 vssd1 vccd1 vccd1 _3221_/D sky130_fd_sc_hd__o211ai_1
XFILLER_8_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2652_ _2652_/A _2655_/B vssd1 vssd1 vccd1 vccd1 _3176_/D sky130_fd_sc_hd__nand2_1
Xoutput426 _2092_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[79] sky130_fd_sc_hd__buf_2
Xoutput415 _2055_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[69] sky130_fd_sc_hd__buf_2
Xoutput404 _2019_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[59] sky130_fd_sc_hd__buf_2
X_1603_ _1496_/C _1590_/X _1602_/Y vssd1 vssd1 vccd1 vccd1 _1603_/Y sky130_fd_sc_hd__o21ai_2
X_2583_ _2466_/X _3488_/Q _2541_/A vssd1 vssd1 vccd1 vccd1 _2583_/X sky130_fd_sc_hd__o21ba_1
Xoutput437 _2128_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[89] sky130_fd_sc_hd__buf_2
Xoutput448 _2168_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[99] sky130_fd_sc_hd__buf_2
X_1534_ _1607_/A vssd1 vssd1 vccd1 vccd1 _1534_/X sky130_fd_sc_hd__clkbuf_2
Xoutput459 _1493_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[18] sky130_fd_sc_hd__buf_2
XFILLER_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3204_ _3368_/CLK _3204_/D vssd1 vssd1 vccd1 vccd1 _3204_/Q sky130_fd_sc_hd__dfxtp_1
X_1465_ _3171_/Q _1462_/X _1464_/Y vssd1 vssd1 vccd1 vccd1 _1465_/X sky130_fd_sc_hd__o21a_2
X_3135_ _3139_/A _3135_/B vssd1 vssd1 vccd1 vccd1 _3472_/D sky130_fd_sc_hd__nor2_1
X_3066_ _3421_/Q _3065_/X _2359_/Y _3061_/X vssd1 vssd1 vccd1 vccd1 _3421_/D sky130_fd_sc_hd__o211a_1
X_2017_ _2017_/A vssd1 vssd1 vccd1 vccd1 _2018_/C sky130_fd_sc_hd__clkinv_2
XFILLER_35_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2919_ _3330_/Q _2907_/X _2903_/X _2058_/Y vssd1 vssd1 vccd1 vccd1 _3330_/D sky130_fd_sc_hd__o211a_1
XFILLER_10_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_24_CLK_A clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_39_CLK_A clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input125_A core_imem_request_put[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input90_A core_dmem_request_put[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1752__A _1752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2704_ _3208_/Q _2695_/X _1588_/Y _2696_/X vssd1 vssd1 vccd1 vccd1 _3208_/D sky130_fd_sc_hd__o211a_1
X_2635_ _3168_/Q _2623_/X _1452_/Y vssd1 vssd1 vccd1 vccd1 _2636_/A sky130_fd_sc_hd__o21ai_1
X_2566_ _2566_/A _2556_/X vssd1 vssd1 vccd1 vccd1 _2566_/X sky130_fd_sc_hd__or2b_1
X_1517_ _3186_/Q _1514_/X _1516_/Y vssd1 vssd1 vccd1 vccd1 _1517_/X sky130_fd_sc_hd__o21a_2
Xoutput278 _2170_/X vssd1 vssd1 vccd1 vccd1 RDY_fmc_dmem_request_get sky130_fd_sc_hd__buf_2
Xoutput289 _2528_/Y vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[12] sky130_fd_sc_hd__buf_2
X_2497_ input6/X vssd1 vssd1 vccd1 vccd1 _2541_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__1662__A _1662_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2758__A _2760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1448_ _3167_/Q _1441_/X _1447_/Y vssd1 vssd1 vccd1 vccd1 _1448_/X sky130_fd_sc_hd__o21a_2
XFILLER_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3118_ _2225_/A _2186_/X _3117_/Y vssd1 vssd1 vccd1 vccd1 _3118_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_82_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3049_ _3091_/A vssd1 vssd1 vccd1 vccd1 _3049_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input242_A ram_imem_response_put[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2221__A1 _1847_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2772__A2 _2772_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output461_A _1430_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2420_ _3443_/Q _2411_/X _2419_/Y vssd1 vssd1 vccd1 vccd1 _2420_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2351_ _2351_/A vssd1 vssd1 vccd1 vccd1 _2351_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2524__A2 _3136_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2282_ _3105_/A vssd1 vssd1 vccd1 vccd1 _2397_/A sky130_fd_sc_hd__buf_2
XANTENNA__1913__C _1913_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1997_ _2018_/A _2026_/B _1997_/C vssd1 vssd1 vccd1 vccd1 _1997_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__2971__B1_N _2959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2618_ _2618_/A vssd1 vssd1 vccd1 vccd1 _2660_/A sky130_fd_sc_hd__buf_2
X_2549_ _2549_/A _2513_/X vssd1 vssd1 vccd1 vccd1 _2549_/X sky130_fd_sc_hd__or2b_1
XANTENNA__2515__A2 _3134_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2279__A1 _1924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input192_A fmc_imem_response_put[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input53_A core_dmem_request_put[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1920_ _1927_/A _1935_/B _1920_/C vssd1 vssd1 vccd1 vccd1 _1920_/Y sky130_fd_sc_hd__nand3_1
X_1851_ _3274_/Q _1834_/X _1850_/Y vssd1 vssd1 vccd1 vccd1 _1851_/X sky130_fd_sc_hd__o21a_1
X_1782_ _2815_/A vssd1 vssd1 vccd1 vccd1 _2950_/A sky130_fd_sc_hd__buf_2
X_3452_ _3452_/CLK _3452_/D vssd1 vssd1 vccd1 vccd1 _3452_/Q sky130_fd_sc_hd__dfxtp_1
X_3383_ _3397_/CLK _3383_/D vssd1 vssd1 vccd1 vccd1 _3383_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3155__C1 _3130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2403_ _2398_/X _2380_/X _3438_/Q vssd1 vssd1 vccd1 vccd1 _2403_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__2101__A _2101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2334_ _2327_/X _2328_/X _2329_/X _1993_/C _2320_/X vssd1 vssd1 vccd1 vccd1 _2334_/Y
+ sky130_fd_sc_hd__o311ai_4
XFILLER_57_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2265_ _2351_/A vssd1 vssd1 vccd1 vccd1 _2265_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1940__A _2049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2196_ _2225_/A vssd1 vssd1 vccd1 vccd1 _2196_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2771__A _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2736__A2 _2736_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input205_A fmc_imem_response_put[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2681__A _2709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2727__A2 _1527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output424_A _2085_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2050_ _2050_/A vssd1 vssd1 vccd1 vccd1 _2051_/C sky130_fd_sc_hd__inv_2
XFILLER_81_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2591__A _2591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2952_ _2952_/A _2952_/B vssd1 vssd1 vccd1 vccd1 _3347_/D sky130_fd_sc_hd__nand2_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2966__A2 _2779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1903_ _2104_/A vssd1 vssd1 vccd1 vccd1 _2049_/A sky130_fd_sc_hd__buf_2
X_2883_ _2959_/A vssd1 vssd1 vccd1 vccd1 _2969_/B sky130_fd_sc_hd__clkbuf_2
X_1834_ _1871_/A vssd1 vssd1 vccd1 vccd1 _1834_/X sky130_fd_sc_hd__clkbuf_2
X_1765_ _1735_/X _3256_/Q _1743_/X vssd1 vssd1 vccd1 vccd1 _1765_/X sky130_fd_sc_hd__o21ba_1
X_3435_ _3449_/CLK _3435_/D vssd1 vssd1 vccd1 vccd1 _3435_/Q sky130_fd_sc_hd__dfxtp_1
X_1696_ _1670_/X _3239_/Q _1671_/X vssd1 vssd1 vccd1 vccd1 _1696_/X sky130_fd_sc_hd__o21ba_1
X_3366_ _3368_/CLK _3366_/D vssd1 vssd1 vccd1 vccd1 _3366_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ _2312_/X _2294_/X _3408_/Q vssd1 vssd1 vccd1 vccd1 _2317_/Y sky130_fd_sc_hd__o21ai_2
X_3297_ _3297_/CLK _3297_/D vssd1 vssd1 vccd1 vccd1 _3297_/Q sky130_fd_sc_hd__dfxtp_1
X_2248_ _3383_/Q _2239_/X _2247_/Y vssd1 vssd1 vccd1 vccd1 _2248_/X sky130_fd_sc_hd__o21a_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2179_ _2179_/A vssd1 vssd1 vccd1 vccd1 _2300_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2957__A2 _2950_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2006__A _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1845__A _2408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput101 core_dmem_request_put[89] vssd1 vssd1 vccd1 vccd1 _2126_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3134__A2 _3134_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input155_A fmc_dmem_response_put[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput123 core_imem_request_put[18] vssd1 vssd1 vccd1 vccd1 _1491_/A sky130_fd_sc_hd__clkbuf_1
Xinput134 core_imem_request_put[28] vssd1 vssd1 vccd1 vccd1 _1526_/A sky130_fd_sc_hd__clkbuf_1
Xinput112 core_dmem_request_put[99] vssd1 vssd1 vccd1 vccd1 _1789_/A sky130_fd_sc_hd__clkbuf_2
Xinput145 core_imem_request_put[9] vssd1 vssd1 vccd1 vccd1 _1459_/A sky130_fd_sc_hd__clkbuf_1
Xinput167 fmc_dmem_response_put[29] vssd1 vssd1 vccd1 vccd1 _2613_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput178 fmc_imem_response_put[0] vssd1 vssd1 vccd1 vccd1 _1639_/A2 sky130_fd_sc_hd__buf_4
Xinput156 fmc_dmem_response_put[19] vssd1 vssd1 vccd1 vccd1 _3147_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_63_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput189 fmc_imem_response_put[1] vssd1 vssd1 vccd1 vccd1 _2736_/A2 sky130_fd_sc_hd__buf_4
XANTENNA_input16_A core_dmem_request_put[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3070__A1 _2033_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output374_A _1918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput608 _1561_/X vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[4] sky130_fd_sc_hd__buf_2
X_1550_ _3194_/Q _1545_/X _1549_/Y vssd1 vssd1 vccd1 vccd1 _1550_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1755__A _1755_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1481_ _3176_/Q _1478_/X _1480_/Y vssd1 vssd1 vccd1 vccd1 _1481_/X sky130_fd_sc_hd__o21a_2
X_3220_ _3384_/CLK _3220_/D vssd1 vssd1 vccd1 vccd1 _3220_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3125__A2 _3125_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3151_ _3140_/X _3151_/A2 _2573_/X _2574_/X _3141_/X vssd1 vssd1 vccd1 vccd1 _3485_/D
+ sky130_fd_sc_hd__a221o_1
X_2102_ _2109_/A _2117_/B _2102_/C vssd1 vssd1 vccd1 vccd1 _2102_/Y sky130_fd_sc_hd__nand3_1
XFILLER_67_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1490__A _2675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3082_ _2062_/C _3077_/X _3081_/X _2389_/Y vssd1 vssd1 vccd1 vccd1 _3432_/D sky130_fd_sc_hd__o211ai_1
X_2033_ _2054_/A _2062_/B _2033_/C vssd1 vssd1 vccd1 vccd1 _2033_/Y sky130_fd_sc_hd__nand3_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2935_ _3339_/Q _2931_/X _2091_/Y vssd1 vssd1 vccd1 vccd1 _2937_/A sky130_fd_sc_hd__o21ai_1
X_2866_ _3303_/Q _2854_/X _1960_/Y vssd1 vssd1 vccd1 vccd1 _2867_/A sky130_fd_sc_hd__o21ai_1
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1817_ _2163_/A vssd1 vssd1 vccd1 vccd1 _2097_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2797_ _2797_/A _2797_/B vssd1 vssd1 vccd1 vccd1 _3267_/D sky130_fd_sc_hd__nand2_1
X_1748_ _1748_/A _1644_/A vssd1 vssd1 vccd1 vccd1 _1748_/X sky130_fd_sc_hd__or2b_1
X_1679_ _1670_/X _3235_/Q _1671_/X vssd1 vssd1 vccd1 vccd1 _1679_/X sky130_fd_sc_hd__o21ba_1
XFILLER_89_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3418_ _3420_/CLK _3418_/D vssd1 vssd1 vccd1 vccd1 _3418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3349_ _3452_/CLK _3349_/D vssd1 vssd1 vccd1 vccd1 _3349_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_input8_A EN_fmc_imem_response_put vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1678__A2 _2742_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input272_A ram_imem_response_put[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3107__A2 _2174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2315__B1 _1971_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2720_ _3220_/Q _2709_/X _1621_/Y _2710_/X vssd1 vssd1 vccd1 vccd1 _3220_/D sky130_fd_sc_hd__o211a_1
XFILLER_73_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2651_ _3176_/Q _2644_/X _1480_/Y vssd1 vssd1 vccd1 vccd1 _2652_/A sky130_fd_sc_hd__o21ai_1
X_1602_ _1591_/X _1597_/X _3213_/Q vssd1 vssd1 vccd1 vccd1 _1602_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2582_ _2563_/X _3153_/A2 _2580_/X _2581_/X vssd1 vssd1 vccd1 vccd1 _2582_/X sky130_fd_sc_hd__a22o_1
Xoutput416 _1822_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[6] sky130_fd_sc_hd__buf_2
Xoutput405 _1816_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[5] sky130_fd_sc_hd__buf_2
X_1533_ _1533_/A vssd1 vssd1 vccd1 vccd1 _1607_/A sky130_fd_sc_hd__buf_2
Xoutput427 _1825_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[7] sky130_fd_sc_hd__buf_2
Xoutput438 _1830_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[8] sky130_fd_sc_hd__buf_2
Xoutput449 _1833_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[9] sky130_fd_sc_hd__buf_2
X_1464_ _1476_/A _1484_/B _1464_/C vssd1 vssd1 vccd1 vccd1 _1464_/Y sky130_fd_sc_hd__nand3_1
X_3203_ _3225_/CLK _3203_/D vssd1 vssd1 vccd1 vccd1 _3203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3134_ _3127_/X _3134_/A2 _2512_/X _2514_/X _3128_/X vssd1 vssd1 vccd1 vccd1 _3471_/D
+ sky130_fd_sc_hd__a221o_1
X_3065_ _3093_/A vssd1 vssd1 vccd1 vccd1 _3065_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2016_ _3318_/Q _2002_/X _2015_/Y vssd1 vssd1 vccd1 vccd1 _2016_/X sky130_fd_sc_hd__o21a_1
XFILLER_70_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2085__A2 _2075_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2918_ _2918_/A _2933_/B vssd1 vssd1 vccd1 vccd1 _3329_/D sky130_fd_sc_hd__nand2_1
XFILLER_12_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2849_ _2868_/A vssd1 vssd1 vccd1 vccd1 _2849_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input118_A core_imem_request_put[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1587__A1 _1473_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input83_A core_dmem_request_put[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3025__A _3067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output337_A _1760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2864__A _2864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2703_ _1473_/C _2693_/X _2698_/X _1586_/Y vssd1 vssd1 vccd1 vccd1 _3207_/D sky130_fd_sc_hd__o211ai_1
X_2634_ _3167_/Q _2619_/X _2621_/X _1447_/Y vssd1 vssd1 vccd1 vccd1 _3167_/D sky130_fd_sc_hd__o211a_1
X_2565_ _2564_/X _3483_/Q _2529_/X vssd1 vssd1 vccd1 vccd1 _2565_/X sky130_fd_sc_hd__o21ba_1
X_1516_ _1516_/A _1523_/B _1516_/C vssd1 vssd1 vccd1 vccd1 _1516_/Y sky130_fd_sc_hd__nand3_1
XFILLER_87_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2496_ _2471_/X _3129_/A2 _2494_/X _2495_/X vssd1 vssd1 vccd1 vccd1 _2496_/X sky130_fd_sc_hd__a22o_1
Xoutput279 _3490_/A vssd1 vssd1 vccd1 vccd1 RDY_fmc_dmem_response_put sky130_fd_sc_hd__buf_2
XFILLER_59_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1447_ _1476_/A _1447_/B _1447_/C vssd1 vssd1 vccd1 vccd1 _1447_/Y sky130_fd_sc_hd__nand3_1
X_3117_ _3459_/Q vssd1 vssd1 vccd1 vccd1 _3117_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3048_ _3409_/Q _3037_/X _2321_/Y _3047_/X vssd1 vssd1 vccd1 vccd1 _3409_/D sky130_fd_sc_hd__o211a_1
XFILLER_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2014__A _2014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input235_A ram_dmem_response_put[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2859__A _2878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output454_A _1474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2350_ _3419_/Q _2326_/X _2349_/Y vssd1 vssd1 vccd1 vccd1 _2350_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2281_ _3395_/Q _2268_/X _2280_/Y vssd1 vssd1 vccd1 vccd1 _2281_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_23_CLK_A clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_38_CLK_A clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1996_ _1996_/A vssd1 vssd1 vccd1 vccd1 _1997_/C sky130_fd_sc_hd__inv_2
XFILLER_9_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2617_ _2617_/A vssd1 vssd1 vccd1 vccd1 _3160_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__1673__A _1673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2548_ _2521_/X _3479_/Q _2529_/X vssd1 vssd1 vccd1 vccd1 _2548_/X sky130_fd_sc_hd__o21ba_1
XFILLER_75_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2479_ _2479_/A _2478_/X vssd1 vssd1 vccd1 vccd1 _2479_/X sky130_fd_sc_hd__or2b_1
XFILLER_68_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1653__B_N _1637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input185_A fmc_imem_response_put[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input46_A core_dmem_request_put[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2442__A2 _1801_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1850_ _1850_/A _1859_/B _1850_/C vssd1 vssd1 vccd1 vccd1 _1850_/Y sky130_fd_sc_hd__nand3_2
X_1781_ _2175_/A _2177_/A _2179_/A input1/X vssd1 vssd1 vccd1 vccd1 _2815_/A sky130_fd_sc_hd__nor4b_2
X_3451_ _3457_/CLK _3451_/D vssd1 vssd1 vccd1 vccd1 _3451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2402_ _3437_/Q _2383_/X _2401_/Y vssd1 vssd1 vccd1 vccd1 _2402_/X sky130_fd_sc_hd__o21a_1
X_3382_ _3384_/CLK _3382_/D vssd1 vssd1 vccd1 vccd1 _3382_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1924__C _1924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2333_ _1990_/C _2311_/X _2332_/Y vssd1 vssd1 vccd1 vccd1 _2333_/Y sky130_fd_sc_hd__o21ai_4
X_2264_ _3389_/Q _2239_/X _2263_/Y vssd1 vssd1 vccd1 vccd1 _2264_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2195_ _2253_/A vssd1 vssd1 vccd1 vccd1 _2195_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2433__A2 _2426_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1668__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2771__B _2771_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1979_ _3308_/Q _1965_/X _1978_/Y vssd1 vssd1 vccd1 vccd1 _1979_/X sky130_fd_sc_hd__o21a_1
XFILLER_88_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2672__A2 _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input100_A core_dmem_request_put[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2188__A1 _1801_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2663__A2 _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2951_ _3347_/Q _2950_/X _2120_/Y vssd1 vssd1 vccd1 vccd1 _2952_/A sky130_fd_sc_hd__o21ai_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1902_ _3287_/Q _1892_/X _1901_/Y vssd1 vssd1 vccd1 vccd1 _1902_/X sky130_fd_sc_hd__o21a_2
X_2882_ _2882_/A _2895_/B vssd1 vssd1 vccd1 vccd1 _3311_/D sky130_fd_sc_hd__nand2_1
X_1833_ _3269_/Q _1813_/X _1832_/Y vssd1 vssd1 vccd1 vccd1 _1833_/X sky130_fd_sc_hd__o21a_1
X_1764_ _2769_/B vssd1 vssd1 vccd1 vccd1 _1764_/Y sky130_fd_sc_hd__inv_2
X_3434_ _3436_/CLK _3434_/D vssd1 vssd1 vccd1 vccd1 _3434_/Q sky130_fd_sc_hd__dfxtp_1
X_1695_ _1691_/X _2749_/A2 _1693_/X _1694_/X vssd1 vssd1 vccd1 vccd1 _1695_/X sky130_fd_sc_hd__a22o_1
XANTENNA__2112__A _2112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3365_ _3461_/CLK _3365_/D vssd1 vssd1 vccd1 vccd1 _3365_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1951__A _1951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2316_ _3407_/Q _2297_/X _2315_/Y vssd1 vssd1 vccd1 vccd1 _2316_/X sky130_fd_sc_hd__o21a_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _3304_/CLK _3296_/D vssd1 vssd1 vccd1 vccd1 _3296_/Q sky130_fd_sc_hd__dfxtp_1
X_2247_ _2240_/X _2241_/X _2242_/X _1880_/C _2232_/X vssd1 vssd1 vccd1 vccd1 _2247_/Y
+ sky130_fd_sc_hd__o311ai_4
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2178_ _2299_/A vssd1 vssd1 vccd1 vccd1 _2178_/X sky130_fd_sc_hd__buf_2
XFILLER_65_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1829__C _1829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2590__A1 _2466_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput102 core_dmem_request_put[8] vssd1 vssd1 vccd1 vccd1 _1828_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput113 core_dmem_request_put[9] vssd1 vssd1 vccd1 vccd1 _1831_/A sky130_fd_sc_hd__clkbuf_1
Xinput124 core_imem_request_put[19] vssd1 vssd1 vccd1 vccd1 _1495_/A sky130_fd_sc_hd__clkbuf_1
Xinput135 core_imem_request_put[29] vssd1 vssd1 vccd1 vccd1 _1533_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_input148_A fmc_dmem_response_put[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput168 fmc_dmem_response_put[2] vssd1 vssd1 vccd1 vccd1 _2483_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput157 fmc_dmem_response_put[1] vssd1 vssd1 vccd1 vccd1 _3123_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput146 fmc_dmem_response_put[0] vssd1 vssd1 vccd1 vccd1 _2468_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_91_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput179 fmc_imem_response_put[10] vssd1 vssd1 vccd1 vccd1 _1689_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput609 _1565_/Y vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[5] sky130_fd_sc_hd__buf_2
XANTENNA_output367_A _1895_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1480_ _1480_/A _1488_/B _1480_/C vssd1 vssd1 vccd1 vccd1 _1480_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__1771__A _2771_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2333__A1 _1990_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3150_ _3152_/A _3150_/B vssd1 vssd1 vccd1 vccd1 _3484_/D sky130_fd_sc_hd__nor2_1
X_2101_ _2101_/A vssd1 vssd1 vccd1 vccd1 _2102_/C sky130_fd_sc_hd__inv_2
X_3081_ _3095_/A vssd1 vssd1 vccd1 vccd1 _3081_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2032_ _2032_/A vssd1 vssd1 vccd1 vccd1 _2033_/C sky130_fd_sc_hd__inv_2
XFILLER_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1844__B1 _1843_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2934_ _3338_/Q _2926_/X _2922_/X _2088_/Y vssd1 vssd1 vccd1 vccd1 _3338_/D sky130_fd_sc_hd__o211a_1
XFILLER_15_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2865_ _3302_/Q _2849_/X _2864_/X _1956_/Y vssd1 vssd1 vccd1 vccd1 _3302_/D sky130_fd_sc_hd__o211a_1
X_1816_ _3265_/Q _1813_/X _1815_/Y vssd1 vssd1 vccd1 vccd1 _1816_/X sky130_fd_sc_hd__o21a_1
X_2796_ _3267_/Q _2795_/X _1824_/Y vssd1 vssd1 vccd1 vccd1 _2797_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__2167__A4 _2165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1747_ _1713_/X _3251_/Q _1714_/X vssd1 vssd1 vccd1 vccd1 _1747_/X sky130_fd_sc_hd__o21ba_1
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1678_ _1642_/X _2742_/A2 _1676_/X _1677_/X vssd1 vssd1 vccd1 vccd1 _1678_/X sky130_fd_sc_hd__a22o_1
X_3417_ _3457_/CLK _3417_/D vssd1 vssd1 vccd1 vccd1 _3417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2777__A _2936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3348_ _3356_/CLK _3348_/D vssd1 vssd1 vccd1 vccd1 _3348_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ _3288_/CLK _3279_/D vssd1 vssd1 vccd1 vccd1 _3279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2017__A _2017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1856__A _2319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input265_A ram_imem_response_put[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2251__B1 _1888_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2650_ _3175_/Q _2641_/X _2642_/X _1476_/Y vssd1 vssd1 vccd1 vccd1 _3175_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1766__A _1766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1601_ _3212_/Q _1576_/X _1600_/Y vssd1 vssd1 vccd1 vccd1 _1601_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput417 _2059_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[70] sky130_fd_sc_hd__buf_2
Xoutput406 _2023_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[60] sky130_fd_sc_hd__buf_2
X_2581_ _2581_/A _2556_/X vssd1 vssd1 vccd1 vccd1 _2581_/X sky130_fd_sc_hd__or2b_1
Xoutput428 _2096_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[80] sky130_fd_sc_hd__buf_2
Xoutput439 _2132_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[90] sky130_fd_sc_hd__buf_2
X_1532_ _1606_/A vssd1 vssd1 vccd1 vccd1 _2725_/B sky130_fd_sc_hd__clkbuf_2
X_1463_ _1463_/A vssd1 vssd1 vccd1 vccd1 _1464_/C sky130_fd_sc_hd__inv_2
XFILLER_79_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3202_ _3226_/CLK _3202_/D vssd1 vssd1 vccd1 vccd1 _3202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3133_ _3139_/A _3133_/B vssd1 vssd1 vccd1 vccd1 _3470_/D sky130_fd_sc_hd__nor2_1
XFILLER_27_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3064_ _2018_/C _3063_/X _3053_/X _2352_/Y vssd1 vssd1 vccd1 vccd1 _3420_/D sky130_fd_sc_hd__o211ai_1
XFILLER_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2015_ _2036_/A _2044_/B _2015_/C vssd1 vssd1 vccd1 vccd1 _2015_/Y sky130_fd_sc_hd__nand3_1
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2917_ _2936_/A vssd1 vssd1 vccd1 vccd1 _2933_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_2848_ _2848_/A _2856_/B vssd1 vssd1 vccd1 vccd1 _3293_/D sky130_fd_sc_hd__nand2_1
X_2779_ _2950_/A vssd1 vssd1 vccd1 vccd1 _2779_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_85_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2233__B1 _1866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input76_A core_dmem_request_put[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_10_CLK clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3384_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2702_ _3206_/Q _2695_/X _1584_/Y _2696_/X vssd1 vssd1 vccd1 vccd1 _3206_/D sky130_fd_sc_hd__o211a_1
XFILLER_13_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1927__C _1927_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2633_ _2633_/A _2636_/B vssd1 vssd1 vccd1 vccd1 _3166_/D sky130_fd_sc_hd__nand2_1
X_2564_ _2564_/A vssd1 vssd1 vccd1 vccd1 _2564_/X sky130_fd_sc_hd__clkbuf_2
X_1515_ _1515_/A vssd1 vssd1 vccd1 vccd1 _1516_/C sky130_fd_sc_hd__clkinv_4
X_2495_ _2495_/A _2478_/X vssd1 vssd1 vccd1 vccd1 _2495_/X sky130_fd_sc_hd__or2b_1
X_1446_ _1446_/A vssd1 vssd1 vccd1 vccd1 _1447_/C sky130_fd_sc_hd__inv_2
XFILLER_95_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3116_ _3116_/A _3116_/B vssd1 vssd1 vccd1 vccd1 _3116_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3047_ _3075_/A vssd1 vssd1 vccd1 vccd1 _3047_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3126__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1741__A2 _1741_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input130_A core_imem_request_put[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input228_A ram_dmem_response_put[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output447_A _2167_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2280_ _2269_/X _2270_/X _2271_/X _1927_/C _2262_/X vssd1 vssd1 vccd1 vccd1 _2280_/Y
+ sky130_fd_sc_hd__o311ai_4
XANTENNA__1732__A2 _1732_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2996__A1 _1840_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1995_ _2031_/A vssd1 vssd1 vccd1 vccd1 _2026_/B sky130_fd_sc_hd__clkbuf_2
X_2616_ _3130_/A _2616_/B vssd1 vssd1 vccd1 vccd1 _2617_/A sky130_fd_sc_hd__and2b_1
X_2547_ _3144_/B vssd1 vssd1 vccd1 vccd1 _2547_/Y sky130_fd_sc_hd__inv_2
X_2478_ _2564_/A vssd1 vssd1 vccd1 vccd1 _2478_/X sky130_fd_sc_hd__buf_2
X_1429_ _1443_/A _1452_/B _1429_/C vssd1 vssd1 vccd1 vccd1 _1429_/Y sky130_fd_sc_hd__nand3_1
XFILLER_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2987__A1 _1824_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1864__A _2967_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input178_A fmc_imem_response_put[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2695__A _2709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input39_A core_dmem_request_put[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2723__B_N _2682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1780_ _1789_/C vssd1 vssd1 vccd1 vccd1 _2179_/A sky130_fd_sc_hd__buf_4
XFILLER_6_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1774__A _1774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3450_ _3452_/CLK _3450_/D vssd1 vssd1 vccd1 vccd1 _3450_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3155__A1 _2462_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3381_ _3397_/CLK _3381_/D vssd1 vssd1 vccd1 vccd1 _3381_/Q sky130_fd_sc_hd__dfxtp_1
X_2401_ _2384_/X _2385_/X _2386_/X _2081_/C _2377_/X vssd1 vssd1 vccd1 vccd1 _2401_/Y
+ sky130_fd_sc_hd__o311ai_2
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2332_ _2312_/X _2323_/X _3412_/Q vssd1 vssd1 vccd1 vccd1 _2332_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2263_ _2240_/X _2241_/X _2242_/X _1906_/C _2262_/X vssd1 vssd1 vccd1 vccd1 _2263_/Y
+ sky130_fd_sc_hd__o311ai_2
X_2194_ _3365_/Q _2174_/X _2193_/Y vssd1 vssd1 vccd1 vccd1 _2194_/X sky130_fd_sc_hd__o21a_1
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2197__A2 _2186_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1978_ _2000_/A _2008_/B _1978_/C vssd1 vssd1 vccd1 vccd1 _1978_/Y sky130_fd_sc_hd__nand3_1
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2011__C _2011_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1850__C _1850_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2121__A2 _2111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2962__B _2965_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2188__A2 _2185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_22_CLK_A clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_37_CLK_A clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1769__A _1769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2950_ _2950_/A vssd1 vssd1 vccd1 vccd1 _2950_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2881_ _3311_/Q _2873_/X _1990_/Y vssd1 vssd1 vccd1 vccd1 _2882_/A sky130_fd_sc_hd__o21ai_1
X_1901_ _1909_/A _1917_/B _1901_/C vssd1 vssd1 vccd1 vccd1 _1901_/Y sky130_fd_sc_hd__nand3_1
XFILLER_30_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1832_ _1832_/A _1840_/B _1832_/C vssd1 vssd1 vccd1 vccd1 _1832_/Y sky130_fd_sc_hd__nand3_1
XFILLER_30_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1763_ _1691_/A _1763_/A2 _1761_/X _1762_/X vssd1 vssd1 vccd1 vccd1 _2769_/B sky130_fd_sc_hd__a22oi_4
XANTENNA__1935__C _1935_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1694_ _1694_/A _1684_/X vssd1 vssd1 vccd1 vccd1 _1694_/X sky130_fd_sc_hd__or2b_1
X_3433_ _3447_/CLK _3433_/D vssd1 vssd1 vccd1 vccd1 _3433_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _3368_/CLK _3364_/D vssd1 vssd1 vccd1 vccd1 _3364_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2315_ _2298_/X _2299_/X _2300_/X _1971_/C _2291_/X vssd1 vssd1 vccd1 vccd1 _2315_/Y
+ sky130_fd_sc_hd__o311ai_4
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _3297_/CLK _3295_/D vssd1 vssd1 vccd1 vccd1 _3295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2246_ _1877_/C _2224_/X _2245_/Y vssd1 vssd1 vccd1 vccd1 _2246_/Y sky130_fd_sc_hd__o21ai_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2103__A2 _2093_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2177_ _2177_/A vssd1 vssd1 vccd1 vccd1 _2299_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput103 core_dmem_request_put[90] vssd1 vssd1 vccd1 vccd1 _2130_/A sky130_fd_sc_hd__buf_2
Xinput125 core_imem_request_put[1] vssd1 vssd1 vccd1 vccd1 _1428_/A sky130_fd_sc_hd__clkbuf_1
Xinput136 core_imem_request_put[2] vssd1 vssd1 vccd1 vccd1 _1431_/A sky130_fd_sc_hd__clkbuf_1
Xinput114 core_imem_request_put[0] vssd1 vssd1 vccd1 vccd1 _1422_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput169 fmc_dmem_response_put[30] vssd1 vssd1 vccd1 vccd1 _2599_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput147 fmc_dmem_response_put[10] vssd1 vssd1 vccd1 vccd1 _2518_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput158 fmc_dmem_response_put[20] vssd1 vssd1 vccd1 vccd1 _2561_/A2 sky130_fd_sc_hd__buf_2
XFILLER_29_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input210_A ram_dmem_response_put[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2869__B1 _2864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3080_ _3431_/Q _3079_/X _2387_/Y _3075_/X vssd1 vssd1 vccd1 vccd1 _3431_/D sky130_fd_sc_hd__o211a_1
X_2100_ _3341_/Q _2093_/X _2099_/Y vssd1 vssd1 vccd1 vccd1 _2100_/X sky130_fd_sc_hd__o21a_2
XFILLER_94_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2031_ _2031_/A vssd1 vssd1 vccd1 vccd1 _2062_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__2883__A _2959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2933_ _2933_/A _2933_/B vssd1 vssd1 vccd1 vccd1 _3337_/D sky130_fd_sc_hd__nand2_1
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2864_ _2864_/A vssd1 vssd1 vccd1 vccd1 _2864_/X sky130_fd_sc_hd__buf_2
X_1815_ _1832_/A _1840_/B _1815_/C vssd1 vssd1 vccd1 vccd1 _1815_/Y sky130_fd_sc_hd__nand3_1
X_2795_ _2945_/A vssd1 vssd1 vccd1 vccd1 _2795_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2591__B_N _2473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2123__A _2123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1746_ _1734_/X _2764_/A2 _1744_/X _1745_/X vssd1 vssd1 vccd1 vccd1 _1746_/X sky130_fd_sc_hd__a22o_1
X_1677_ _1677_/A _1649_/X vssd1 vssd1 vccd1 vccd1 _1677_/X sky130_fd_sc_hd__or2b_1
X_3416_ _3420_/CLK _3416_/D vssd1 vssd1 vccd1 vccd1 _3416_/Q sky130_fd_sc_hd__dfxtp_1
X_3347_ _3448_/CLK _3347_/D vssd1 vssd1 vccd1 vccd1 _3347_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3278_ _3360_/CLK _3278_/D vssd1 vssd1 vccd1 vccd1 _3278_/Q sky130_fd_sc_hd__dfxtp_1
X_2229_ _3377_/Q _2210_/X _2228_/Y vssd1 vssd1 vccd1 vccd1 _2229_/X sky130_fd_sc_hd__o21a_1
XFILLER_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input258_A ram_imem_response_put[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input160_A fmc_dmem_response_put[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input21_A core_dmem_request_put[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3039__A _3067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1600_ _1577_/X _1578_/X _1579_/X _1492_/C _1594_/X vssd1 vssd1 vccd1 vccd1 _1600_/Y
+ sky130_fd_sc_hd__o311ai_4
XANTENNA_output477_A _1444_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput407 _2027_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[61] sky130_fd_sc_hd__buf_2
X_2580_ _2564_/X _3487_/Q _2572_/X vssd1 vssd1 vccd1 vccd1 _2580_/X sky130_fd_sc_hd__o21ba_1
Xoutput429 _2100_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[81] sky130_fd_sc_hd__buf_2
Xoutput418 _2063_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[71] sky130_fd_sc_hd__buf_2
X_1531_ _1531_/A vssd1 vssd1 vccd1 vccd1 _1606_/A sky130_fd_sc_hd__buf_2
XANTENNA__2878__A _2878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1462_ _1514_/A vssd1 vssd1 vccd1 vccd1 _1462_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3201_ _3226_/CLK _3201_/D vssd1 vssd1 vccd1 vccd1 _3201_/Q sky130_fd_sc_hd__dfxtp_1
X_3132_ _3127_/X _3132_/A2 _2505_/X _2506_/X _3128_/X vssd1 vssd1 vccd1 vccd1 _3469_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_94_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3063_ _3091_/A vssd1 vssd1 vccd1 vccd1 _3063_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2014_ _2014_/A vssd1 vssd1 vccd1 vccd1 _2015_/C sky130_fd_sc_hd__inv_2
XFILLER_23_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2916_ _3329_/Q _2912_/X _2054_/Y vssd1 vssd1 vccd1 vccd1 _2918_/A sky130_fd_sc_hd__o21ai_1
X_2847_ _3293_/Q _2835_/X _1924_/Y vssd1 vssd1 vccd1 vccd1 _2848_/A sky130_fd_sc_hd__o21ai_1
X_2778_ _3260_/Q _2145_/X _2965_/B _1794_/Y vssd1 vssd1 vccd1 vccd1 _3260_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2788__A _2794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1729_ _1691_/X _2759_/A2 _1726_/X _1728_/X vssd1 vssd1 vccd1 vccd1 _1729_/X sky130_fd_sc_hd__a22o_1
XANTENNA__2487__B_N _2478_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2028__A _2028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2481__A1 _2464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input69_A core_dmem_request_put[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2536__A2 _2536_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2701_ _1467_/C _2693_/X _2698_/X _1582_/Y vssd1 vssd1 vccd1 vccd1 _3205_/D sky130_fd_sc_hd__o211ai_1
XFILLER_13_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2632_ _3166_/Q _2623_/X _1443_/Y vssd1 vssd1 vccd1 vccd1 _2633_/A sky130_fd_sc_hd__o21ai_1
X_2563_ _3140_/A vssd1 vssd1 vccd1 vccd1 _2563_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2527__A2 _2527_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1514_ _1514_/A vssd1 vssd1 vccd1 vccd1 _1514_/X sky130_fd_sc_hd__buf_2
XFILLER_87_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2494_ _2473_/X _3467_/Q _2485_/X vssd1 vssd1 vccd1 vccd1 _2494_/X sky130_fd_sc_hd__o21ba_1
X_1445_ _1541_/A vssd1 vssd1 vccd1 vccd1 _1476_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3115_ _2169_/X _2162_/X _3105_/X _3458_/Q _3114_/X vssd1 vssd1 vccd1 vccd1 _3458_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3046_ _1974_/C _3035_/X _3039_/X _2317_/Y vssd1 vssd1 vccd1 vccd1 _3408_/D sky130_fd_sc_hd__o211ai_1
XFILLER_82_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2766__A2 _2766_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2518__A2 _2518_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2311__A _2397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2965__B _2965_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input123_A core_imem_request_put[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output342_A _1775_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output607_A _1559_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1994_ _3312_/Q _1984_/X _1993_/Y vssd1 vssd1 vccd1 vccd1 _1994_/X sky130_fd_sc_hd__o21a_1
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1938__C _1938_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2615_ _2601_/X _2615_/A2 _2602_/X _2603_/X _3154_/A vssd1 vssd1 vccd1 vccd1 _3159_/D
+ sky130_fd_sc_hd__a221o_1
X_2546_ _2541_/X _2546_/A2 _2544_/X _2545_/X vssd1 vssd1 vccd1 vccd1 _3144_/B sky130_fd_sc_hd__a22oi_4
XANTENNA__1970__A _1970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2477_ _2605_/B vssd1 vssd1 vccd1 vccd1 _2564_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1428_ _1428_/A vssd1 vssd1 vccd1 vccd1 _1429_/C sky130_fd_sc_hd__clkinv_4
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3029_ _3395_/Q _3023_/X _2280_/Y _3019_/X vssd1 vssd1 vccd1 vccd1 _3395_/D sky130_fd_sc_hd__o211a_1
XFILLER_83_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2987__A2 _2451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput590 _1599_/Y vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[17] sky130_fd_sc_hd__buf_2
XFILLER_78_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input240_A ram_dmem_response_put[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2400_ _2077_/C _2397_/X _2399_/Y vssd1 vssd1 vccd1 vccd1 _2400_/Y sky130_fd_sc_hd__o21ai_4
X_3380_ _3384_/CLK _3380_/D vssd1 vssd1 vccd1 vccd1 _3380_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3155__A2 _3155_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2331_ _3411_/Q _2326_/X _2330_/Y vssd1 vssd1 vccd1 vccd1 _2331_/X sky130_fd_sc_hd__o21a_1
X_2262_ _2291_/A vssd1 vssd1 vccd1 vccd1 _2262_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2193_ _2176_/X _2178_/X _2180_/X _1811_/C _2152_/A vssd1 vssd1 vccd1 vccd1 _2193_/Y
+ sky130_fd_sc_hd__o311ai_2
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2418__A1 _2099_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2126__A _2126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1977_ _1977_/A vssd1 vssd1 vccd1 vccd1 _1978_/C sky130_fd_sc_hd__inv_2
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2529_ _2572_/A vssd1 vssd1 vccd1 vccd1 _2529_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3082__A1 _2062_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1875__A _1951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input190_A fmc_imem_response_put[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input51_A core_dmem_request_put[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2880_ _3310_/Q _2868_/X _2864_/X _1986_/Y vssd1 vssd1 vccd1 vccd1 _3310_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1623__A2 _1452_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1900_ _1900_/A vssd1 vssd1 vccd1 vccd1 _1901_/C sky130_fd_sc_hd__clkinv_4
XFILLER_15_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1488__C _1488_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1831_ _1831_/A vssd1 vssd1 vccd1 vccd1 _1832_/C sky130_fd_sc_hd__inv_4
XFILLER_30_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1785__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1762_ _1762_/A _1644_/A vssd1 vssd1 vccd1 vccd1 _1762_/X sky130_fd_sc_hd__or2b_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1693_ _1692_/X _3238_/Q _1656_/X vssd1 vssd1 vccd1 vccd1 _1693_/X sky130_fd_sc_hd__o21ba_1
X_3432_ _3432_/CLK _3432_/D vssd1 vssd1 vccd1 vccd1 _3432_/Q sky130_fd_sc_hd__dfxtp_1
X_3363_ _3372_/CLK _3363_/D vssd1 vssd1 vccd1 vccd1 _3363_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2314_ _1967_/C _2311_/X _2313_/Y vssd1 vssd1 vccd1 vccd1 _2314_/Y sky130_fd_sc_hd__o21ai_4
X_3294_ _3304_/CLK _3294_/D vssd1 vssd1 vccd1 vccd1 _3294_/Q sky130_fd_sc_hd__dfxtp_1
X_2245_ _2225_/X _2236_/X _3382_/Q vssd1 vssd1 vccd1 vccd1 _2245_/Y sky130_fd_sc_hd__o21ai_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2176_ _2298_/A vssd1 vssd1 vccd1 vccd1 _2176_/X sky130_fd_sc_hd__buf_2
XFILLER_53_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput115 core_imem_request_put[10] vssd1 vssd1 vccd1 vccd1 _1463_/A sky130_fd_sc_hd__clkbuf_1
Xinput126 core_imem_request_put[20] vssd1 vssd1 vccd1 vccd1 _1499_/A sky130_fd_sc_hd__clkbuf_1
Xinput104 core_dmem_request_put[91] vssd1 vssd1 vccd1 vccd1 _2133_/A sky130_fd_sc_hd__clkbuf_2
Xinput137 core_imem_request_put[30] vssd1 vssd1 vccd1 vccd1 _1531_/A sky130_fd_sc_hd__clkbuf_4
Xinput148 fmc_dmem_response_put[11] vssd1 vssd1 vccd1 vccd1 _3136_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput159 fmc_dmem_response_put[21] vssd1 vssd1 vccd1 vccd1 _3149_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_56_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input203_A fmc_imem_response_put[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input99_A core_dmem_request_put[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2030__A2 _2020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output422_A _2078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2030_ _3322_/Q _2020_/X _2029_/Y vssd1 vssd1 vccd1 vccd1 _2030_/X sky130_fd_sc_hd__o21a_1
XFILLER_47_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3046__A1 _1974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2932_ _3337_/Q _2931_/X _2084_/Y vssd1 vssd1 vccd1 vccd1 _2933_/A sky130_fd_sc_hd__o21ai_1
XFILLER_30_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2863_ _2863_/A _2875_/B vssd1 vssd1 vccd1 vccd1 _3301_/D sky130_fd_sc_hd__nand2_1
X_1814_ _1814_/A vssd1 vssd1 vccd1 vccd1 _1815_/C sky130_fd_sc_hd__inv_4
X_2794_ _2794_/A vssd1 vssd1 vccd1 vccd1 _2945_/A sky130_fd_sc_hd__clkbuf_4
X_1745_ _1745_/A _1727_/X vssd1 vssd1 vccd1 vccd1 _1745_/X sky130_fd_sc_hd__or2b_1
XFILLER_7_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2309__B1 _1963_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1676_ _1644_/X _3234_/Q _1656_/X vssd1 vssd1 vccd1 vccd1 _1676_/X sky130_fd_sc_hd__o21ba_1
X_3415_ _3457_/CLK _3415_/D vssd1 vssd1 vccd1 vccd1 _3415_/Q sky130_fd_sc_hd__dfxtp_1
X_3346_ _3356_/CLK _3346_/D vssd1 vssd1 vccd1 vccd1 _3346_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ _3360_/CLK _3277_/D vssd1 vssd1 vccd1 vccd1 _3277_/Q sky130_fd_sc_hd__dfxtp_1
X_2228_ _2211_/X _2212_/X _2213_/X _1859_/C _2203_/X vssd1 vssd1 vccd1 vccd1 _2228_/Y
+ sky130_fd_sc_hd__o311ai_4
XANTENNA_clkbuf_leaf_21_CLK_A clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2159_ _2159_/A vssd1 vssd1 vccd1 vccd1 _3116_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1599__A1 _1488_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_36_CLK_A clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2012__A2 _2002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input153_A fmc_dmem_response_put[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input14_A core_dmem_request_put[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3028__A1 _1924_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput408 _2030_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[62] sky130_fd_sc_hd__buf_2
Xoutput419 _2066_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[72] sky130_fd_sc_hd__buf_2
X_1530_ _1605_/A vssd1 vssd1 vccd1 vccd1 _1530_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1461_ _3170_/Q _1441_/X _1460_/Y vssd1 vssd1 vccd1 vccd1 _1461_/X sky130_fd_sc_hd__o21a_2
X_3200_ _3226_/CLK _3200_/D vssd1 vssd1 vccd1 vccd1 _3200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3131_ _3139_/A _3131_/B vssd1 vssd1 vccd1 vccd1 _3468_/D sky130_fd_sc_hd__nor2_1
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3062_ _3419_/Q _3051_/X _2349_/Y _3061_/X vssd1 vssd1 vccd1 vccd1 _3419_/D sky130_fd_sc_hd__o211a_1
XFILLER_67_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2013_ _2049_/A vssd1 vssd1 vccd1 vccd1 _2044_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2778__B1 _2965_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2915_ _3328_/Q _2907_/X _2903_/X _2051_/Y vssd1 vssd1 vccd1 vccd1 _3328_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2134__A _2169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2846_ _3292_/Q _2830_/X _2845_/X _1920_/Y vssd1 vssd1 vccd1 vccd1 _3292_/D sky130_fd_sc_hd__o211a_1
X_2777_ _2936_/A vssd1 vssd1 vccd1 vccd1 _2965_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__1753__A1 _1734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1728_ _1728_/A _1727_/X vssd1 vssd1 vccd1 vccd1 _1728_/X sky130_fd_sc_hd__or2b_1
X_1659_ _1642_/X _2738_/A2 _1657_/X _1658_/X vssd1 vssd1 vccd1 vccd1 _1659_/X sky130_fd_sc_hd__a22o_1
XANTENNA_input6_A EN_fmc_dmem_response_put vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3329_ _3436_/CLK _3329_/D vssd1 vssd1 vccd1 vccd1 _3329_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input270_A ram_imem_response_put[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2700_ _3204_/Q _2695_/X _1580_/Y _2696_/X vssd1 vssd1 vccd1 vccd1 _3204_/D sky130_fd_sc_hd__o211a_1
XFILLER_9_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1496__C _1496_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2631_ _3165_/Q _2619_/X _2621_/X _1438_/Y vssd1 vssd1 vccd1 vccd1 _3165_/D sky130_fd_sc_hd__o211a_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2562_ _3148_/B vssd1 vssd1 vccd1 vccd1 _2562_/Y sky130_fd_sc_hd__inv_2
X_1513_ _3185_/Q _1498_/X _1512_/Y vssd1 vssd1 vccd1 vccd1 _1513_/X sky130_fd_sc_hd__o21a_2
X_2493_ _3126_/B vssd1 vssd1 vccd1 vccd1 _2493_/Y sky130_fd_sc_hd__inv_2
X_1444_ _3166_/Q _1441_/X _1443_/Y vssd1 vssd1 vccd1 vccd1 _1444_/X sky130_fd_sc_hd__o21a_2
XFILLER_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3114_ input9/X _2682_/B vssd1 vssd1 vccd1 vccd1 _3114_/X sky130_fd_sc_hd__or2b_1
X_3045_ _3407_/Q _3037_/X _2315_/Y _3033_/X vssd1 vssd1 vccd1 vccd1 _3407_/D sky130_fd_sc_hd__o211a_1
XFILLER_82_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2829_ _2829_/A _2837_/B vssd1 vssd1 vccd1 vccd1 _3283_/D sky130_fd_sc_hd__nand2_1
XFILLER_78_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input116_A core_imem_request_put[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input81_A core_dmem_request_put[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2502__A _2502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2390__A1 _2062_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output335_A _1753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2445__A2 _2439_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1993_ _2000_/A _2008_/B _1993_/C vssd1 vssd1 vccd1 vccd1 _1993_/Y sky130_fd_sc_hd__nand3_1
XFILLER_20_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2614_ _3126_/A _2614_/B vssd1 vssd1 vccd1 vccd1 _3158_/D sky130_fd_sc_hd__nor2_1
X_2545_ _2545_/A _2534_/X vssd1 vssd1 vccd1 vccd1 _2545_/X sky130_fd_sc_hd__or2b_1
XFILLER_87_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2476_ _2473_/X _3463_/Q _3140_/A vssd1 vssd1 vccd1 vccd1 _2476_/X sky130_fd_sc_hd__o21ba_1
XFILLER_87_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1427_ _1597_/A vssd1 vssd1 vccd1 vccd1 _1452_/B sky130_fd_sc_hd__buf_2
XFILLER_55_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3028_ _1924_/C _3021_/X _3025_/X _2278_/Y vssd1 vssd1 vccd1 vccd1 _3394_/D sky130_fd_sc_hd__o211ai_1
XFILLER_51_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2372__A1 _2040_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput580 _2458_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[99] sky130_fd_sc_hd__buf_2
Xoutput591 _1601_/X vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[18] sky130_fd_sc_hd__buf_2
XFILLER_78_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input233_A ram_dmem_response_put[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output452_A _1468_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2330_ _2327_/X _2328_/X _2329_/X _1986_/C _2320_/X vssd1 vssd1 vccd1 vccd1 _2330_/Y
+ sky130_fd_sc_hd__o311ai_2
X_2261_ _1901_/C _2253_/X _2260_/Y vssd1 vssd1 vccd1 vccd1 _2261_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__3063__A _3091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2192_ _1808_/C _2185_/X _2191_/Y vssd1 vssd1 vccd1 vccd1 _2192_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2666__A2 _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1949__C _1949_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1976_ _2049_/A vssd1 vssd1 vccd1 vccd1 _2008_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2142__A _2142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2528_ _3137_/B vssd1 vssd1 vccd1 vccd1 _2528_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2459_ _3461_/Q _2459_/B vssd1 vssd1 vccd1 vccd1 _2460_/A sky130_fd_sc_hd__or2_1
XFILLER_68_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1859__C _1859_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input183_A fmc_imem_response_put[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1891__A _2794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input44_A core_dmem_request_put[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1608__B1 _1500_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1830_ _3268_/Q _1813_/X _1829_/Y vssd1 vssd1 vccd1 vccd1 _1830_/X sky130_fd_sc_hd__o21a_1
XFILLER_30_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1761_ _1637_/X _3255_/Q _1712_/A vssd1 vssd1 vccd1 vccd1 _1761_/X sky130_fd_sc_hd__o21ba_1
X_1692_ _1735_/A vssd1 vssd1 vccd1 vccd1 _1692_/X sky130_fd_sc_hd__clkbuf_2
X_3431_ _3431_/CLK _3431_/D vssd1 vssd1 vccd1 vccd1 _3431_/Q sky130_fd_sc_hd__dfxtp_1
X_3362_ _3368_/CLK _3362_/D vssd1 vssd1 vccd1 vccd1 _3362_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ _2312_/X _2294_/X _3406_/Q vssd1 vssd1 vccd1 vccd1 _2313_/Y sky130_fd_sc_hd__o21ai_2
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _3297_/CLK _3293_/D vssd1 vssd1 vccd1 vccd1 _3293_/Q sky130_fd_sc_hd__dfxtp_1
X_2244_ _3381_/Q _2239_/X _2243_/Y vssd1 vssd1 vccd1 vccd1 _2244_/X sky130_fd_sc_hd__o21a_1
XFILLER_85_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2175_ _2175_/A vssd1 vssd1 vccd1 vccd1 _2298_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2272__B1 _1913_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1976__A _2049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1959_ _1959_/A vssd1 vssd1 vccd1 vccd1 _1960_/C sky130_fd_sc_hd__inv_2
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput116 core_imem_request_put[11] vssd1 vssd1 vccd1 vccd1 _1466_/A sky130_fd_sc_hd__clkbuf_1
Xinput127 core_imem_request_put[21] vssd1 vssd1 vccd1 vccd1 _1502_/A sky130_fd_sc_hd__clkbuf_1
Xinput105 core_dmem_request_put[92] vssd1 vssd1 vccd1 vccd1 _2136_/A sky130_fd_sc_hd__buf_2
XFILLER_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput138 core_imem_request_put[31] vssd1 vssd1 vccd1 vccd1 _1529_/A sky130_fd_sc_hd__clkbuf_4
Xinput149 fmc_dmem_response_put[12] vssd1 vssd1 vccd1 vccd1 _2527_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_29_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2263__B1 _1906_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2318__A1 _1974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_40_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3297_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2869__A2 _2868_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output415_A _2055_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2931_ _2950_/A vssd1 vssd1 vccd1 vccd1 _2931_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1796__A _2319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2862_ _3301_/Q _2854_/X _1953_/Y vssd1 vssd1 vccd1 vccd1 _2863_/A sky130_fd_sc_hd__o21ai_1
X_2793_ _3266_/Q _2789_/X _2784_/X _1821_/Y vssd1 vssd1 vccd1 vccd1 _3266_/D sky130_fd_sc_hd__o211a_1
X_1813_ _1871_/A vssd1 vssd1 vccd1 vccd1 _1813_/X sky130_fd_sc_hd__clkbuf_2
X_1744_ _1735_/X _3250_/Q _1743_/X vssd1 vssd1 vccd1 vccd1 _1744_/X sky130_fd_sc_hd__o21ba_1
X_3414_ _3456_/CLK _3414_/D vssd1 vssd1 vccd1 vccd1 _3414_/Q sky130_fd_sc_hd__dfxtp_1
X_1675_ _2741_/B vssd1 vssd1 vccd1 vccd1 _1675_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_31_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3448_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_58_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3345_ _3440_/CLK _3345_/D vssd1 vssd1 vccd1 vccd1 _3345_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ _3337_/CLK _3276_/D vssd1 vssd1 vccd1 vccd1 _3276_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ _1854_/C _2224_/X _2226_/Y vssd1 vssd1 vccd1 vccd1 _2227_/Y sky130_fd_sc_hd__o21ai_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2158_ _2413_/A vssd1 vssd1 vccd1 vccd1 _2159_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_26_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2089_ _3338_/Q _2075_/X _2088_/Y vssd1 vssd1 vccd1 vccd1 _2089_/X sky130_fd_sc_hd__o21a_1
XFILLER_26_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2033__C _2033_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3356_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_1_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2181__C1 _2152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input146_A fmc_dmem_response_put[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput409 _2034_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[63] sky130_fd_sc_hd__buf_2
XANTENNA_output365_A _1886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_CLK clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3404_/CLK sky130_fd_sc_hd__clkbuf_16
X_1460_ _1480_/A _1488_/B _1460_/C vssd1 vssd1 vccd1 vccd1 _1460_/Y sky130_fd_sc_hd__nand3_1
X_3130_ _3130_/A vssd1 vssd1 vccd1 vccd1 _3139_/A sky130_fd_sc_hd__clkbuf_2
X_3061_ _3075_/A vssd1 vssd1 vccd1 vccd1 _3061_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2012_ _3317_/Q _2002_/X _2011_/Y vssd1 vssd1 vccd1 vccd1 _2012_/X sky130_fd_sc_hd__o21a_2
XFILLER_90_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2914_ _2914_/A _2914_/B vssd1 vssd1 vccd1 vccd1 _3327_/D sky130_fd_sc_hd__nand2_1
X_2845_ _2864_/A vssd1 vssd1 vccd1 vccd1 _2845_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2776_ _2959_/A vssd1 vssd1 vccd1 vccd1 _2936_/A sky130_fd_sc_hd__buf_2
X_1727_ _1735_/A vssd1 vssd1 vccd1 vccd1 _1727_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1753__A2 _2766_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1658_ _1658_/A _1649_/X vssd1 vssd1 vccd1 vccd1 _1658_/X sky130_fd_sc_hd__or2b_1
X_1589_ _3208_/Q _1576_/X _1588_/Y vssd1 vssd1 vccd1 vccd1 _1589_/X sky130_fd_sc_hd__o21a_1
X_3328_ _3330_/CLK _3328_/D vssd1 vssd1 vccd1 vccd1 _3328_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3259_ _3259_/CLK _3259_/D vssd1 vssd1 vccd1 vccd1 _3259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2218__B1 _1843_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input263_A ram_imem_response_put[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2995__A _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2457__B1 _2185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_2_CLK clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3221_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2630_ _2630_/A _2636_/B vssd1 vssd1 vccd1 vccd1 _3164_/D sky130_fd_sc_hd__nand2_1
X_2561_ _2541_/X _2561_/A2 _2559_/X _2560_/X vssd1 vssd1 vccd1 vccd1 _3148_/B sky130_fd_sc_hd__a22oi_4
XANTENNA_clkbuf_leaf_20_CLK_A clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1512_ _1512_/A _1520_/B _1512_/C vssd1 vssd1 vccd1 vccd1 _1512_/Y sky130_fd_sc_hd__nand3_1
X_2492_ _2462_/X _2492_/A2 _2489_/X _2491_/X vssd1 vssd1 vccd1 vccd1 _3126_/B sky130_fd_sc_hd__a22oi_2
XFILLER_4_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1443_ _1443_/A _1452_/B _1443_/C vssd1 vssd1 vccd1 vccd1 _1443_/Y sky130_fd_sc_hd__nand3_1
XFILLER_4_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_35_CLK_A clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3113_ _3457_/Q _2174_/A _2454_/Y _3103_/X vssd1 vssd1 vccd1 vccd1 _3457_/D sky130_fd_sc_hd__o211a_1
XFILLER_67_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2448__B1 _2143_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3044_ _1967_/C _3035_/X _3039_/X _2313_/Y vssd1 vssd1 vccd1 vccd1 _3406_/D sky130_fd_sc_hd__o211ai_1
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2828_ _3283_/Q _2816_/X _1885_/Y vssd1 vssd1 vccd1 vccd1 _2829_/A sky130_fd_sc_hd__o21ai_1
X_2759_ _2757_/X _2759_/A2 _1726_/X _1728_/X _2758_/X vssd1 vssd1 vccd1 vccd1 _3246_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_2_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2687__B1 _2686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input109_A core_dmem_request_put[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input74_A core_dmem_request_put[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1717__A2 _1717_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output328_A _1729_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1992_ _1992_/A vssd1 vssd1 vccd1 vccd1 _1993_/C sky130_fd_sc_hd__inv_2
XFILLER_9_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2613_ _2601_/X _2613_/A2 _2594_/X _2595_/X _3154_/A vssd1 vssd1 vccd1 vccd1 _3157_/D
+ sky130_fd_sc_hd__a221o_1
X_2544_ _2542_/X _3478_/Q _2543_/X vssd1 vssd1 vccd1 vccd1 _2544_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__2131__C _2131_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2475_ _2572_/A vssd1 vssd1 vccd1 vccd1 _3140_/A sky130_fd_sc_hd__clkbuf_2
X_1426_ _1426_/A vssd1 vssd1 vccd1 vccd1 _1597_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3027_ _3393_/Q _3023_/X _2276_/Y _3019_/X vssd1 vssd1 vccd1 vccd1 _3393_/D sky130_fd_sc_hd__o211a_1
XFILLER_36_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2603__A _2603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput581 _2208_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[9] sky130_fd_sc_hd__buf_2
Xoutput570 _2205_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[8] sky130_fd_sc_hd__buf_2
XFILLER_78_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1580__B1 _1464_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput592 _1603_/Y vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[19] sky130_fd_sc_hd__buf_2
XANTENNA__1880__C _1880_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input226_A ram_dmem_response_put[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2260_ _2255_/X _2236_/X _3388_/Q vssd1 vssd1 vccd1 vccd1 _2260_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_69_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2191_ _2165_/X _2186_/X _3364_/Q vssd1 vssd1 vccd1 vccd1 _2191_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_65_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1799__A _2408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1975_ _3307_/Q _1965_/X _1974_/Y vssd1 vssd1 vccd1 vccd1 _1975_/X sky130_fd_sc_hd__o21a_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2527_ _2498_/X _2527_/A2 _2525_/X _2526_/X vssd1 vssd1 vccd1 vccd1 _3137_/B sky130_fd_sc_hd__a22oi_4
XFILLER_88_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2458_ _2169_/X _2156_/X _2185_/X _3460_/Q vssd1 vssd1 vccd1 vccd1 _2458_/X sky130_fd_sc_hd__a22o_2
XFILLER_75_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1409_ _3259_/Q vssd1 vssd1 vccd1 vccd1 _3491_/A sky130_fd_sc_hd__inv_6
XFILLER_68_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2389_ _2370_/X _2380_/X _3432_/Q vssd1 vssd1 vccd1 vccd1 _2389_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_83_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2290__A1 _1938_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input176_A fmc_dmem_response_put[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input37_A core_dmem_request_put[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2467__B_N _2466_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1412__A _3461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1760_ _1734_/X _2768_/A2 _1758_/X _1759_/X vssd1 vssd1 vccd1 vccd1 _1760_/X sky130_fd_sc_hd__a22o_2
X_1691_ _1691_/A vssd1 vssd1 vccd1 vccd1 _1691_/X sky130_fd_sc_hd__clkbuf_2
X_3430_ _3448_/CLK _3430_/D vssd1 vssd1 vccd1 vccd1 _3430_/Q sky130_fd_sc_hd__dfxtp_1
X_3361_ _3372_/CLK _3361_/D vssd1 vssd1 vccd1 vccd1 _3361_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2312_ _2370_/A vssd1 vssd1 vccd1 vccd1 _2312_/X sky130_fd_sc_hd__buf_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ _3432_/CLK _3292_/D vssd1 vssd1 vccd1 vccd1 _3292_/Q sky130_fd_sc_hd__dfxtp_1
X_2243_ _2240_/X _2241_/X _2242_/X _1873_/C _2232_/X vssd1 vssd1 vccd1 vccd1 _2243_/Y
+ sky130_fd_sc_hd__o311ai_4
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2174_ _2174_/A vssd1 vssd1 vccd1 vccd1 _2174_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2575__A2 _3151_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1958_ _2031_/A vssd1 vssd1 vccd1 vccd1 _1990_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__1992__A _1992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1889_ _3284_/Q _1871_/X _1888_/Y vssd1 vssd1 vccd1 vccd1 _1889_/X sky130_fd_sc_hd__o21a_2
XFILLER_88_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput117 core_imem_request_put[12] vssd1 vssd1 vccd1 vccd1 _1469_/A sky130_fd_sc_hd__clkbuf_1
Xinput106 core_dmem_request_put[93] vssd1 vssd1 vccd1 vccd1 _2139_/A sky130_fd_sc_hd__buf_2
XFILLER_88_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput139 core_imem_request_put[3] vssd1 vssd1 vccd1 vccd1 _1434_/A sky130_fd_sc_hd__clkbuf_1
Xinput128 core_imem_request_put[22] vssd1 vssd1 vccd1 vccd1 _1505_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2930_ _3336_/Q _2926_/X _2922_/X _2081_/Y vssd1 vssd1 vccd1 vccd1 _3336_/D sky130_fd_sc_hd__o211a_1
X_2861_ _3300_/Q _2849_/X _2845_/X _1949_/Y vssd1 vssd1 vccd1 vccd1 _3300_/D sky130_fd_sc_hd__o211a_1
X_1812_ _3264_/Q _1784_/X _1811_/Y vssd1 vssd1 vccd1 vccd1 _1812_/X sky130_fd_sc_hd__o21a_1
X_2792_ _2792_/A _2797_/B vssd1 vssd1 vccd1 vccd1 _3265_/D sky130_fd_sc_hd__nand2_1
X_1743_ _1743_/A vssd1 vssd1 vccd1 vccd1 _1743_/X sky130_fd_sc_hd__clkbuf_2
X_1674_ _1669_/X _1674_/A2 _1672_/X _1673_/X vssd1 vssd1 vccd1 vccd1 _2741_/B sky130_fd_sc_hd__a22oi_4
X_3413_ _3413_/CLK _3413_/D vssd1 vssd1 vccd1 vccd1 _3413_/Q sky130_fd_sc_hd__dfxtp_1
X_3344_ _3356_/CLK _3344_/D vssd1 vssd1 vccd1 vccd1 _3344_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _3360_/CLK _3275_/D vssd1 vssd1 vccd1 vccd1 _3275_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ _2225_/X _2206_/X _3376_/Q vssd1 vssd1 vccd1 vccd1 _2226_/Y sky130_fd_sc_hd__o21ai_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2157_ _2177_/A vssd1 vssd1 vccd1 vccd1 _2413_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2088_ _2109_/A _2117_/B _2088_/C vssd1 vssd1 vccd1 vccd1 _2088_/Y sky130_fd_sc_hd__nand3_1
XFILLER_41_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2611__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2181__B1 _1794_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input139_A core_imem_request_put[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output358_A _1863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output525_A _2325_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3060_ _2011_/C _3049_/X _3053_/X _2346_/Y vssd1 vssd1 vccd1 vccd1 _3418_/D sky130_fd_sc_hd__o211ai_1
XFILLER_94_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2011_ _2018_/A _2026_/B _2011_/C vssd1 vssd1 vccd1 vccd1 _2011_/Y sky130_fd_sc_hd__nand3_1
XFILLER_63_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2227__A1 _1854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2778__A2 _2145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2913_ _3327_/Q _2912_/X _2047_/Y vssd1 vssd1 vccd1 vccd1 _2914_/A sky130_fd_sc_hd__o21ai_1
X_2844_ _2844_/A _2856_/B vssd1 vssd1 vccd1 vccd1 _3291_/D sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_9_CLK_A clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2775_ input5/X _2975_/B vssd1 vssd1 vccd1 vccd1 _2959_/A sky130_fd_sc_hd__nor2b_2
X_1726_ _1692_/X _3246_/Q _1700_/X vssd1 vssd1 vccd1 vccd1 _1726_/X sky130_fd_sc_hd__o21ba_1
X_1657_ _1644_/X _3230_/Q _1656_/X vssd1 vssd1 vccd1 vccd1 _1657_/X sky130_fd_sc_hd__o21ba_1
X_1588_ _1577_/X _1578_/X _1579_/X _1476_/C _1566_/X vssd1 vssd1 vccd1 vccd1 _1588_/Y
+ sky130_fd_sc_hd__o311ai_4
X_3327_ _3436_/CLK _3327_/D vssd1 vssd1 vccd1 vccd1 _3327_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3258_ _3258_/CLK _3258_/D vssd1 vssd1 vccd1 vccd1 _3258_/Q sky130_fd_sc_hd__dfxtp_1
X_2209_ _2973_/A vssd1 vssd1 vccd1 vccd1 _2326_/A sky130_fd_sc_hd__clkbuf_2
X_3189_ _3388_/CLK _3189_/D vssd1 vssd1 vccd1 vccd1 _3189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2341__A _2370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input256_A ram_imem_response_put[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2457__A1 _2169_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output475_A _1436_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2560_ _2560_/A _2534_/X vssd1 vssd1 vccd1 vccd1 _2560_/X sky130_fd_sc_hd__or2b_1
X_1511_ _1511_/A vssd1 vssd1 vccd1 vccd1 _1512_/C sky130_fd_sc_hd__inv_2
X_2491_ _2491_/A _2490_/X vssd1 vssd1 vccd1 vccd1 _2491_/X sky130_fd_sc_hd__or2b_1
XFILLER_4_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1442_ _1442_/A vssd1 vssd1 vccd1 vccd1 _1443_/C sky130_fd_sc_hd__clkinv_4
XFILLER_67_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3112_ _2147_/C _3105_/X _3003_/A _2452_/Y vssd1 vssd1 vccd1 vccd1 _3456_/D sky130_fd_sc_hd__o211ai_1
X_3043_ _3405_/Q _3037_/X _2309_/Y _3033_/X vssd1 vssd1 vccd1 vccd1 _3405_/D sky130_fd_sc_hd__o211a_1
XFILLER_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2426__A _3035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2827_ _3282_/Q _2810_/X _2826_/X _1880_/Y vssd1 vssd1 vccd1 vccd1 _3282_/D sky130_fd_sc_hd__o211a_1
X_2758_ _2760_/A vssd1 vssd1 vccd1 vccd1 _2758_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1709_ _1692_/X _3242_/Q _1700_/X vssd1 vssd1 vccd1 vccd1 _1709_/X sky130_fd_sc_hd__o21ba_1
X_2689_ _1435_/C _1618_/X _2686_/X _1558_/Y vssd1 vssd1 vccd1 vccd1 _3197_/D sky130_fd_sc_hd__o211ai_1
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2687__A1 _1429_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2975__A_N input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2071__A _2071_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input67_A core_dmem_request_put[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1415__A _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1991_ _3311_/Q _1984_/X _1990_/Y vssd1 vssd1 vccd1 vccd1 _1991_/X sky130_fd_sc_hd__o21a_2
XFILLER_20_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2602__A1 _2478_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3077__A _3091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2612_ _3143_/A vssd1 vssd1 vccd1 vccd1 _3154_/A sky130_fd_sc_hd__clkbuf_4
X_2543_ input6/X vssd1 vssd1 vccd1 vccd1 _2543_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2474_ input6/X vssd1 vssd1 vccd1 vccd1 _2572_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1425_ _1486_/A vssd1 vssd1 vccd1 vccd1 _1443_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3026_ _1917_/C _3021_/X _3025_/X _2274_/Y vssd1 vssd1 vccd1 vccd1 _3392_/D sky130_fd_sc_hd__o211ai_1
XFILLER_36_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3149__A2 _3149_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput560 _2416_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[80] sky130_fd_sc_hd__buf_2
Xoutput571 _2441_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[90] sky130_fd_sc_hd__buf_2
Xoutput582 _1550_/X vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[0] sky130_fd_sc_hd__buf_2
Xoutput593 _1555_/Y vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[1] sky130_fd_sc_hd__buf_2
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1744__B1_N _1743_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input219_A ram_dmem_response_put[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input121_A core_imem_request_put[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_34_CLK_A clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1571__A1 _1452_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_49_CLK_A clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2190_ _3363_/Q _2174_/X _2189_/Y vssd1 vssd1 vccd1 vccd1 _2190_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output605_A _1628_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1974_ _1981_/A _1990_/B _1974_/C vssd1 vssd1 vccd1 vccd1 _1974_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__3000__A1 _1854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2526_ _2526_/A _2490_/X vssd1 vssd1 vccd1 vccd1 _2526_/X sky130_fd_sc_hd__or2b_1
XANTENNA__1981__C _1981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2457_ _2169_/X _3116_/B _2185_/X _3459_/Q vssd1 vssd1 vccd1 vccd1 _2457_/X sky130_fd_sc_hd__a22o_2
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2388_ _3431_/Q _2383_/X _2387_/Y vssd1 vssd1 vccd1 vccd1 _2388_/X sky130_fd_sc_hd__o21a_1
XFILLER_56_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3009_ _3009_/A vssd1 vssd1 vccd1 vccd1 _3067_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2614__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input169_A fmc_dmem_response_put[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput390 _1972_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[46] sky130_fd_sc_hd__buf_2
XFILLER_74_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3058__A1 _2004_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1412__B _3360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output388_A _1964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1690_ _2748_/B vssd1 vssd1 vccd1 vccd1 _1690_/Y sky130_fd_sc_hd__inv_2
X_3360_ _3360_/CLK _3360_/D vssd1 vssd1 vccd1 vccd1 _3360_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2311_ _2397_/A vssd1 vssd1 vccd1 vccd1 _2311_/X sky130_fd_sc_hd__clkbuf_4
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _3486_/CLK _3291_/D vssd1 vssd1 vccd1 vccd1 _3291_/Q sky130_fd_sc_hd__dfxtp_1
X_2242_ _2300_/A vssd1 vssd1 vccd1 vccd1 _2242_/X sky130_fd_sc_hd__buf_2
XFILLER_78_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2173_ _3093_/A vssd1 vssd1 vccd1 vccd1 _2174_/A sky130_fd_sc_hd__buf_2
XANTENNA__2137__C _2137_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1957_ _3302_/Q _1947_/X _1956_/Y vssd1 vssd1 vccd1 vccd1 _1957_/X sky130_fd_sc_hd__o21a_2
X_1888_ _1888_/A _1898_/B _1888_/C vssd1 vssd1 vccd1 vccd1 _1888_/Y sky130_fd_sc_hd__nand3_1
XFILLER_88_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2509_ _2509_/A _2490_/X vssd1 vssd1 vccd1 vccd1 _2509_/X sky130_fd_sc_hd__or2b_1
XFILLER_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput118 core_imem_request_put[13] vssd1 vssd1 vccd1 vccd1 _1472_/A sky130_fd_sc_hd__clkbuf_1
Xinput107 core_dmem_request_put[94] vssd1 vssd1 vccd1 vccd1 _2142_/A sky130_fd_sc_hd__buf_2
X_3489_ _3489_/CLK _3489_/D vssd1 vssd1 vccd1 vccd1 _3489_/Q sky130_fd_sc_hd__dfxtp_1
Xinput129 core_imem_request_put[23] vssd1 vssd1 vccd1 vccd1 _1508_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2047__C _2047_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2584__B_N _2473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1423__A _2725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2860_ _2860_/A _2875_/B vssd1 vssd1 vccd1 vccd1 _3299_/D sky130_fd_sc_hd__nand2_1
XFILLER_43_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1811_ _3116_/A _1821_/B _1811_/C vssd1 vssd1 vccd1 vccd1 _1811_/Y sky130_fd_sc_hd__nand3_2
X_2791_ _3265_/Q _2779_/X _1815_/Y vssd1 vssd1 vccd1 vccd1 _2792_/A sky130_fd_sc_hd__o21ai_1
X_1742_ _2763_/B vssd1 vssd1 vccd1 vccd1 _1742_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_1_1_0_CLK_A clkbuf_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1673_ _1673_/A _1661_/X vssd1 vssd1 vccd1 vccd1 _1673_/X sky130_fd_sc_hd__or2b_1
X_3412_ _3456_/CLK _3412_/D vssd1 vssd1 vccd1 vccd1 _3412_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _3440_/CLK _3343_/D vssd1 vssd1 vccd1 vccd1 _3343_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _3337_/CLK _3274_/D vssd1 vssd1 vccd1 vccd1 _3274_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ _2225_/A vssd1 vssd1 vccd1 vccd1 _2225_/X sky130_fd_sc_hd__clkbuf_2
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2156_ _2156_/A vssd1 vssd1 vccd1 vccd1 _2156_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2087_ _2087_/A vssd1 vssd1 vccd1 vccd1 _2088_/C sky130_fd_sc_hd__inv_2
XFILLER_53_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2989_ _3003_/A vssd1 vssd1 vccd1 vccd1 _2989_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1756__A1 _1691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input201_A fmc_imem_response_put[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2074__A _2794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input97_A core_dmem_request_put[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output420_A _2070_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2010_ _2010_/A vssd1 vssd1 vccd1 vccd1 _2011_/C sky130_fd_sc_hd__inv_2
XFILLER_82_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2912_ _2950_/A vssd1 vssd1 vccd1 vccd1 _2912_/X sky130_fd_sc_hd__clkbuf_2
X_2843_ _3291_/Q _2835_/X _1917_/Y vssd1 vssd1 vccd1 vccd1 _2844_/A sky130_fd_sc_hd__o21ai_1
XFILLER_31_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2774_ _2774_/A vssd1 vssd1 vccd1 vccd1 _3259_/D sky130_fd_sc_hd__clkbuf_1
X_1725_ _2756_/B vssd1 vssd1 vccd1 vccd1 _1725_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1738__A1 _1734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1656_ _1743_/A vssd1 vssd1 vccd1 vccd1 _1656_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1587_ _1473_/C _1562_/X _1586_/Y vssd1 vssd1 vccd1 vccd1 _1587_/Y sky130_fd_sc_hd__o21ai_2
X_3326_ _3420_/CLK _3326_/D vssd1 vssd1 vccd1 vccd1 _3326_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3112__B1 _3003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _3297_/CLK _3257_/D vssd1 vssd1 vccd1 vccd1 _3257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2208_ _1832_/C _2195_/X _2207_/Y vssd1 vssd1 vccd1 vccd1 _2208_/Y sky130_fd_sc_hd__o21ai_1
X_3188_ _3221_/CLK _3188_/D vssd1 vssd1 vccd1 vccd1 _3188_/Q sky130_fd_sc_hd__dfxtp_1
X_2139_ _2139_/A vssd1 vssd1 vccd1 vccd1 _2140_/C sky130_fd_sc_hd__inv_2
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input151_A fmc_dmem_response_put[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input249_A ram_imem_response_put[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input12_A EN_ram_imem_response_put vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output468_A _1521_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output370_A _1907_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1510_ _3184_/Q _1498_/X _1509_/Y vssd1 vssd1 vccd1 vccd1 _1510_/X sky130_fd_sc_hd__o21a_2
X_2490_ _2542_/A vssd1 vssd1 vccd1 vccd1 _2490_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1441_ _1514_/A vssd1 vssd1 vccd1 vccd1 _1441_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3111_ _3455_/Q _2174_/A _2448_/Y _3103_/X vssd1 vssd1 vccd1 vccd1 _3455_/D sky130_fd_sc_hd__o211a_1
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3042_ _1960_/C _3035_/X _3039_/X _2307_/Y vssd1 vssd1 vccd1 vccd1 _3404_/D sky130_fd_sc_hd__o211ai_1
XFILLER_48_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2826_ _2864_/A vssd1 vssd1 vccd1 vccd1 _2826_/X sky130_fd_sc_hd__clkbuf_2
X_2757_ _2757_/A vssd1 vssd1 vccd1 vccd1 _2757_/X sky130_fd_sc_hd__buf_2
X_2688_ _3196_/Q _2681_/X _1556_/Y _2684_/X vssd1 vssd1 vccd1 vccd1 _3196_/D sky130_fd_sc_hd__o211a_1
X_1708_ _2752_/B vssd1 vssd1 vccd1 vccd1 _1708_/Y sky130_fd_sc_hd__inv_2
X_1639_ _1633_/X _1639_/A2 _1636_/X _1638_/X vssd1 vssd1 vccd1 vccd1 _2734_/B sky130_fd_sc_hd__a22oi_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A EN_core_imem_response_get vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3309_ _3410_/CLK _3309_/D vssd1 vssd1 vccd1 vccd1 _3309_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1894__C _1894_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input199_A fmc_imem_response_put[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_0_0_CLK_A clkbuf_2_1_0_CLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_CLK_A clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1990_ _2018_/A _1990_/B _1990_/C vssd1 vssd1 vccd1 vccd1 _1990_/Y sky130_fd_sc_hd__nand3_1
XFILLER_60_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2611_ _3126_/A _2611_/B vssd1 vssd1 vccd1 vccd1 _3156_/D sky130_fd_sc_hd__nor2_1
XANTENNA__2366__A1 _2033_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2542_ _2542_/A vssd1 vssd1 vccd1 vccd1 _2542_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2473_ _2473_/A vssd1 vssd1 vccd1 vccd1 _2473_/X sky130_fd_sc_hd__clkbuf_2
X_1424_ _3161_/Q _1415_/X _1423_/Y vssd1 vssd1 vccd1 vccd1 _1424_/X sky130_fd_sc_hd__o21a_2
XANTENNA__2669__A2 _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3025_ _3067_/A vssd1 vssd1 vccd1 vccd1 _3025_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2809_ _2809_/A _2818_/B vssd1 vssd1 vccd1 vccd1 _3273_/D sky130_fd_sc_hd__nand2_1
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput561 _2418_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[81] sky130_fd_sc_hd__buf_2
Xoutput572 _2443_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[91] sky130_fd_sc_hd__buf_2
Xoutput550 _2390_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[71] sky130_fd_sc_hd__buf_2
Xoutput583 _1581_/X vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[10] sky130_fd_sc_hd__buf_2
Xoutput594 _1609_/X vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[20] sky130_fd_sc_hd__buf_2
XFILLER_86_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input114_A core_imem_request_put[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2810__A _2868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output333_A _1746_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1973_ _1973_/A vssd1 vssd1 vccd1 vccd1 _1974_/C sky130_fd_sc_hd__inv_2
X_2525_ _2499_/X _3474_/Q _2500_/X vssd1 vssd1 vccd1 vccd1 _2525_/X sky130_fd_sc_hd__o21ba_1
XFILLER_88_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2456_ _2169_/X _2162_/X _2185_/X _3458_/Q vssd1 vssd1 vccd1 vccd1 _2456_/X sky130_fd_sc_hd__a22o_2
X_2387_ _2384_/X _2385_/X _2386_/X _2058_/C _2377_/X vssd1 vssd1 vccd1 vccd1 _2387_/Y
+ sky130_fd_sc_hd__o311ai_2
XFILLER_68_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3008_ _3381_/Q _3007_/X _2243_/Y _3003_/X vssd1 vssd1 vccd1 vccd1 _3381_/D sky130_fd_sc_hd__o211a_1
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput380 _1939_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[37] sky130_fd_sc_hd__buf_2
Xoutput391 _1975_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[47] sky130_fd_sc_hd__buf_2
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input231_A ram_dmem_response_put[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_43_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3482_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_output450_A _1424_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2310_ _3405_/Q _2297_/X _2309_/Y vssd1 vssd1 vccd1 vccd1 _2310_/X sky130_fd_sc_hd__o21a_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ _3486_/CLK _3290_/D vssd1 vssd1 vccd1 vccd1 _3290_/Q sky130_fd_sc_hd__dfxtp_1
X_2241_ _2299_/A vssd1 vssd1 vccd1 vccd1 _2241_/X sky130_fd_sc_hd__buf_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2172_ _2973_/A vssd1 vssd1 vccd1 vccd1 _3093_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1956_ _1963_/A _1971_/B _1956_/C vssd1 vssd1 vccd1 vccd1 _1956_/Y sky130_fd_sc_hd__nand3_1
X_1887_ _1887_/A vssd1 vssd1 vccd1 vccd1 _1888_/C sky130_fd_sc_hd__clkinv_4
Xclkbuf_leaf_34_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3337_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2193__C1 _2152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2508_ _2499_/X _3470_/Q _2500_/X vssd1 vssd1 vccd1 vccd1 _2508_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__1758__B1_N _1743_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3488_ _3489_/CLK _3488_/D vssd1 vssd1 vccd1 vccd1 _3488_/Q sky130_fd_sc_hd__dfxtp_1
Xinput108 core_dmem_request_put[95] vssd1 vssd1 vccd1 vccd1 _2146_/A sky130_fd_sc_hd__buf_2
XFILLER_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2439_ _2459_/B vssd1 vssd1 vccd1 vccd1 _2439_/X sky130_fd_sc_hd__buf_2
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput119 core_imem_request_put[14] vssd1 vssd1 vccd1 vccd1 _1475_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_84_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_33_CLK_A clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_48_CLK_A clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2625__A _2677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_25_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3452_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_input181_A fmc_imem_response_put[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input42_A core_dmem_request_put[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2535__A _2535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1810_ _1810_/A vssd1 vssd1 vccd1 vccd1 _1811_/C sky130_fd_sc_hd__inv_6
XFILLER_30_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2790_ _3264_/Q _2789_/X _2784_/X _1811_/Y vssd1 vssd1 vccd1 vccd1 _3264_/D sky130_fd_sc_hd__o211a_1
XFILLER_7_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1741_ _1712_/X _1741_/A2 _1739_/X _1740_/X vssd1 vssd1 vccd1 vccd1 _2763_/B sky130_fd_sc_hd__a22oi_4
Xclkbuf_leaf_16_CLK clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3459_/CLK sky130_fd_sc_hd__clkbuf_16
X_1672_ _1670_/X _3233_/Q _1671_/X vssd1 vssd1 vccd1 vccd1 _1672_/X sky130_fd_sc_hd__o21ba_1
X_3411_ _3413_/CLK _3411_/D vssd1 vssd1 vccd1 vccd1 _3411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3342_ _3447_/CLK _3342_/D vssd1 vssd1 vccd1 vccd1 _3342_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1517__A2 _1514_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _3337_/CLK _3273_/D vssd1 vssd1 vccd1 vccd1 _3273_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2224_ _2253_/A vssd1 vssd1 vccd1 vccd1 _2224_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2155_ _2412_/A vssd1 vssd1 vccd1 vccd1 _2156_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_66_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2086_ _2206_/A vssd1 vssd1 vccd1 vccd1 _2117_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2988_ _3095_/A vssd1 vssd1 vccd1 vccd1 _3003_/A sky130_fd_sc_hd__clkbuf_4
X_1939_ _3297_/Q _1929_/X _1938_/Y vssd1 vssd1 vccd1 vccd1 _1939_/X sky130_fd_sc_hd__o21a_2
XANTENNA__1756__A2 _1756_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput90 core_dmem_request_put[79] vssd1 vssd1 vccd1 vccd1 _2090_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__2705__A1 _1480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2355__A _2459_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3121__A1 _3461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output413_A _2048_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2880__B1 _2864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_CLK clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3226_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2265__A _2351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2911_ _3326_/Q _2907_/X _2903_/X _2044_/Y vssd1 vssd1 vccd1 vccd1 _3326_/D sky130_fd_sc_hd__o211a_1
XFILLER_50_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2842_ _3290_/Q _2830_/X _2826_/X _1913_/Y vssd1 vssd1 vccd1 vccd1 _3290_/D sky130_fd_sc_hd__o211a_1
X_2773_ _2747_/A _2773_/B vssd1 vssd1 vccd1 vccd1 _2774_/A sky130_fd_sc_hd__and2b_1
X_1724_ _1712_/X _1724_/A2 _1722_/X _1723_/X vssd1 vssd1 vccd1 vccd1 _2756_/B sky130_fd_sc_hd__a22oi_4
XANTENNA__1738__A2 _2762_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1655_ _2737_/B vssd1 vssd1 vccd1 vccd1 _1655_/Y sky130_fd_sc_hd__inv_2
X_1586_ _1563_/X _1569_/X _3207_/Q vssd1 vssd1 vccd1 vccd1 _1586_/Y sky130_fd_sc_hd__o21ai_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ _3436_/CLK _3325_/D vssd1 vssd1 vccd1 vccd1 _3325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _3258_/CLK _3256_/D vssd1 vssd1 vccd1 vccd1 _3256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2207_ _2196_/X _2206_/X _3370_/Q vssd1 vssd1 vccd1 vccd1 _2207_/Y sky130_fd_sc_hd__o21ai_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3187_ _3404_/CLK _3187_/D vssd1 vssd1 vccd1 vccd1 _3187_/Q sky130_fd_sc_hd__dfxtp_1
X_2138_ _3352_/Q _2129_/X _2137_/Y vssd1 vssd1 vccd1 vccd1 _2138_/X sky130_fd_sc_hd__o21a_1
XFILLER_66_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2175__A _2175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2069_ _2091_/A _2099_/B _2069_/C vssd1 vssd1 vccd1 vccd1 _2069_/Y sky130_fd_sc_hd__nand3_1
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1729__A2 _2759_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input144_A core_imem_request_put[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1429__A _1443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output363_A _1878_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1440_ _2618_/A vssd1 vssd1 vccd1 vccd1 _1514_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_output530_A _2337_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3110_ _2140_/C _3105_/X _3003_/A _2446_/Y vssd1 vssd1 vccd1 vccd1 _3454_/D sky130_fd_sc_hd__o211ai_1
XFILLER_4_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3041_ _3403_/Q _3037_/X _2305_/Y _3033_/X vssd1 vssd1 vccd1 vccd1 _3403_/D sky130_fd_sc_hd__o211a_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2723__A _2723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2825_ _2825_/A _2837_/B vssd1 vssd1 vccd1 vccd1 _3281_/D sky130_fd_sc_hd__nand2_1
X_2756_ _2756_/A _2756_/B vssd1 vssd1 vccd1 vccd1 _3245_/D sky130_fd_sc_hd__nor2_1
X_2687_ _1429_/C _1618_/X _2686_/X _1554_/Y vssd1 vssd1 vccd1 vccd1 _3195_/D sky130_fd_sc_hd__o211ai_1
X_1707_ _1669_/X _1707_/A2 _1704_/X _1706_/X vssd1 vssd1 vccd1 vccd1 _2752_/B sky130_fd_sc_hd__a22oi_4
X_1638_ _1638_/A _1637_/X vssd1 vssd1 vccd1 vccd1 _1638_/X sky130_fd_sc_hd__or2b_1
X_1569_ _2675_/B vssd1 vssd1 vccd1 vccd1 _1569_/X sky130_fd_sc_hd__clkbuf_2
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3308_ _3394_/CLK _3308_/D vssd1 vssd1 vccd1 vccd1 _3308_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ _3476_/CLK _3239_/D vssd1 vssd1 vccd1 vccd1 _3239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input261_A ram_imem_response_put[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2543__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output480_A _1457_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2610_ _3130_/A vssd1 vssd1 vccd1 vccd1 _3126_/A sky130_fd_sc_hd__buf_2
X_2541_ _2541_/A vssd1 vssd1 vccd1 vccd1 _2541_/X sky130_fd_sc_hd__buf_4
XFILLER_5_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2472_ _2605_/B vssd1 vssd1 vccd1 vccd1 _2473_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2118__A2 _2111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1423_ _2725_/A _1447_/B _1423_/C vssd1 vssd1 vccd1 vccd1 _1423_/Y sky130_fd_sc_hd__nand3_2
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3024_ _3391_/Q _3023_/X _2272_/Y _3019_/X vssd1 vssd1 vccd1 vccd1 _3391_/D sky130_fd_sc_hd__o211a_1
XFILLER_55_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2808_ _3273_/Q _2795_/X _1847_/Y vssd1 vssd1 vccd1 vccd1 _2809_/A sky130_fd_sc_hd__o21ai_1
X_2739_ _2743_/A _2739_/B vssd1 vssd1 vccd1 vccd1 _3231_/D sky130_fd_sc_hd__nor2_1
Xoutput551 _2392_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[72] sky130_fd_sc_hd__buf_2
Xoutput540 _2364_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[62] sky130_fd_sc_hd__buf_2
Xoutput562 _2420_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[82] sky130_fd_sc_hd__buf_2
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput584 _1583_/Y vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[11] sky130_fd_sc_hd__buf_2
Xoutput595 _1611_/Y vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[21] sky130_fd_sc_hd__buf_2
Xoutput573 _2445_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[92] sky130_fd_sc_hd__buf_2
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input107_A core_dmem_request_put[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2596__A2 _2613_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input72_A core_dmem_request_put[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1556__B1 _1432_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output326_A _1721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1972_ _3306_/Q _1965_/X _1971_/Y vssd1 vssd1 vccd1 vccd1 _1972_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2524_ _2520_/X _3136_/A2 _2522_/X _2523_/X vssd1 vssd1 vccd1 vccd1 _2524_/X sky130_fd_sc_hd__a22o_1
X_2455_ _3457_/Q _2439_/X _2454_/Y vssd1 vssd1 vccd1 vccd1 _2455_/X sky130_fd_sc_hd__o21a_1
X_2386_ _2414_/A vssd1 vssd1 vccd1 vccd1 _2386_/X sky130_fd_sc_hd__buf_2
XFILLER_68_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3007_ _3037_/A vssd1 vssd1 vccd1 vccd1 _3007_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2275__A1 _1917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2578__A2 _2578_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_7_CLK_A clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput370 _1907_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[28] sky130_fd_sc_hd__buf_2
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput392 _1979_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[48] sky130_fd_sc_hd__buf_2
Xoutput381 _1943_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[38] sky130_fd_sc_hd__buf_2
XFILLER_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input224_A ram_dmem_response_put[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2821__A _2878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output276_A _1411_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ _2298_/A vssd1 vssd1 vccd1 vccd1 _2240_/X sky130_fd_sc_hd__buf_2
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2171_ _2175_/A _2177_/A _2179_/A _2163_/A vssd1 vssd1 vccd1 vccd1 _2973_/A sky130_fd_sc_hd__o31a_2
XFILLER_38_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2257__A1 _1894_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1955_ _1955_/A vssd1 vssd1 vccd1 vccd1 _1956_/C sky130_fd_sc_hd__clkinv_4
X_1886_ _3283_/Q _1871_/X _1885_/Y vssd1 vssd1 vccd1 vccd1 _1886_/X sky130_fd_sc_hd__o21a_2
XFILLER_88_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2193__B1 _1811_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2507_ _2471_/X _3132_/A2 _2505_/X _2506_/X vssd1 vssd1 vccd1 vccd1 _2507_/X sky130_fd_sc_hd__a22o_1
X_3487_ _3489_/CLK _3487_/D vssd1 vssd1 vccd1 vccd1 _3487_/Q sky130_fd_sc_hd__dfxtp_1
Xinput109 core_dmem_request_put[96] vssd1 vssd1 vccd1 vccd1 _2151_/A sky130_fd_sc_hd__clkbuf_4
X_2438_ _2127_/C _2426_/X _2437_/Y vssd1 vssd1 vccd1 vccd1 _2438_/Y sky130_fd_sc_hd__o21ai_2
X_2369_ _2397_/A vssd1 vssd1 vccd1 vccd1 _2369_/X sky130_fd_sc_hd__buf_4
XFILLER_56_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2641__A _2660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input174_A fmc_dmem_response_put[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input35_A core_dmem_request_put[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1423__C _1423_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2816__A _2893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1720__A _1720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output393_A _1982_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1740_ _1740_/A _1705_/X vssd1 vssd1 vccd1 vccd1 _1740_/X sky130_fd_sc_hd__or2b_1
XFILLER_7_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1671_ _1743_/A vssd1 vssd1 vccd1 vccd1 _1671_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3410_ _3410_/CLK _3410_/D vssd1 vssd1 vccd1 vccd1 _3410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3341_ _3440_/CLK _3341_/D vssd1 vssd1 vccd1 vccd1 _3341_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _3337_/CLK _3272_/D vssd1 vssd1 vccd1 vccd1 _3272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ _3375_/Q _2210_/X _2222_/Y vssd1 vssd1 vccd1 vccd1 _2223_/X sky130_fd_sc_hd__o21a_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2154_ _2175_/A vssd1 vssd1 vccd1 vccd1 _2412_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1630__A _3226_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2085_ _3337_/Q _2075_/X _2084_/Y vssd1 vssd1 vccd1 vccd1 _2085_/X sky130_fd_sc_hd__o21a_2
XFILLER_34_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2987_ _1824_/C _2451_/X _2980_/X _2201_/Y vssd1 vssd1 vccd1 vccd1 _3368_/D sky130_fd_sc_hd__o211ai_1
XANTENNA__2461__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1938_ _1945_/A _1953_/B _1938_/C vssd1 vssd1 vccd1 vccd1 _1938_/Y sky130_fd_sc_hd__nand3_1
X_1869_ _1869_/A _1877_/B _1869_/C vssd1 vssd1 vccd1 vccd1 _1869_/Y sky130_fd_sc_hd__nand3_1
Xinput80 core_dmem_request_put[6] vssd1 vssd1 vccd1 vccd1 _1820_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput91 core_dmem_request_put[7] vssd1 vssd1 vccd1 vccd1 _1823_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_88_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3121__A2 _2439_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2910_ _2910_/A _2914_/B vssd1 vssd1 vccd1 vccd1 _3325_/D sky130_fd_sc_hd__nand2_1
X_2841_ _2841_/A _2856_/B vssd1 vssd1 vccd1 vccd1 _3289_/D sky130_fd_sc_hd__nand2_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2772_ _1633_/X _2772_/A2 _1773_/X _1774_/X _2747_/A vssd1 vssd1 vccd1 vccd1 _3258_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_32_CLK_A clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1723_ _1723_/A _1705_/X vssd1 vssd1 vccd1 vccd1 _1723_/X sky130_fd_sc_hd__or2b_1
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1654_ _1633_/X _1654_/A2 _1652_/X _1653_/X vssd1 vssd1 vccd1 vccd1 _2737_/B sky130_fd_sc_hd__a22oi_2
X_1585_ _3206_/Q _1576_/X _1584_/Y vssd1 vssd1 vccd1 vccd1 _1585_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2699__A1 _1460_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3324_ _3420_/CLK _3324_/D vssd1 vssd1 vccd1 vccd1 _3324_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_47_CLK_A clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _3297_/CLK _3255_/D vssd1 vssd1 vccd1 vccd1 _3255_/Q sky130_fd_sc_hd__dfxtp_1
X_2206_ _2206_/A vssd1 vssd1 vccd1 vccd1 _2206_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3112__A2 _3105_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _3221_/CLK _3186_/D vssd1 vssd1 vccd1 vccd1 _3186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2137_ _2143_/A _2152_/B _2137_/C vssd1 vssd1 vccd1 vccd1 _2137_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__1674__A2 _1674_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2068_ _2068_/A vssd1 vssd1 vccd1 vccd1 _2069_/C sky130_fd_sc_hd__inv_2
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1535__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2069__C _2069_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input137_A core_imem_request_put[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1429__B _1452_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output523_A _2318_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput270 ram_imem_response_put[6] vssd1 vssd1 vccd1 vccd1 _1673_/A sky130_fd_sc_hd__buf_2
X_3040_ _1953_/C _3035_/X _3039_/X _2303_/Y vssd1 vssd1 vccd1 vccd1 _3402_/D sky130_fd_sc_hd__o211ai_1
XFILLER_48_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2824_ _3281_/Q _2816_/X _1877_/Y vssd1 vssd1 vccd1 vccd1 _2825_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__3030__A1 _1931_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2755_ _2744_/X _2755_/A2 _1719_/X _1720_/X _2745_/X vssd1 vssd1 vccd1 vccd1 _3244_/D
+ sky130_fd_sc_hd__a221o_1
X_2686_ _2686_/A vssd1 vssd1 vccd1 vccd1 _2686_/X sky130_fd_sc_hd__clkbuf_2
X_1706_ _1706_/A _1705_/X vssd1 vssd1 vccd1 vccd1 _1706_/X sky130_fd_sc_hd__or2b_1
X_1637_ _1776_/B vssd1 vssd1 vccd1 vccd1 _1637_/X sky130_fd_sc_hd__buf_2
X_1568_ _3200_/Q _1545_/X _1567_/Y vssd1 vssd1 vccd1 vccd1 _1568_/X sky130_fd_sc_hd__o21a_1
X_3307_ _3410_/CLK _3307_/D vssd1 vssd1 vccd1 vccd1 _3307_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1499_ _1499_/A vssd1 vssd1 vccd1 vccd1 _1500_/C sky130_fd_sc_hd__inv_2
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ _3258_/CLK _3238_/D vssd1 vssd1 vccd1 vccd1 _3238_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2186__A _2206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3169_ _3482_/CLK _3169_/D vssd1 vssd1 vccd1 vccd1 _3169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1583__A1 _1467_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input254_A ram_imem_response_put[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2063__A2 _2056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output473_A _1539_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2540_ _2520_/X _3142_/A2 _2538_/X _2539_/X vssd1 vssd1 vccd1 vccd1 _2540_/X sky130_fd_sc_hd__a22o_1
X_2471_ _2520_/A vssd1 vssd1 vccd1 vccd1 _2471_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1422_ _1422_/A vssd1 vssd1 vccd1 vccd1 _1423_/C sky130_fd_sc_hd__clkinv_4
XFILLER_68_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3023_ _3037_/A vssd1 vssd1 vccd1 vccd1 _3023_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2807_ _3272_/Q _2789_/X _2806_/X _1843_/Y vssd1 vssd1 vccd1 vccd1 _3272_/D sky130_fd_sc_hd__o211a_1
XFILLER_3_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2738_ _1772_/X _2738_/A2 _1657_/X _1658_/X _2771_/A vssd1 vssd1 vccd1 vccd1 _3230_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1565__A1 _1443_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput530 _2337_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[53] sky130_fd_sc_hd__buf_2
Xoutput541 _2366_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[63] sky130_fd_sc_hd__buf_2
Xoutput563 _2422_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[83] sky130_fd_sc_hd__buf_2
Xoutput552 _2394_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[73] sky130_fd_sc_hd__buf_2
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2669_ _3186_/Q _1415_/A _1516_/Y vssd1 vssd1 vccd1 vccd1 _2670_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__1516__C _1516_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput585 _1585_/X vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[12] sky130_fd_sc_hd__buf_2
Xoutput574 _2447_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[93] sky130_fd_sc_hd__buf_2
Xoutput596 _1613_/X vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[22] sky130_fd_sc_hd__buf_2
XFILLER_59_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2644__A _2660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2045__A2 _2038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input65_A core_dmem_request_put[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1723__A _1723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1971_ _2000_/A _1971_/B _1971_/C vssd1 vssd1 vccd1 vccd1 _1971_/Y sky130_fd_sc_hd__nand3_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2523_ _2523_/A _2513_/X vssd1 vssd1 vccd1 vccd1 _2523_/X sky130_fd_sc_hd__or2b_1
X_2454_ _2156_/A _2159_/A _2162_/A _2152_/C _2434_/X vssd1 vssd1 vccd1 vccd1 _2454_/Y
+ sky130_fd_sc_hd__o311ai_4
X_2385_ _2413_/A vssd1 vssd1 vccd1 vccd1 _2385_/X sky130_fd_sc_hd__buf_2
XFILLER_56_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput1 EN_core_dmem_request_put vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_4
XFILLER_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3006_ _1869_/C _3005_/X _2995_/X _2237_/Y vssd1 vssd1 vccd1 vccd1 _3380_/D sky130_fd_sc_hd__o211ai_1
XFILLER_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2027__A2 _2020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1527__B _1527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput371 _1910_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[29] sky130_fd_sc_hd__buf_2
Xoutput360 _1870_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[19] sky130_fd_sc_hd__buf_2
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput393 _1982_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[49] sky130_fd_sc_hd__buf_2
Xoutput382 _1946_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[39] sky130_fd_sc_hd__buf_2
XFILLER_59_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2077__C _2077_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input217_A ram_dmem_response_put[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2549__A _2549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2170_ _2169_/X _1821_/B _3360_/Q vssd1 vssd1 vccd1 vccd1 _2170_/X sky130_fd_sc_hd__a21o_1
XFILLER_38_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output603_A _1627_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2284__A _2370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2009__A2 _2002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1954_ _3301_/Q _1947_/X _1953_/Y vssd1 vssd1 vccd1 vccd1 _1954_/X sky130_fd_sc_hd__o21a_2
XANTENNA__2731__B _2975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1768__A1 _1637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1885_ _1909_/A _1917_/B _1885_/C vssd1 vssd1 vccd1 vccd1 _1885_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2506_ _2506_/A _2478_/X vssd1 vssd1 vccd1 vccd1 _2506_/X sky130_fd_sc_hd__or2b_1
X_3486_ _3486_/CLK _3486_/D vssd1 vssd1 vccd1 vccd1 _3486_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2459__A _3461_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2437_ _2427_/X _1801_/B _3450_/Q vssd1 vssd1 vccd1 vccd1 _2437_/Y sky130_fd_sc_hd__o21ai_1
X_2368_ _3425_/Q _2355_/X _2367_/Y vssd1 vssd1 vccd1 vccd1 _2368_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2496__A2 _3129_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2299_ _2299_/A vssd1 vssd1 vccd1 vccd1 _2299_/X sky130_fd_sc_hd__buf_2
XFILLER_71_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input167_A fmc_dmem_response_put[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2369__A _2397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input28_A core_dmem_request_put[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2775__B_N _2975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output386_A _1957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1670_ _1713_/A vssd1 vssd1 vccd1 vccd1 _1670_/X sky130_fd_sc_hd__clkbuf_2
X_3340_ _3447_/CLK _3340_/D vssd1 vssd1 vccd1 vccd1 _3340_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3271_/CLK _3271_/D vssd1 vssd1 vccd1 vccd1 _3271_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _2211_/X _2212_/X _2213_/X _1850_/C _2203_/X vssd1 vssd1 vccd1 vccd1 _2222_/Y
+ sky130_fd_sc_hd__o311ai_4
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2153_ _3356_/Q _2145_/X _2152_/Y vssd1 vssd1 vccd1 vccd1 _2153_/X sky130_fd_sc_hd__o21a_1
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_6_CLK_A clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1630__B _1630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2084_ _2091_/A _2099_/B _2084_/C vssd1 vssd1 vccd1 vccd1 _2084_/Y sky130_fd_sc_hd__nand3_1
XFILLER_61_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2986_ _3367_/Q _2974_/X _2199_/Y _2978_/X vssd1 vssd1 vccd1 vccd1 _3367_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1937_ _1937_/A vssd1 vssd1 vccd1 vccd1 _1938_/C sky130_fd_sc_hd__inv_2
X_1868_ _1868_/A vssd1 vssd1 vccd1 vccd1 _1869_/C sky130_fd_sc_hd__clkinv_4
Xinput70 core_dmem_request_put[60] vssd1 vssd1 vccd1 vccd1 _2021_/A sky130_fd_sc_hd__buf_2
Xinput81 core_dmem_request_put[70] vssd1 vssd1 vccd1 vccd1 _2057_/A sky130_fd_sc_hd__buf_2
X_1799_ _2408_/A vssd1 vssd1 vccd1 vccd1 _1801_/B sky130_fd_sc_hd__clkbuf_4
Xinput92 core_dmem_request_put[80] vssd1 vssd1 vccd1 vccd1 _2094_/A sky130_fd_sc_hd__buf_2
XANTENNA__3115__B1 _3105_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3469_ _3476_/CLK _3469_/D vssd1 vssd1 vccd1 vccd1 _3469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2917__A _2936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1731__A _1731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2880__A2 _2868_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2840_ _2878_/A vssd1 vssd1 vccd1 vccd1 _2856_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2771_ _2771_/A _2771_/B vssd1 vssd1 vccd1 vccd1 _3257_/D sky130_fd_sc_hd__nor2_1
X_1722_ _1713_/X _3245_/Q _1714_/X vssd1 vssd1 vccd1 vccd1 _1722_/X sky130_fd_sc_hd__o21ba_1
X_1653_ _1653_/A _1637_/X vssd1 vssd1 vccd1 vccd1 _1653_/X sky130_fd_sc_hd__or2b_1
X_1584_ _1577_/X _1578_/X _1579_/X _1470_/C _1566_/X vssd1 vssd1 vccd1 vccd1 _1584_/Y
+ sky130_fd_sc_hd__o311ai_4
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3323_ _3432_/CLK _3323_/D vssd1 vssd1 vccd1 vccd1 _3323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3254_ _3410_/CLK _3254_/D vssd1 vssd1 vccd1 vccd1 _3254_/Q sky130_fd_sc_hd__dfxtp_1
X_2205_ _3369_/Q _2174_/X _2204_/Y vssd1 vssd1 vccd1 vccd1 _2205_/X sky130_fd_sc_hd__o21a_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3185_ _3404_/CLK _3185_/D vssd1 vssd1 vccd1 vccd1 _3185_/Q sky130_fd_sc_hd__dfxtp_1
X_2136_ _2136_/A vssd1 vssd1 vccd1 vccd1 _2137_/C sky130_fd_sc_hd__clkinv_2
XFILLER_19_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2067_ _2104_/A vssd1 vssd1 vccd1 vccd1 _2099_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2472__A _2605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2969_ _2969_/A _2969_/B _3358_/Q vssd1 vssd1 vccd1 vccd1 _2970_/A sky130_fd_sc_hd__and3_1
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input95_A core_dmem_request_put[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1429__C _1429_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput271 ram_imem_response_put[7] vssd1 vssd1 vccd1 vccd1 _1677_/A sky130_fd_sc_hd__clkbuf_2
Xinput260 ram_imem_response_put[26] vssd1 vssd1 vccd1 vccd1 _1755_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2557__A _2557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2823_ _3280_/Q _2810_/X _2806_/X _1873_/Y vssd1 vssd1 vccd1 vccd1 _3280_/D sky130_fd_sc_hd__o211a_1
X_2754_ _2756_/A _2754_/B vssd1 vssd1 vccd1 vccd1 _3243_/D sky130_fd_sc_hd__nor2_1
X_1705_ _1713_/A vssd1 vssd1 vccd1 vccd1 _1705_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2685_ _3194_/Q _2681_/X _1549_/Y _2684_/X vssd1 vssd1 vccd1 vccd1 _3194_/D sky130_fd_sc_hd__o211a_1
X_1636_ _1635_/X _3227_/Q _1641_/A vssd1 vssd1 vccd1 vccd1 _1636_/X sky130_fd_sc_hd__o21ba_1
X_1567_ _1546_/X _1547_/X _1548_/X _1447_/C _1566_/X vssd1 vssd1 vccd1 vccd1 _1567_/Y
+ sky130_fd_sc_hd__o311ai_4
X_3306_ _3456_/CLK _3306_/D vssd1 vssd1 vccd1 vccd1 _3306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ _1514_/A vssd1 vssd1 vccd1 vccd1 _1498_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2467__A _2467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3237_ _3472_/CLK _3237_/D vssd1 vssd1 vccd1 vccd1 _3237_/Q sky130_fd_sc_hd__dfxtp_1
X_3168_ _3482_/CLK _3168_/D vssd1 vssd1 vccd1 vccd1 _3168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2119_ _2119_/A vssd1 vssd1 vccd1 vccd1 _2120_/C sky130_fd_sc_hd__inv_2
X_3099_ _3445_/Q _3093_/X _2423_/Y _3089_/X vssd1 vssd1 vccd1 vccd1 _3445_/D sky130_fd_sc_hd__o211a_1
XFILLER_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input247_A ram_imem_response_put[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input10_A EN_ram_dmem_response_put vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_31_CLK_A clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2599__A1 _2520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_46_CLK_A clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2840__A _2878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2470_ _2470_/A vssd1 vssd1 vccd1 vccd1 _2520_/A sky130_fd_sc_hd__buf_4
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1421_ _2675_/B vssd1 vssd1 vccd1 vccd1 _1447_/B sky130_fd_sc_hd__buf_2
XFILLER_95_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2287__B1 _1935_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3022_ _1909_/C _3021_/X _3010_/X _2266_/Y vssd1 vssd1 vccd1 vccd1 _3390_/D sky130_fd_sc_hd__o211ai_1
XFILLER_24_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2806_ _2864_/A vssd1 vssd1 vccd1 vccd1 _2806_/X sky130_fd_sc_hd__clkbuf_2
X_2737_ _2743_/A _2737_/B vssd1 vssd1 vccd1 vccd1 _3229_/D sky130_fd_sc_hd__nor2_1
Xoutput520 _2310_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[44] sky130_fd_sc_hd__buf_2
X_2668_ _3185_/Q _2660_/X _2661_/X _1512_/Y vssd1 vssd1 vccd1 vccd1 _3185_/D sky130_fd_sc_hd__o211a_1
Xoutput531 _2339_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[54] sky130_fd_sc_hd__buf_2
Xoutput553 _2396_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[74] sky130_fd_sc_hd__buf_2
Xoutput542 _2368_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[64] sky130_fd_sc_hd__buf_2
X_1619_ _1563_/A _1597_/X _3219_/Q vssd1 vssd1 vccd1 vccd1 _1619_/Y sky130_fd_sc_hd__o21ai_2
Xoutput575 _2449_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[94] sky130_fd_sc_hd__buf_2
Xoutput586 _1587_/Y vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[13] sky130_fd_sc_hd__buf_2
Xoutput564 _2424_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[84] sky130_fd_sc_hd__buf_2
XFILLER_59_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2599_ _2520_/A _2599_/A2 _2597_/X _2598_/X vssd1 vssd1 vccd1 vccd1 _2614_/B sky130_fd_sc_hd__a22oi_4
Xoutput597 _1615_/Y vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[23] sky130_fd_sc_hd__buf_2
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input2_A EN_core_dmem_response_get vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input197_A fmc_imem_response_put[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2660__A _2660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input58_A core_dmem_request_put[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3491__A _3491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2835__A _2893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1970_ _1970_/A vssd1 vssd1 vccd1 vccd1 _1971_/C sky130_fd_sc_hd__clkinv_2
XFILLER_21_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2992__A1 _1832_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_46_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3476_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2522_ _2521_/X _3473_/Q _2485_/X vssd1 vssd1 vccd1 vccd1 _2522_/X sky130_fd_sc_hd__o21ba_1
X_2453_ _2147_/C _2451_/X _2452_/Y vssd1 vssd1 vccd1 vccd1 _2453_/Y sky130_fd_sc_hd__o21ai_4
X_2384_ _2412_/A vssd1 vssd1 vccd1 vccd1 _2384_/X sky130_fd_sc_hd__buf_2
XFILLER_83_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput2 EN_core_dmem_response_get vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3005_ _3035_/A vssd1 vssd1 vccd1 vccd1 _3005_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2745__A _2760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2983__A1 _1808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3288_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1527__C _1527_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput361 _1802_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[1] sky130_fd_sc_hd__buf_2
Xoutput350 _1795_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[0] sky130_fd_sc_hd__buf_2
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput383 _1809_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[3] sky130_fd_sc_hd__buf_2
Xoutput372 _1805_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[2] sky130_fd_sc_hd__buf_2
Xoutput394 _1812_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[4] sky130_fd_sc_hd__buf_2
XFILLER_74_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input112_A core_dmem_request_put[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3410_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output331_A _1738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output429_A _2100_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1953_ _1981_/A _1953_/B _1953_/C vssd1 vssd1 vccd1 vccd1 _1953_/Y sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_19_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3431_/CLK sky130_fd_sc_hd__clkbuf_16
X_1884_ _1884_/A vssd1 vssd1 vccd1 vccd1 _1885_/C sky130_fd_sc_hd__clkinv_4
XANTENNA__2717__A1 _1509_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2505_ _2473_/X _3469_/Q _2485_/X vssd1 vssd1 vccd1 vccd1 _2505_/X sky130_fd_sc_hd__o21ba_1
X_3485_ _3485_/CLK _3485_/D vssd1 vssd1 vccd1 vccd1 _3485_/Q sky130_fd_sc_hd__dfxtp_1
X_2436_ _3449_/Q _2411_/X _2435_/Y vssd1 vssd1 vccd1 vccd1 _2436_/X sky130_fd_sc_hd__o21a_1
XFILLER_88_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1644__A _1644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2459__B _2459_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2367_ _2356_/X _2357_/X _2358_/X _2036_/C _2348_/X vssd1 vssd1 vccd1 vccd1 _2367_/Y
+ sky130_fd_sc_hd__o311ai_4
XFILLER_56_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2298_ _2298_/A vssd1 vssd1 vccd1 vccd1 _2298_/X sky130_fd_sc_hd__buf_2
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2577__B_N _2473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1819__A _2169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2708__A1 _1488_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output379_A _1936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output281_A _3491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3270_ _3337_/CLK _3270_/D vssd1 vssd1 vccd1 vccd1 _3270_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _1847_/C _2195_/X _2220_/Y vssd1 vssd1 vccd1 vccd1 _2221_/Y sky130_fd_sc_hd__o21ai_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_8_CLK clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3461_/CLK sky130_fd_sc_hd__clkbuf_16
X_2152_ _2152_/A _2152_/B _2152_/C vssd1 vssd1 vccd1 vccd1 _2152_/Y sky130_fd_sc_hd__nand3_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2083_ _2083_/A vssd1 vssd1 vccd1 vccd1 _2084_/C sky130_fd_sc_hd__clkinv_2
XFILLER_81_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2985_ _1815_/C _2451_/X _2980_/X _2197_/Y vssd1 vssd1 vccd1 vccd1 _3366_/D sky130_fd_sc_hd__o211ai_1
X_1936_ _3296_/Q _1929_/X _1935_/Y vssd1 vssd1 vccd1 vccd1 _1936_/X sky130_fd_sc_hd__o21a_2
X_1867_ _3278_/Q _1852_/X _1866_/Y vssd1 vssd1 vccd1 vccd1 _1867_/X sky130_fd_sc_hd__o21a_1
Xinput60 core_dmem_request_put[51] vssd1 vssd1 vccd1 vccd1 _1989_/A sky130_fd_sc_hd__clkbuf_1
Xinput71 core_dmem_request_put[61] vssd1 vssd1 vccd1 vccd1 _2025_/A sky130_fd_sc_hd__clkbuf_1
Xinput82 core_dmem_request_put[71] vssd1 vssd1 vccd1 vccd1 _2061_/A sky130_fd_sc_hd__clkbuf_1
X_1798_ _2235_/A vssd1 vssd1 vccd1 vccd1 _2408_/A sky130_fd_sc_hd__clkbuf_2
Xinput93 core_dmem_request_put[81] vssd1 vssd1 vccd1 vccd1 _2098_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3115__A1 _2169_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3468_ _3472_/CLK _3468_/D vssd1 vssd1 vccd1 vccd1 _3468_/Q sky130_fd_sc_hd__dfxtp_1
X_3399_ _3459_/CLK _3399_/D vssd1 vssd1 vccd1 vccd1 _3399_/Q sky130_fd_sc_hd__dfxtp_1
X_2419_ _2412_/X _2413_/X _2414_/X _2102_/C _2405_/X vssd1 vssd1 vccd1 vccd1 _2419_/Y
+ sky130_fd_sc_hd__o311ai_4
XFILLER_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input40_A core_dmem_request_put[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2865__B1 _2864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2770_ _1633_/X _2770_/A2 _1765_/X _1766_/X _2747_/A vssd1 vssd1 vccd1 vccd1 _3256_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_7_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1721_ _1691_/X _2755_/A2 _1719_/X _1720_/X vssd1 vssd1 vccd1 vccd1 _1721_/X sky130_fd_sc_hd__a22o_2
X_1652_ _1635_/X _3229_/Q _1641_/A vssd1 vssd1 vccd1 vccd1 _1652_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__2148__A2 _2145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1583_ _1467_/C _1562_/X _1582_/Y vssd1 vssd1 vccd1 vccd1 _1583_/Y sky130_fd_sc_hd__o21ai_2
X_3322_ _3330_/CLK _3322_/D vssd1 vssd1 vccd1 vccd1 _3322_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _3297_/CLK _3253_/D vssd1 vssd1 vccd1 vccd1 _3253_/Q sky130_fd_sc_hd__dfxtp_1
X_2204_ _2176_/X _2178_/X _2180_/X _1829_/C _2203_/X vssd1 vssd1 vccd1 vccd1 _2204_/Y
+ sky130_fd_sc_hd__o311ai_2
X_3184_ _3221_/CLK _3184_/D vssd1 vssd1 vccd1 vccd1 _3184_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2135_ _3351_/Q _2129_/X _2134_/Y vssd1 vssd1 vccd1 vccd1 _2135_/X sky130_fd_sc_hd__o21a_1
XFILLER_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2066_ _3332_/Q _2056_/X _2065_/Y vssd1 vssd1 vccd1 vccd1 _2066_/X sky130_fd_sc_hd__o21a_1
XFILLER_26_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2968_ _2969_/A _3357_/Q _2959_/X vssd1 vssd1 vccd1 vccd1 _3357_/D sky130_fd_sc_hd__a21bo_1
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1919_ _1919_/A vssd1 vssd1 vccd1 vccd1 _1920_/C sky130_fd_sc_hd__clkinv_4
XANTENNA__1595__B1 _1484_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2899_ _2899_/A _2914_/B vssd1 vssd1 vccd1 vccd1 _3319_/D sky130_fd_sc_hd__nand2_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input88_A core_dmem_request_put[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_CLK_A clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2550__A2 _3145_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput272 ram_imem_response_put[8] vssd1 vssd1 vccd1 vccd1 _1680_/A sky130_fd_sc_hd__buf_2
Xinput261 ram_imem_response_put[27] vssd1 vssd1 vccd1 vccd1 _1759_/A sky130_fd_sc_hd__clkbuf_2
Xinput250 ram_imem_response_put[17] vssd1 vssd1 vccd1 vccd1 _1720_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output411_A _2041_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2822_ _2822_/A _2837_/B vssd1 vssd1 vccd1 vccd1 _3279_/D sky130_fd_sc_hd__nand2_1
XFILLER_31_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2753_ _2744_/X _2753_/A2 _1709_/X _1710_/X _2745_/X vssd1 vssd1 vccd1 vccd1 _3242_/D
+ sky130_fd_sc_hd__a221o_1
X_1704_ _1670_/X _3241_/Q _1671_/X vssd1 vssd1 vccd1 vccd1 _1704_/X sky130_fd_sc_hd__o21ba_1
X_2684_ _2712_/A vssd1 vssd1 vccd1 vccd1 _2684_/X sky130_fd_sc_hd__clkbuf_2
X_1635_ _1713_/A vssd1 vssd1 vccd1 vccd1 _1635_/X sky130_fd_sc_hd__clkbuf_2
X_1566_ _2675_/A vssd1 vssd1 vccd1 vccd1 _1566_/X sky130_fd_sc_hd__buf_4
XFILLER_86_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3305_ _3410_/CLK _3305_/D vssd1 vssd1 vccd1 vccd1 _3305_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1497_ _3180_/Q _1478_/X _1496_/Y vssd1 vssd1 vccd1 vccd1 _1497_/X sky130_fd_sc_hd__o21a_2
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _3258_/CLK _3236_/D vssd1 vssd1 vccd1 vccd1 _3236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3167_ _3482_/CLK _3167_/D vssd1 vssd1 vccd1 vccd1 _3167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2118_ _3346_/Q _2111_/X _2117_/Y vssd1 vssd1 vccd1 vccd1 _2118_/X sky130_fd_sc_hd__o21a_1
XFILLER_54_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3098_ _2106_/C _3091_/X _3095_/X _2421_/Y vssd1 vssd1 vccd1 vccd1 _3444_/D sky130_fd_sc_hd__o211ai_1
XFILLER_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2049_ _2049_/A vssd1 vssd1 vccd1 vccd1 _2081_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_54_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1827__A _2967_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2780__A2 _2779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2532__A2 _3138_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input142_A core_imem_request_put[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2296__A1 _1945_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2599__A2 _2599_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1737__A _1737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output459_A _1493_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1420_ _1426_/A vssd1 vssd1 vccd1 vccd1 _2675_/B sky130_fd_sc_hd__buf_2
XFILLER_79_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3021_ _3035_/A vssd1 vssd1 vccd1 vccd1 _3021_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2805_ _2805_/A _2818_/B vssd1 vssd1 vccd1 vccd1 _3271_/D sky130_fd_sc_hd__nand2_1
X_2736_ _1772_/X _2736_/A2 _1647_/X _1650_/X _2771_/A vssd1 vssd1 vccd1 vccd1 _3228_/D
+ sky130_fd_sc_hd__a221o_1
Xoutput510 _2286_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[35] sky130_fd_sc_hd__buf_2
X_2667_ _2667_/A _2673_/B vssd1 vssd1 vccd1 vccd1 _3184_/D sky130_fd_sc_hd__nand2_1
XANTENNA__2762__A2 _2762_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput554 _2400_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[75] sky130_fd_sc_hd__buf_2
Xoutput521 _2314_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[45] sky130_fd_sc_hd__buf_2
Xoutput532 _2343_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[55] sky130_fd_sc_hd__buf_2
Xoutput543 _2372_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[65] sky130_fd_sc_hd__buf_2
X_1618_ _2707_/A vssd1 vssd1 vccd1 vccd1 _1618_/X sky130_fd_sc_hd__clkbuf_4
Xoutput587 _1589_/X vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[14] sky130_fd_sc_hd__buf_2
Xoutput565 _2429_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[85] sky130_fd_sc_hd__buf_2
Xoutput576 _2453_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[95] sky130_fd_sc_hd__buf_2
X_2598_ _2598_/A _2473_/A vssd1 vssd1 vccd1 vccd1 _2598_/X sky130_fd_sc_hd__or2b_1
Xoutput598 _1617_/X vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[24] sky130_fd_sc_hd__buf_2
X_1549_ _1546_/X _1547_/X _1548_/X _1423_/C _1527_/A vssd1 vssd1 vccd1 vccd1 _1549_/Y
+ sky130_fd_sc_hd__o311ai_4
X_3219_ _3388_/CLK _3219_/D vssd1 vssd1 vccd1 vccd1 _3219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2738__C1 _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2202__A1 _1824_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2753__A2 _2753_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1467__A _1480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2521_ _2564_/A vssd1 vssd1 vccd1 vccd1 _2521_/X sky130_fd_sc_hd__clkbuf_2
X_2452_ _2225_/A _1801_/B _3456_/Q vssd1 vssd1 vccd1 vccd1 _2452_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2383_ _2459_/B vssd1 vssd1 vccd1 vccd1 _2383_/X sky130_fd_sc_hd__clkbuf_2
X_3004_ _3379_/Q _2993_/X _2233_/Y _3003_/X vssd1 vssd1 vccd1 vccd1 _3379_/D sky130_fd_sc_hd__o211a_1
XFILLER_49_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput3 EN_core_imem_request_put vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_4
XFILLER_36_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2983__A2 _2451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1808__C _1808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2719_ _1516_/C _2707_/X _2712_/X _1619_/Y vssd1 vssd1 vccd1 vccd1 _3219_/D sky130_fd_sc_hd__o211ai_1
XANTENNA_clkbuf_leaf_30_CLK_A clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput340 _1655_/Y vssd1 vssd1 vccd1 vccd1 core_imem_response_get[2] sky130_fd_sc_hd__buf_2
Xoutput351 _1837_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[10] sky130_fd_sc_hd__buf_2
Xoutput362 _1874_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[20] sky130_fd_sc_hd__buf_2
Xoutput395 _1987_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[50] sky130_fd_sc_hd__buf_2
Xoutput384 _1950_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[40] sky130_fd_sc_hd__buf_2
Xoutput373 _1914_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[30] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_45_CLK_A clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2936__A _2936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input105_A core_dmem_request_put[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input70_A core_dmem_request_put[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3151__A2 _3151_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1750__A _2765_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output324_A _1711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2581__A _2581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1952_ _1952_/A vssd1 vssd1 vccd1 vccd1 _1953_/C sky130_fd_sc_hd__inv_2
XFILLER_33_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1883_ _2031_/A vssd1 vssd1 vccd1 vccd1 _1917_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_2504_ _3131_/B vssd1 vssd1 vccd1 vccd1 _2504_/Y sky130_fd_sc_hd__inv_2
X_3484_ _3486_/CLK _3484_/D vssd1 vssd1 vccd1 vccd1 _3484_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2435_ _2412_/X _2413_/X _2414_/X _2124_/C _2434_/X vssd1 vssd1 vccd1 vccd1 _2435_/Y
+ sky130_fd_sc_hd__o311ai_4
XANTENNA__3142__A2 _3142_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2366_ _2033_/C _2340_/X _2365_/Y vssd1 vssd1 vccd1 vccd1 _2366_/Y sky130_fd_sc_hd__o21ai_2
X_2297_ _2326_/A vssd1 vssd1 vccd1 vccd1 _2297_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2491__A _2491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1695__A2 _2749_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input222_A ram_dmem_response_put[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1745__A _1745_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output441_A _2138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output539_A _2362_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2220_ _2196_/X _2206_/X _3374_/Q vssd1 vssd1 vccd1 vccd1 _2220_/Y sky130_fd_sc_hd__o21ai_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2151_ _2151_/A vssd1 vssd1 vccd1 vccd1 _2152_/C sky130_fd_sc_hd__inv_2
XANTENNA__1480__A _1480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1686__A2 _2746_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2082_ _3336_/Q _2075_/X _2081_/Y vssd1 vssd1 vccd1 vccd1 _2082_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2984_ _3365_/Q _2974_/X _2193_/Y _2978_/X vssd1 vssd1 vccd1 vccd1 _3365_/D sky130_fd_sc_hd__o211a_1
XFILLER_61_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1769__B_N _1644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3060__A1 _2011_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1935_ _1963_/A _1935_/B _1935_/C vssd1 vssd1 vccd1 vccd1 _1935_/Y sky130_fd_sc_hd__nand3_1
X_1866_ _1888_/A _1898_/B _1866_/C vssd1 vssd1 vccd1 vccd1 _1866_/Y sky130_fd_sc_hd__nand3_2
Xinput50 core_dmem_request_put[42] vssd1 vssd1 vccd1 vccd1 _1955_/A sky130_fd_sc_hd__clkbuf_1
X_1797_ _1951_/A vssd1 vssd1 vccd1 vccd1 _1832_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput61 core_dmem_request_put[52] vssd1 vssd1 vccd1 vccd1 _1992_/A sky130_fd_sc_hd__buf_2
Xinput72 core_dmem_request_put[62] vssd1 vssd1 vccd1 vccd1 _2028_/A sky130_fd_sc_hd__buf_2
Xinput94 core_dmem_request_put[82] vssd1 vssd1 vccd1 vccd1 _2101_/A sky130_fd_sc_hd__buf_2
Xinput83 core_dmem_request_put[72] vssd1 vssd1 vccd1 vccd1 _2064_/A sky130_fd_sc_hd__buf_2
XFILLER_1_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3467_ _3473_/CLK _3467_/D vssd1 vssd1 vccd1 vccd1 _3467_/Q sky130_fd_sc_hd__dfxtp_1
X_3398_ _3404_/CLK _3398_/D vssd1 vssd1 vccd1 vccd1 _3398_/Q sky130_fd_sc_hd__dfxtp_1
X_2418_ _2099_/C _2397_/X _2417_/Y vssd1 vssd1 vccd1 vccd1 _2418_/Y sky130_fd_sc_hd__o21ai_4
X_2349_ _2327_/X _2328_/X _2329_/X _2015_/C _2348_/X vssd1 vssd1 vccd1 vccd1 _2349_/Y
+ sky130_fd_sc_hd__o311ai_2
XFILLER_29_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1821__C _1821_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input172_A fmc_dmem_response_put[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3106__A2 _3105_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2099__C _2099_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input33_A core_dmem_request_put[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output391_A _1975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3042__A1 _1960_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1720_ _1720_/A _1684_/X vssd1 vssd1 vccd1 vccd1 _1720_/X sky130_fd_sc_hd__or2b_1
XFILLER_7_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1651_ _1642_/X _2736_/A2 _1647_/X _1650_/X vssd1 vssd1 vccd1 vccd1 _1651_/X sky130_fd_sc_hd__a22o_2
XANTENNA__1906__C _1906_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1582_ _1563_/X _1569_/X _3205_/Q vssd1 vssd1 vccd1 vccd1 _1582_/Y sky130_fd_sc_hd__o21ai_1
X_3321_ _3432_/CLK _3321_/D vssd1 vssd1 vccd1 vccd1 _3321_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _3252_/CLK _3252_/D vssd1 vssd1 vccd1 vccd1 _3252_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2305__B1 _1956_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2203_ _2291_/A vssd1 vssd1 vccd1 vccd1 _2203_/X sky130_fd_sc_hd__buf_2
X_3183_ _3404_/CLK _3183_/D vssd1 vssd1 vccd1 vccd1 _3183_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1659__A2 _2738_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2134_ _2169_/A _2134_/B _2134_/C vssd1 vssd1 vccd1 vccd1 _2134_/Y sky130_fd_sc_hd__nand3_1
XFILLER_54_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2065_ _2072_/A _2081_/B _2065_/C vssd1 vssd1 vccd1 vccd1 _2065_/Y sky130_fd_sc_hd__nand3_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2967_ _2967_/A _2967_/B vssd1 vssd1 vccd1 vccd1 _2969_/A sky130_fd_sc_hd__nand2_1
X_2898_ _2936_/A vssd1 vssd1 vccd1 vccd1 _2914_/B sky130_fd_sc_hd__clkbuf_2
X_1918_ _3291_/Q _1911_/X _1917_/Y vssd1 vssd1 vccd1 vccd1 _1918_/X sky130_fd_sc_hd__o21a_2
X_1849_ _1849_/A vssd1 vssd1 vccd1 vccd1 _1850_/C sky130_fd_sc_hd__inv_4
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput240 ram_dmem_response_put[8] vssd1 vssd1 vccd1 vccd1 _2509_/A sky130_fd_sc_hd__buf_2
Xinput251 ram_imem_response_put[18] vssd1 vssd1 vccd1 vccd1 _1723_/A sky130_fd_sc_hd__clkbuf_2
Xinput262 ram_imem_response_put[28] vssd1 vssd1 vccd1 vccd1 _1762_/A sky130_fd_sc_hd__buf_2
Xinput273 ram_imem_response_put[9] vssd1 vssd1 vccd1 vccd1 _1685_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output404_A _2019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2854__A _2893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2066__A2 _2056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3015__A1 _1894_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2821_ _2878_/A vssd1 vssd1 vccd1 vccd1 _2837_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2752_ _2756_/A _2752_/B vssd1 vssd1 vccd1 vccd1 _3241_/D sky130_fd_sc_hd__nor2_1
X_1703_ _1691_/X _2751_/A2 _1701_/X _1702_/X vssd1 vssd1 vccd1 vccd1 _1703_/X sky130_fd_sc_hd__a22o_1
X_2683_ _2686_/A vssd1 vssd1 vccd1 vccd1 _2712_/A sky130_fd_sc_hd__clkbuf_2
X_1634_ _1776_/B vssd1 vssd1 vccd1 vccd1 _1713_/A sky130_fd_sc_hd__clkbuf_2
X_1565_ _1443_/C _1562_/X _1564_/Y vssd1 vssd1 vccd1 vccd1 _1565_/Y sky130_fd_sc_hd__o21ai_2
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1933__A _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3304_ _3304_/CLK _3304_/D vssd1 vssd1 vccd1 vccd1 _3304_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3235_ _3472_/CLK _3235_/D vssd1 vssd1 vccd1 vccd1 _3235_/Q sky130_fd_sc_hd__dfxtp_1
X_1496_ _1516_/A _1523_/B _1496_/C vssd1 vssd1 vccd1 vccd1 _1496_/Y sky130_fd_sc_hd__nand3_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3166_ _3477_/CLK _3166_/D vssd1 vssd1 vccd1 vccd1 _3166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3097_ _3443_/Q _3093_/X _2419_/Y _3089_/X vssd1 vssd1 vccd1 vccd1 _3443_/D sky130_fd_sc_hd__o211a_1
X_2117_ _2143_/A _2117_/B _2117_/C vssd1 vssd1 vccd1 vccd1 _2117_/Y sky130_fd_sc_hd__nand3_1
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2048_ _3327_/Q _2038_/X _2047_/Y vssd1 vssd1 vccd1 vccd1 _2048_/X sky130_fd_sc_hd__o21a_2
XFILLER_22_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3006__A1 _1869_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input135_A core_imem_request_put[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2048__A2 _2038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1559__A1 _1435_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1456__C _1456_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2849__A _2868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output521_A _2314_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3020_ _3389_/Q _3007_/X _2263_/Y _3019_/X vssd1 vssd1 vccd1 vccd1 _3389_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2584__A _2584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2804_ _3271_/Q _2795_/X _1840_/Y vssd1 vssd1 vccd1 vccd1 _2805_/A sky130_fd_sc_hd__o21ai_1
X_2735_ _2760_/A vssd1 vssd1 vccd1 vccd1 _2771_/A sky130_fd_sc_hd__buf_2
Xoutput511 _2288_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[36] sky130_fd_sc_hd__buf_2
Xoutput500 _2259_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[26] sky130_fd_sc_hd__buf_2
X_2666_ _3184_/Q _1415_/A _1509_/Y vssd1 vssd1 vccd1 vccd1 _2667_/A sky130_fd_sc_hd__o21ai_1
Xoutput522 _2316_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[46] sky130_fd_sc_hd__buf_2
Xoutput533 _2345_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[56] sky130_fd_sc_hd__buf_2
Xoutput544 _2374_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[66] sky130_fd_sc_hd__buf_2
X_1617_ _3218_/Q _1604_/X _1616_/Y vssd1 vssd1 vccd1 vccd1 _1617_/X sky130_fd_sc_hd__o21a_1
Xoutput566 _2431_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[86] sky130_fd_sc_hd__buf_2
Xoutput577 _2455_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[96] sky130_fd_sc_hd__buf_2
Xoutput555 _2402_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[76] sky130_fd_sc_hd__buf_2
X_2597_ _2466_/X _3158_/Q _2541_/A vssd1 vssd1 vccd1 vccd1 _2597_/X sky130_fd_sc_hd__o21ba_1
Xoutput588 _1593_/Y vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[15] sky130_fd_sc_hd__buf_2
Xoutput599 _1620_/Y vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[25] sky130_fd_sc_hd__buf_2
X_1548_ _1607_/A vssd1 vssd1 vccd1 vccd1 _1548_/X sky130_fd_sc_hd__buf_4
X_1479_ _1479_/A vssd1 vssd1 vccd1 vccd1 _1480_/C sky130_fd_sc_hd__inv_2
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3218_ _3388_/CLK _3218_/D vssd1 vssd1 vccd1 vccd1 _3218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3149_ _3140_/X _3149_/A2 _2565_/X _2566_/X _3141_/X vssd1 vssd1 vccd1 vccd1 _3483_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_27_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_4_CLK_A clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1838__A _1951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input252_A ram_imem_response_put[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2441__A2 _2439_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1748__A _1748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output569_A _2438_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output471_A _1538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2520_ _2520_/A vssd1 vssd1 vccd1 vccd1 _2520_/X sky130_fd_sc_hd__clkbuf_2
X_2451_ _3091_/A vssd1 vssd1 vccd1 vccd1 _2451_/X sky130_fd_sc_hd__buf_4
XFILLER_5_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2382_ _2054_/C _2369_/X _2381_/Y vssd1 vssd1 vccd1 vccd1 _2382_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3003_ _3003_/A vssd1 vssd1 vccd1 vccd1 _3003_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput4 EN_core_imem_response_get vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2680__A2 _1514_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1658__A _1658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2718_ _3218_/Q _2709_/X _1616_/Y _2710_/X vssd1 vssd1 vccd1 vccd1 _3218_/D sky130_fd_sc_hd__o211a_1
XFILLER_10_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput330 _1733_/Y vssd1 vssd1 vccd1 vccd1 core_imem_response_get[20] sky130_fd_sc_hd__buf_2
Xoutput341 _1771_/Y vssd1 vssd1 vccd1 vccd1 core_imem_response_get[30] sky130_fd_sc_hd__buf_2
Xoutput352 _1841_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[11] sky130_fd_sc_hd__buf_2
X_2649_ _2649_/A _2655_/B vssd1 vssd1 vccd1 vccd1 _3174_/D sky130_fd_sc_hd__nand2_1
XFILLER_87_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput385 _1954_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[41] sky130_fd_sc_hd__buf_2
Xoutput396 _1991_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[51] sky130_fd_sc_hd__buf_2
Xoutput374 _1918_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[31] sky130_fd_sc_hd__buf_2
XANTENNA__1824__C _1824_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput363 _1878_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[21] sky130_fd_sc_hd__buf_2
XFILLER_19_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2187__A1 _2165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input63_A core_dmem_request_put[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1951_ _1951_/A vssd1 vssd1 vccd1 vccd1 _1981_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1909__C _1909_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1882_ _2235_/A vssd1 vssd1 vccd1 vccd1 _2031_/A sky130_fd_sc_hd__buf_2
X_2503_ _2498_/X _2503_/A2 _2501_/X _2502_/X vssd1 vssd1 vccd1 vccd1 _3131_/B sky130_fd_sc_hd__a22oi_4
X_3483_ _3485_/CLK _3483_/D vssd1 vssd1 vccd1 vccd1 _3483_/Q sky130_fd_sc_hd__dfxtp_1
X_2434_ _2434_/A vssd1 vssd1 vccd1 vccd1 _2434_/X sky130_fd_sc_hd__buf_4
XFILLER_69_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2365_ _2341_/X _2351_/X _3424_/Q vssd1 vssd1 vccd1 vccd1 _2365_/Y sky130_fd_sc_hd__o21ai_1
X_2296_ _1945_/C _2283_/X _2295_/Y vssd1 vssd1 vccd1 vccd1 _2296_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_56_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input215_A ram_dmem_response_put[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3018__A _3095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1464__C _1464_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2150_ _2291_/A vssd1 vssd1 vccd1 vccd1 _2152_/A sky130_fd_sc_hd__buf_4
XFILLER_66_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2081_ _2109_/A _2081_/B _2081_/C vssd1 vssd1 vccd1 vccd1 _2081_/Y sky130_fd_sc_hd__nand3_1
XANTENNA_output601_A _1624_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2983_ _1808_/C _2451_/X _2980_/X _2191_/Y vssd1 vssd1 vccd1 vccd1 _3364_/D sky130_fd_sc_hd__o211ai_1
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1934_ _1934_/A vssd1 vssd1 vccd1 vccd1 _1935_/C sky130_fd_sc_hd__clkinv_4
XANTENNA_clkbuf_leaf_44_CLK_A clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput40 core_dmem_request_put[33] vssd1 vssd1 vccd1 vccd1 _1923_/A sky130_fd_sc_hd__clkbuf_1
X_1865_ _1865_/A vssd1 vssd1 vccd1 vccd1 _1866_/C sky130_fd_sc_hd__inv_4
Xinput62 core_dmem_request_put[53] vssd1 vssd1 vccd1 vccd1 _1996_/A sky130_fd_sc_hd__clkbuf_1
Xinput51 core_dmem_request_put[43] vssd1 vssd1 vccd1 vccd1 _1959_/A sky130_fd_sc_hd__clkbuf_1
Xinput73 core_dmem_request_put[63] vssd1 vssd1 vccd1 vccd1 _2032_/A sky130_fd_sc_hd__clkbuf_1
X_1796_ _2319_/A vssd1 vssd1 vccd1 vccd1 _1951_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2166__A4 _2165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput84 core_dmem_request_put[73] vssd1 vssd1 vccd1 vccd1 _2068_/A sky130_fd_sc_hd__clkbuf_1
Xinput95 core_dmem_request_put[83] vssd1 vssd1 vccd1 vccd1 _2105_/A sky130_fd_sc_hd__clkbuf_1
X_3466_ _3466_/CLK _3466_/D vssd1 vssd1 vccd1 vccd1 _3466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2417_ _2398_/X _2408_/X _3442_/Q vssd1 vssd1 vccd1 vccd1 _2417_/Y sky130_fd_sc_hd__o21ai_2
X_3397_ _3397_/CLK _3397_/D vssd1 vssd1 vccd1 vccd1 _3397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2348_ _2434_/A vssd1 vssd1 vccd1 vccd1 _2348_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2279_ _1924_/C _2253_/X _2278_/Y vssd1 vssd1 vccd1 vccd1 _2279_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2007__A _2007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input165_A fmc_dmem_response_put[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2314__A1 _1967_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input26_A core_dmem_request_put[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output384_A _1950_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1650_ _1650_/A _1649_/X vssd1 vssd1 vccd1 vccd1 _1650_/X sky130_fd_sc_hd__or2b_1
X_1581_ _3204_/Q _1576_/X _1580_/Y vssd1 vssd1 vccd1 vccd1 _1581_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3320_ _3330_/CLK _3320_/D vssd1 vssd1 vccd1 vccd1 _3320_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3297_/CLK _3251_/D vssd1 vssd1 vccd1 vccd1 _3251_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2202_ _1824_/C _2195_/X _2201_/Y vssd1 vssd1 vccd1 vccd1 _2202_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3182_ _3244_/CLK _3182_/D vssd1 vssd1 vccd1 vccd1 _3182_/Q sky130_fd_sc_hd__dfxtp_1
X_2133_ _2133_/A vssd1 vssd1 vccd1 vccd1 _2134_/C sky130_fd_sc_hd__inv_2
XFILLER_93_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2064_ _2064_/A vssd1 vssd1 vccd1 vccd1 _2065_/C sky130_fd_sc_hd__inv_2
XFILLER_62_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2966_ _3356_/Q _2779_/X _2959_/X _2152_/Y vssd1 vssd1 vccd1 vccd1 _3356_/D sky130_fd_sc_hd__o211a_1
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1917_ _1945_/A _1917_/B _1917_/C vssd1 vssd1 vccd1 vccd1 _1917_/Y sky130_fd_sc_hd__nand3_1
XFILLER_30_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2897_ _3319_/Q _2893_/X _2018_/Y vssd1 vssd1 vccd1 vccd1 _2899_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__1666__A _1666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1848_ _3273_/Q _1834_/X _1847_/Y vssd1 vssd1 vccd1 vccd1 _1848_/X sky130_fd_sc_hd__o21a_1
X_1779_ _1789_/B vssd1 vssd1 vccd1 vccd1 _2177_/A sky130_fd_sc_hd__buf_4
XFILLER_89_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3449_ _3449_/CLK _3449_/D vssd1 vssd1 vccd1 vccd1 _3449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2497__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1832__C _1832_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1576__A _1630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput241 ram_dmem_response_put[9] vssd1 vssd1 vccd1 vccd1 _2514_/A sky130_fd_sc_hd__clkbuf_4
Xinput263 ram_imem_response_put[29] vssd1 vssd1 vccd1 vccd1 _1766_/A sky130_fd_sc_hd__clkbuf_4
Xinput230 ram_dmem_response_put[28] vssd1 vssd1 vccd1 vccd1 _2591_/A sky130_fd_sc_hd__buf_2
Xinput252 ram_imem_response_put[19] vssd1 vssd1 vccd1 vccd1 _1728_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output599_A _1620_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2820_ _3279_/Q _2816_/X _1869_/Y vssd1 vssd1 vccd1 vccd1 _2822_/A sky130_fd_sc_hd__o21ai_1
XFILLER_31_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2751_ _2744_/X _2751_/A2 _1701_/X _1702_/X _2745_/X vssd1 vssd1 vccd1 vccd1 _3240_/D
+ sky130_fd_sc_hd__a221o_1
X_2682_ _2723_/A _2682_/B vssd1 vssd1 vccd1 vccd1 _2686_/A sky130_fd_sc_hd__and2b_1
XANTENNA__1917__C _1917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1702_ _1702_/A _1684_/X vssd1 vssd1 vccd1 vccd1 _1702_/X sky130_fd_sc_hd__or2b_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1633_ _1641_/A vssd1 vssd1 vccd1 vccd1 _1633_/X sky130_fd_sc_hd__buf_2
X_1564_ _1563_/X _1527_/B _3199_/Q vssd1 vssd1 vccd1 vccd1 _1564_/Y sky130_fd_sc_hd__o21ai_1
X_1495_ _1495_/A vssd1 vssd1 vccd1 vccd1 _1496_/C sky130_fd_sc_hd__inv_2
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3303_ _3410_/CLK _3303_/D vssd1 vssd1 vccd1 vccd1 _3303_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _3241_/CLK _3234_/D vssd1 vssd1 vccd1 vccd1 _3234_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3165_ _3485_/CLK _3165_/D vssd1 vssd1 vccd1 vccd1 _3165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2116_ _2116_/A vssd1 vssd1 vccd1 vccd1 _2117_/C sky130_fd_sc_hd__inv_2
XFILLER_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3096_ _2099_/C _3091_/X _3095_/X _2417_/Y vssd1 vssd1 vccd1 vccd1 _3442_/D sky130_fd_sc_hd__o211ai_1
X_2047_ _2054_/A _2062_/B _2047_/C vssd1 vssd1 vccd1 vccd1 _2047_/Y sky130_fd_sc_hd__nand3_1
XFILLER_22_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2214__B1 _1836_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2949_ _3346_/Q _2945_/X _2941_/X _2117_/Y vssd1 vssd1 vccd1 vccd1 _3346_/D sky130_fd_sc_hd__o211a_1
XFILLER_89_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3116__A _3116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input128_A core_imem_request_put[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input93_A core_dmem_request_put[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output514_A _2296_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2444__B1 _2137_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_49_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3472_/CLK sky130_fd_sc_hd__clkbuf_16
X_2803_ _3270_/Q _2789_/X _2784_/X _1836_/Y vssd1 vssd1 vccd1 vccd1 _3270_/D sky130_fd_sc_hd__o211a_1
X_2734_ _2743_/A _2734_/B vssd1 vssd1 vccd1 vccd1 _3227_/D sky130_fd_sc_hd__nor2_1
Xoutput501 _2261_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[27] sky130_fd_sc_hd__buf_2
X_2665_ _3183_/Q _2660_/X _2661_/X _1506_/Y vssd1 vssd1 vccd1 vccd1 _3183_/D sky130_fd_sc_hd__o211a_1
Xoutput512 _2290_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[37] sky130_fd_sc_hd__buf_2
Xoutput523 _2318_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[47] sky130_fd_sc_hd__buf_2
Xoutput534 _2347_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[57] sky130_fd_sc_hd__buf_2
Xoutput545 _2376_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[67] sky130_fd_sc_hd__buf_2
X_1616_ _1605_/X _1606_/X _1607_/X _1512_/C _1594_/X vssd1 vssd1 vccd1 vccd1 _1616_/Y
+ sky130_fd_sc_hd__o311ai_4
X_2596_ _2563_/X _2613_/A2 _2594_/X _2595_/X vssd1 vssd1 vccd1 vccd1 _2596_/X sky130_fd_sc_hd__a22o_1
Xoutput578 _2456_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[97] sky130_fd_sc_hd__buf_2
Xoutput567 _2433_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[87] sky130_fd_sc_hd__buf_2
Xoutput556 _2404_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[77] sky130_fd_sc_hd__buf_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput589 _1596_/X vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[16] sky130_fd_sc_hd__buf_2
XFILLER_59_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1547_ _1606_/A vssd1 vssd1 vccd1 vccd1 _1547_/X sky130_fd_sc_hd__buf_4
XFILLER_86_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1478_ _1514_/A vssd1 vssd1 vccd1 vccd1 _1478_/X sky130_fd_sc_hd__clkbuf_2
X_3217_ _3388_/CLK _3217_/D vssd1 vssd1 vccd1 vccd1 _3217_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2775__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3148_ _3152_/A _3148_/B vssd1 vssd1 vccd1 vccd1 _3482_/D sky130_fd_sc_hd__nor2_1
XFILLER_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3079_ _3093_/A vssd1 vssd1 vccd1 vccd1 _3079_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2199__C1 _2152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input245_A ram_imem_response_put[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2729__A1 _2725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1467__C _1467_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2450_ _3105_/A vssd1 vssd1 vccd1 vccd1 _3091_/A sky130_fd_sc_hd__buf_2
XFILLER_5_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2381_ _2370_/X _2380_/X _3430_/Q vssd1 vssd1 vccd1 vccd1 _2381_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__2595__A _2595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3002_ _1862_/C _2991_/X _2995_/X _2230_/Y vssd1 vssd1 vccd1 vccd1 _3378_/D sky130_fd_sc_hd__o211ai_1
Xinput5 EN_fmc_dmem_request_get vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2717_ _1509_/C _2707_/X _2712_/X _1614_/Y vssd1 vssd1 vccd1 vccd1 _3217_/D sky130_fd_sc_hd__o211ai_1
Xoutput331 _1738_/X vssd1 vssd1 vccd1 vccd1 core_imem_response_get[21] sky130_fd_sc_hd__buf_2
Xoutput342 _1775_/X vssd1 vssd1 vccd1 vccd1 core_imem_response_get[31] sky130_fd_sc_hd__buf_2
Xoutput320 _1695_/X vssd1 vssd1 vccd1 vccd1 core_imem_response_get[11] sky130_fd_sc_hd__buf_2
X_2648_ _3174_/Q _2644_/X _1473_/Y vssd1 vssd1 vccd1 vccd1 _2649_/A sky130_fd_sc_hd__o21ai_1
Xoutput353 _1844_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[12] sky130_fd_sc_hd__buf_2
Xoutput386 _1957_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[42] sky130_fd_sc_hd__buf_2
Xoutput375 _1921_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[32] sky130_fd_sc_hd__buf_2
X_2579_ _3152_/B vssd1 vssd1 vccd1 vccd1 _2579_/Y sky130_fd_sc_hd__inv_2
Xoutput364 _1881_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[22] sky130_fd_sc_hd__buf_2
Xoutput397 _1994_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[52] sky130_fd_sc_hd__buf_2
XFILLER_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1840__C _1840_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input195_A fmc_imem_response_put[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2187__A2 _2186_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input56_A core_dmem_request_put[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1759__A _1759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1950_ _3300_/Q _1947_/X _1949_/Y vssd1 vssd1 vccd1 vccd1 _1950_/X sky130_fd_sc_hd__o21a_2
X_1881_ _3282_/Q _1871_/X _1880_/Y vssd1 vssd1 vccd1 vccd1 _1881_/X sky130_fd_sc_hd__o21a_1
X_2502_ _2502_/A _2490_/X vssd1 vssd1 vccd1 vccd1 _2502_/X sky130_fd_sc_hd__or2b_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3482_ _3482_/CLK _3482_/D vssd1 vssd1 vccd1 vccd1 _3482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_3_CLK_A clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2433_ _2120_/C _2426_/X _2432_/Y vssd1 vssd1 vccd1 vccd1 _2433_/Y sky130_fd_sc_hd__o21ai_4
X_2364_ _3423_/Q _2355_/X _2363_/Y vssd1 vssd1 vccd1 vccd1 _2364_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2295_ _2284_/X _2294_/X _3400_/Q vssd1 vssd1 vccd1 vccd1 _2295_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_56_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3118__A1 _2225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3124__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input110_A core_dmem_request_put[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input208_A fmc_imem_response_put[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2682__B _2682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2080_ _2080_/A vssd1 vssd1 vccd1 vccd1 _2081_/C sky130_fd_sc_hd__inv_2
XANTENNA__1480__C _1480_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2873__A _2893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2982_ _3363_/Q _2974_/X _2189_/Y _2978_/X vssd1 vssd1 vccd1 vccd1 _3363_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1933_ _2006_/A vssd1 vssd1 vccd1 vccd1 _1963_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput30 core_dmem_request_put[24] vssd1 vssd1 vccd1 vccd1 _1887_/A sky130_fd_sc_hd__clkbuf_1
X_1864_ _2967_/B vssd1 vssd1 vccd1 vccd1 _1898_/B sky130_fd_sc_hd__clkbuf_2
Xinput52 core_dmem_request_put[44] vssd1 vssd1 vccd1 vccd1 _1962_/A sky130_fd_sc_hd__clkbuf_1
Xinput41 core_dmem_request_put[34] vssd1 vssd1 vccd1 vccd1 _1926_/A sky130_fd_sc_hd__clkbuf_1
Xinput63 core_dmem_request_put[54] vssd1 vssd1 vccd1 vccd1 _1999_/A sky130_fd_sc_hd__buf_2
X_1795_ _3260_/Q _1784_/X _1794_/Y vssd1 vssd1 vccd1 vccd1 _1795_/X sky130_fd_sc_hd__o21a_1
Xinput96 core_dmem_request_put[84] vssd1 vssd1 vccd1 vccd1 _2108_/A sky130_fd_sc_hd__buf_2
Xinput85 core_dmem_request_put[74] vssd1 vssd1 vccd1 vccd1 _2071_/A sky130_fd_sc_hd__buf_2
Xinput74 core_dmem_request_put[64] vssd1 vssd1 vccd1 vccd1 _2035_/A sky130_fd_sc_hd__buf_2
XFILLER_6_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3465_ _3473_/CLK _3465_/D vssd1 vssd1 vccd1 vccd1 _3465_/Q sky130_fd_sc_hd__dfxtp_1
X_2416_ _3441_/Q _2411_/X _2415_/Y vssd1 vssd1 vccd1 vccd1 _2416_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3396_ _3404_/CLK _3396_/D vssd1 vssd1 vccd1 vccd1 _3396_/Q sky130_fd_sc_hd__dfxtp_1
X_2347_ _2011_/C _2340_/X _2346_/Y vssd1 vssd1 vccd1 vccd1 _2347_/Y sky130_fd_sc_hd__o21ai_2
X_2278_ _2255_/X _2265_/X _3394_/Q vssd1 vssd1 vccd1 vccd1 _2278_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2783__A _2959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input158_A fmc_dmem_response_put[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2677__B _2677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input19_A core_dmem_request_put[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2250__A1 _1885_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output377_A _1928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1580_ _1577_/X _1578_/X _1579_/X _1464_/C _1566_/X vssd1 vssd1 vccd1 vccd1 _1580_/Y
+ sky130_fd_sc_hd__o311ai_4
XANTENNA__2553__A2 _2553_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2868__A _2868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3252_/CLK _3250_/D vssd1 vssd1 vccd1 vccd1 _3250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2201_ _2196_/X _2186_/X _3368_/Q vssd1 vssd1 vccd1 vccd1 _2201_/Y sky130_fd_sc_hd__o21ai_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _3252_/CLK _3181_/D vssd1 vssd1 vccd1 vccd1 _3181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2132_ _3350_/Q _2129_/X _2131_/Y vssd1 vssd1 vccd1 vccd1 _2132_/X sky130_fd_sc_hd__o21a_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2063_ _3331_/Q _2056_/X _2062_/Y vssd1 vssd1 vccd1 vccd1 _2063_/X sky130_fd_sc_hd__o21a_2
XFILLER_62_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2108__A _2108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2965_ _2965_/A _2965_/B vssd1 vssd1 vccd1 vccd1 _3355_/D sky130_fd_sc_hd__nand2_1
X_2896_ _3318_/Q _2888_/X _2884_/X _2015_/Y vssd1 vssd1 vccd1 vccd1 _3318_/D sky130_fd_sc_hd__o211a_1
X_1916_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1917_/C sky130_fd_sc_hd__inv_2
X_1847_ _1869_/A _1877_/B _1847_/C vssd1 vssd1 vccd1 vccd1 _1847_/Y sky130_fd_sc_hd__nand3_1
X_1778_ _1789_/A vssd1 vssd1 vccd1 vccd1 _2175_/A sky130_fd_sc_hd__buf_4
X_3448_ _3448_/CLK _3448_/D vssd1 vssd1 vccd1 vccd1 _3448_/Q sky130_fd_sc_hd__dfxtp_1
X_3379_ _3397_/CLK _3379_/D vssd1 vssd1 vccd1 vccd1 _3379_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1857__A _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput220 ram_dmem_response_put[19] vssd1 vssd1 vccd1 vccd1 _2557_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput231 ram_dmem_response_put[29] vssd1 vssd1 vccd1 vccd1 _2595_/A sky130_fd_sc_hd__clkbuf_4
Xinput253 ram_imem_response_put[1] vssd1 vssd1 vccd1 vccd1 _1650_/A sky130_fd_sc_hd__clkbuf_2
Xinput242 ram_imem_response_put[0] vssd1 vssd1 vccd1 vccd1 _1638_/A sky130_fd_sc_hd__buf_2
XFILLER_0_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_43_CLK_A clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput264 ram_imem_response_put[2] vssd1 vssd1 vccd1 vccd1 _1653_/A sky130_fd_sc_hd__buf_2
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2750_ _2756_/A _2750_/B vssd1 vssd1 vccd1 vccd1 _3239_/D sky130_fd_sc_hd__nor2_1
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2681_ _2709_/A vssd1 vssd1 vccd1 vccd1 _2681_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1701_ _1692_/X _3240_/Q _1700_/X vssd1 vssd1 vccd1 vccd1 _1701_/X sky130_fd_sc_hd__o21ba_1
XFILLER_8_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1632_ input8/X vssd1 vssd1 vccd1 vccd1 _1641_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1563_ _1563_/A vssd1 vssd1 vccd1 vccd1 _1563_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2598__A _2598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3302_ _3432_/CLK _3302_/D vssd1 vssd1 vccd1 vccd1 _3302_/Q sky130_fd_sc_hd__dfxtp_1
X_1494_ _1597_/A vssd1 vssd1 vccd1 vccd1 _1523_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_79_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _3472_/CLK _3233_/D vssd1 vssd1 vccd1 vccd1 _3233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3164_ _3485_/CLK _3164_/D vssd1 vssd1 vccd1 vccd1 _3164_/Q sky130_fd_sc_hd__dfxtp_1
X_2115_ _2967_/A vssd1 vssd1 vccd1 vccd1 _2143_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3095_ _3095_/A vssd1 vssd1 vccd1 vccd1 _3095_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2046_ _2046_/A vssd1 vssd1 vccd1 vccd1 _2047_/C sky130_fd_sc_hd__inv_2
XFILLER_35_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1677__A _1677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2948_ _2948_/A _2952_/B vssd1 vssd1 vccd1 vccd1 _3345_/D sky130_fd_sc_hd__nand2_1
XFILLER_13_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2879_ _2879_/A _2895_/B vssd1 vssd1 vccd1 vccd1 _3309_/D sky130_fd_sc_hd__nand2_1
XANTENNA__2004__C _2004_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1843__C _1843_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2955__B _2965_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input86_A core_dmem_request_put[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2802_ _2802_/A _2818_/B vssd1 vssd1 vccd1 vccd1 _3269_/D sky130_fd_sc_hd__nand2_1
X_2733_ _2747_/A vssd1 vssd1 vccd1 vccd1 _2743_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput502 _2264_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[28] sky130_fd_sc_hd__buf_2
X_2664_ _2664_/A _2673_/B vssd1 vssd1 vccd1 vccd1 _3182_/D sky130_fd_sc_hd__nand2_1
Xoutput513 _2293_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[38] sky130_fd_sc_hd__buf_2
Xoutput524 _2322_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[48] sky130_fd_sc_hd__buf_2
Xoutput535 _2350_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[58] sky130_fd_sc_hd__buf_2
X_1615_ _1509_/C _1590_/X _1614_/Y vssd1 vssd1 vccd1 vccd1 _1615_/Y sky130_fd_sc_hd__o21ai_2
X_2595_ _2595_/A _2464_/X vssd1 vssd1 vccd1 vccd1 _2595_/X sky130_fd_sc_hd__or2b_1
Xoutput568 _2436_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[88] sky130_fd_sc_hd__buf_2
Xoutput546 _2379_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[68] sky130_fd_sc_hd__buf_2
Xoutput557 _2407_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[78] sky130_fd_sc_hd__buf_2
X_1546_ _1605_/A vssd1 vssd1 vccd1 vccd1 _1546_/X sky130_fd_sc_hd__buf_4
Xoutput579 _2457_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[98] sky130_fd_sc_hd__buf_2
X_1477_ _3175_/Q _1462_/X _1476_/Y vssd1 vssd1 vccd1 vccd1 _1477_/X sky130_fd_sc_hd__o21a_2
XFILLER_67_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3216_ _3222_/CLK _3216_/D vssd1 vssd1 vccd1 vccd1 _3216_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3147_ _3140_/X _3147_/A2 _2555_/X _2557_/X _3141_/X vssd1 vssd1 vccd1 vccd1 _3481_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3078_ _2054_/C _3077_/X _3067_/X _2381_/Y vssd1 vssd1 vccd1 vccd1 _3430_/D sky130_fd_sc_hd__o211ai_1
XFILLER_82_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2029_ _2036_/A _2044_/B _2029_/C vssd1 vssd1 vccd1 vccd1 _2029_/Y sky130_fd_sc_hd__nand3_1
XFILLER_24_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2199__B1 _1821_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2738__A2 _2738_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input238_A ram_dmem_response_put[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input140_A core_imem_request_put[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2206__A _2206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output457_A _1485_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2380_ _2408_/A vssd1 vssd1 vccd1 vccd1 _2380_/X sky130_fd_sc_hd__buf_2
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3001_ _3377_/Q _2993_/X _2228_/Y _2989_/X vssd1 vssd1 vccd1 vccd1 _3377_/D sky130_fd_sc_hd__o211a_1
XFILLER_49_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput6 EN_fmc_dmem_response_put vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_4
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1625__C1 _1443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2116__A _2116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2716_ _3216_/Q _2709_/X _1612_/Y _2710_/X vssd1 vssd1 vccd1 vccd1 _3216_/D sky130_fd_sc_hd__o211a_1
Xoutput310 _2604_/X vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[31] sky130_fd_sc_hd__buf_2
X_2647_ _3173_/Q _2641_/X _2642_/X _1470_/Y vssd1 vssd1 vccd1 vccd1 _3173_/D sky130_fd_sc_hd__o211a_1
Xoutput343 _1659_/X vssd1 vssd1 vccd1 vccd1 core_imem_response_get[3] sky130_fd_sc_hd__buf_2
Xoutput321 _1699_/Y vssd1 vssd1 vccd1 vccd1 core_imem_response_get[12] sky130_fd_sc_hd__buf_2
Xoutput332 _1742_/Y vssd1 vssd1 vccd1 vccd1 core_imem_response_get[22] sky130_fd_sc_hd__buf_2
XANTENNA__3145__A2 _3145_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput387 _1961_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[43] sky130_fd_sc_hd__buf_2
Xoutput376 _1925_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[33] sky130_fd_sc_hd__buf_2
X_2578_ _2541_/X _2578_/A2 _2576_/X _2577_/X vssd1 vssd1 vccd1 vccd1 _3152_/B sky130_fd_sc_hd__a22oi_4
Xoutput354 _1848_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[13] sky130_fd_sc_hd__buf_2
Xoutput365 _1886_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[23] sky130_fd_sc_hd__buf_2
XFILLER_87_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput398 _1998_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[53] sky130_fd_sc_hd__buf_2
X_1529_ _1529_/A vssd1 vssd1 vccd1 vccd1 _1605_/A sky130_fd_sc_hd__buf_2
XFILLER_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input188_A fmc_imem_response_put[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3136__A2 _3136_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1698__A2 _1698_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input49_A core_dmem_request_put[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3072__A1 _2040_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1880_ _1888_/A _1898_/B _1880_/C vssd1 vssd1 vccd1 vccd1 _1880_/Y sky130_fd_sc_hd__nand3_1
XANTENNA_output574_A _2447_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2501_ _2499_/X _3468_/Q _2500_/X vssd1 vssd1 vccd1 vccd1 _2501_/X sky130_fd_sc_hd__o21ba_1
X_3481_ _3485_/CLK _3481_/D vssd1 vssd1 vccd1 vccd1 _3481_/Q sky130_fd_sc_hd__dfxtp_1
X_2432_ _2427_/X _2408_/X _3448_/Q vssd1 vssd1 vccd1 vccd1 _2432_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2363_ _2356_/X _2357_/X _2358_/X _2029_/C _2348_/X vssd1 vssd1 vccd1 vccd1 _2363_/Y
+ sky130_fd_sc_hd__o311ai_4
XANTENNA__1689__A2 _1689_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2294_ _2351_/A vssd1 vssd1 vccd1 vccd1 _2294_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1685__A _1685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3118__A2 _2186_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input103_A core_dmem_request_put[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3054__A1 _1990_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3109__A2 _2174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output322_A _1703_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2096__A2 _2093_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2981_ _1801_/C _2451_/X _2980_/X _2187_/Y vssd1 vssd1 vccd1 vccd1 _3362_/D sky130_fd_sc_hd__o211ai_1
X_1932_ _3295_/Q _1929_/X _1931_/Y vssd1 vssd1 vccd1 vccd1 _1932_/X sky130_fd_sc_hd__o21a_2
X_1863_ _3277_/Q _1852_/X _1862_/Y vssd1 vssd1 vccd1 vccd1 _1863_/X sky130_fd_sc_hd__o21a_2
Xinput20 core_dmem_request_put[15] vssd1 vssd1 vccd1 vccd1 _1853_/A sky130_fd_sc_hd__clkbuf_1
Xinput31 core_dmem_request_put[25] vssd1 vssd1 vccd1 vccd1 _1893_/A sky130_fd_sc_hd__clkbuf_1
Xinput53 core_dmem_request_put[45] vssd1 vssd1 vccd1 vccd1 _1966_/A sky130_fd_sc_hd__clkbuf_1
Xinput42 core_dmem_request_put[35] vssd1 vssd1 vccd1 vccd1 _1930_/A sky130_fd_sc_hd__clkbuf_1
X_1794_ _3116_/A _1821_/B _1794_/C vssd1 vssd1 vccd1 vccd1 _1794_/Y sky130_fd_sc_hd__nand3_2
Xinput64 core_dmem_request_put[55] vssd1 vssd1 vccd1 vccd1 _2003_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_0_CLK_A CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput97 core_dmem_request_put[85] vssd1 vssd1 vccd1 vccd1 _2112_/A sky130_fd_sc_hd__clkbuf_2
Xinput86 core_dmem_request_put[75] vssd1 vssd1 vccd1 vccd1 _2076_/A sky130_fd_sc_hd__clkbuf_1
Xinput75 core_dmem_request_put[65] vssd1 vssd1 vccd1 vccd1 _2039_/A sky130_fd_sc_hd__clkbuf_1
X_3464_ _3466_/CLK _3464_/D vssd1 vssd1 vccd1 vccd1 _3464_/Q sky130_fd_sc_hd__dfxtp_1
X_2415_ _2412_/X _2413_/X _2414_/X _2095_/C _2405_/X vssd1 vssd1 vccd1 vccd1 _2415_/Y
+ sky130_fd_sc_hd__o311ai_4
X_3395_ _3459_/CLK _3395_/D vssd1 vssd1 vccd1 vccd1 _3395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2346_ _2341_/X _2323_/X _3418_/Q vssd1 vssd1 vccd1 vccd1 _2346_/Y sky130_fd_sc_hd__o21ai_1
X_2277_ _3393_/Q _2268_/X _2276_/Y vssd1 vssd1 vccd1 vccd1 _2277_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3036__A1 _1945_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2958__B _2965_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1770__A1 _1691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input220_A ram_dmem_response_put[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2078__A2 _2075_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_2_CLK_A clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1761__A1 _1637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2200_ _3367_/Q _2174_/X _2199_/Y vssd1 vssd1 vccd1 vccd1 _2200_/X sky130_fd_sc_hd__o21a_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3180_ _3244_/CLK _3180_/D vssd1 vssd1 vccd1 vccd1 _3180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2131_ _2143_/A _2152_/B _2131_/C vssd1 vssd1 vccd1 vccd1 _2131_/Y sky130_fd_sc_hd__nand3_1
X_2062_ _2091_/A _2062_/B _2062_/C vssd1 vssd1 vccd1 vccd1 _2062_/Y sky130_fd_sc_hd__nand3_1
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2964_ _3355_/Q _2950_/X _2147_/Y vssd1 vssd1 vccd1 vccd1 _2965_/A sky130_fd_sc_hd__o21ai_1
X_1915_ _1951_/A vssd1 vssd1 vccd1 vccd1 _1945_/A sky130_fd_sc_hd__clkbuf_2
X_2895_ _2895_/A _2895_/B vssd1 vssd1 vccd1 vccd1 _3317_/D sky130_fd_sc_hd__nand2_1
X_1846_ _1846_/A vssd1 vssd1 vccd1 vccd1 _1847_/C sky130_fd_sc_hd__inv_4
XFILLER_30_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1777_ _1777_/A vssd1 vssd1 vccd1 vccd1 _2773_/B sky130_fd_sc_hd__clkbuf_2
X_3447_ _3447_/CLK _3447_/D vssd1 vssd1 vccd1 vccd1 _3447_/Q sky130_fd_sc_hd__dfxtp_1
X_3378_ _3384_/CLK _3378_/D vssd1 vssd1 vccd1 vccd1 _3378_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2329_ _2414_/A vssd1 vssd1 vccd1 vccd1 _2329_/X sky130_fd_sc_hd__clkbuf_4
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2794__A _2794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2480__A2 _3123_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input170_A fmc_dmem_response_put[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input268_A ram_imem_response_put[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput210 ram_dmem_response_put[0] vssd1 vssd1 vccd1 vccd1 _2467_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput232 ram_dmem_response_put[2] vssd1 vssd1 vccd1 vccd1 _2482_/A sky130_fd_sc_hd__buf_2
Xinput221 ram_dmem_response_put[1] vssd1 vssd1 vccd1 vccd1 _2479_/A sky130_fd_sc_hd__clkbuf_4
Xinput243 ram_imem_response_put[10] vssd1 vssd1 vccd1 vccd1 _1688_/A sky130_fd_sc_hd__buf_2
Xinput254 ram_imem_response_put[20] vssd1 vssd1 vccd1 vccd1 _1731_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input31_A core_dmem_request_put[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput265 ram_imem_response_put[30] vssd1 vssd1 vccd1 vccd1 _1769_/A sky130_fd_sc_hd__buf_2
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2680_ _3193_/Q _1514_/X _2636_/B vssd1 vssd1 vccd1 vccd1 _3193_/D sky130_fd_sc_hd__o21a_1
X_1700_ _1743_/A vssd1 vssd1 vccd1 vccd1 _1700_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1631_ _1631_/A vssd1 vssd1 vccd1 vccd1 _1631_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1783__A _2950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1562_ _1562_/A vssd1 vssd1 vccd1 vccd1 _1562_/X sky130_fd_sc_hd__buf_2
X_3301_ _3410_/CLK _3301_/D vssd1 vssd1 vccd1 vccd1 _3301_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1493_ _3179_/Q _1478_/X _1492_/Y vssd1 vssd1 vccd1 vccd1 _1493_/X sky130_fd_sc_hd__o21a_2
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ _3472_/CLK _3232_/D vssd1 vssd1 vccd1 vccd1 _3232_/Q sky130_fd_sc_hd__dfxtp_1
X_3163_ _3482_/CLK _3163_/D vssd1 vssd1 vccd1 vccd1 _3163_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2114_ _3345_/Q _2111_/X _2113_/Y vssd1 vssd1 vccd1 vccd1 _2114_/X sky130_fd_sc_hd__o21a_2
XFILLER_94_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3094_ _3441_/Q _3093_/X _2415_/Y _3089_/X vssd1 vssd1 vccd1 vccd1 _3441_/D sky130_fd_sc_hd__o211a_1
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2045_ _3326_/Q _2038_/X _2044_/Y vssd1 vssd1 vccd1 vccd1 _2045_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2947_ _3345_/Q _2931_/X _2113_/Y vssd1 vssd1 vccd1 vccd1 _2948_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__2789__A _2868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2878_ _2878_/A vssd1 vssd1 vccd1 vccd1 _2895_/B sky130_fd_sc_hd__clkbuf_2
X_1829_ _1850_/A _1859_/B _1829_/C vssd1 vssd1 vccd1 vccd1 _1829_/Y sky130_fd_sc_hd__nand3_2
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2453__A2 _2451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input79_A core_dmem_request_put[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output402_A _2012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2801_ _2878_/A vssd1 vssd1 vccd1 vccd1 _2818_/B sky130_fd_sc_hd__clkbuf_2
X_2732_ _2760_/A vssd1 vssd1 vccd1 vccd1 _2747_/A sky130_fd_sc_hd__buf_2
XFILLER_8_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2663_ _3182_/Q _1415_/A _1503_/Y vssd1 vssd1 vccd1 vccd1 _2664_/A sky130_fd_sc_hd__o21ai_1
Xoutput503 _2267_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[29] sky130_fd_sc_hd__buf_2
Xoutput514 _2296_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[39] sky130_fd_sc_hd__buf_2
Xoutput525 _2325_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[49] sky130_fd_sc_hd__buf_2
Xoutput536 _2353_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[59] sky130_fd_sc_hd__buf_2
X_1614_ _1591_/X _1597_/X _3217_/Q vssd1 vssd1 vccd1 vccd1 _1614_/Y sky130_fd_sc_hd__o21ai_1
X_2594_ _2564_/X _3157_/Q _2572_/X vssd1 vssd1 vccd1 vccd1 _2594_/X sky130_fd_sc_hd__o21ba_1
Xoutput558 _2410_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[79] sky130_fd_sc_hd__buf_2
Xoutput569 _2438_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[89] sky130_fd_sc_hd__buf_2
Xoutput547 _2382_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[69] sky130_fd_sc_hd__buf_2
X_1545_ _1630_/B vssd1 vssd1 vccd1 vccd1 _1545_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3215_ _3388_/CLK _3215_/D vssd1 vssd1 vccd1 vccd1 _3215_/Q sky130_fd_sc_hd__dfxtp_1
X_1476_ _1476_/A _1484_/B _1476_/C vssd1 vssd1 vccd1 vccd1 _1476_/Y sky130_fd_sc_hd__nand3_1
X_3146_ _3152_/A _3146_/B vssd1 vssd1 vccd1 vccd1 _3480_/D sky130_fd_sc_hd__nor2_1
X_3077_ _3091_/A vssd1 vssd1 vccd1 vccd1 _3077_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2028_ _2028_/A vssd1 vssd1 vccd1 vccd1 _2029_/C sky130_fd_sc_hd__clkinv_2
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1688__A _1688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_42_CLK_A clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2312__A _2370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1854__C _1854_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input133_A core_imem_request_put[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2362__A1 _2026_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3053__A _3067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3000_ _1854_/C _2991_/X _2995_/X _2226_/Y vssd1 vssd1 vccd1 vccd1 _3376_/D sky130_fd_sc_hd__o211ai_1
XFILLER_49_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 EN_fmc_imem_request_get vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_2
XFILLER_64_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1625__B1 _1527_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2715_ _1503_/C _2707_/X _2712_/X _1610_/Y vssd1 vssd1 vccd1 vccd1 _3215_/D sky130_fd_sc_hd__o211ai_1
Xoutput300 _2571_/Y vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[22] sky130_fd_sc_hd__buf_2
X_2646_ _2646_/A _2655_/B vssd1 vssd1 vccd1 vccd1 _3172_/D sky130_fd_sc_hd__nand2_1
Xoutput344 _1664_/Y vssd1 vssd1 vccd1 vccd1 core_imem_response_get[4] sky130_fd_sc_hd__buf_2
Xoutput322 _1703_/X vssd1 vssd1 vccd1 vccd1 core_imem_response_get[13] sky130_fd_sc_hd__buf_2
Xoutput311 _2488_/X vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[3] sky130_fd_sc_hd__buf_2
Xoutput333 _1746_/X vssd1 vssd1 vccd1 vccd1 core_imem_response_get[23] sky130_fd_sc_hd__buf_2
Xoutput377 _1928_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[34] sky130_fd_sc_hd__buf_2
X_2577_ _2577_/A _2473_/A vssd1 vssd1 vccd1 vccd1 _2577_/X sky130_fd_sc_hd__or2b_1
Xoutput355 _1851_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[14] sky130_fd_sc_hd__buf_2
Xoutput366 _1889_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[24] sky130_fd_sc_hd__buf_2
Xoutput399 _2001_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[54] sky130_fd_sc_hd__buf_2
Xoutput388 _1964_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[44] sky130_fd_sc_hd__buf_2
X_1528_ _3189_/Q _1514_/X _1527_/Y vssd1 vssd1 vccd1 vccd1 _1528_/X sky130_fd_sc_hd__o21a_2
X_1459_ _1459_/A vssd1 vssd1 vccd1 vccd1 _1460_/C sky130_fd_sc_hd__clkinv_4
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3129_ _3127_/X _3129_/A2 _2494_/X _2495_/X _3128_/X vssd1 vssd1 vccd1 vccd1 _3467_/D
+ sky130_fd_sc_hd__a221o_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1616__B1 _1512_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2592__A1 _2520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2977__A _3095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input250_A ram_imem_response_put[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_3_0_CLK_A clkbuf_2_3_0_CLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2280__B1 _1927_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output567_A _2433_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2583__A1 _2466_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2500_ _2572_/A vssd1 vssd1 vccd1 vccd1 _2500_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3480_ _3482_/CLK _3480_/D vssd1 vssd1 vccd1 vccd1 _3480_/Q sky130_fd_sc_hd__dfxtp_1
X_2431_ _3447_/Q _2411_/X _2430_/Y vssd1 vssd1 vccd1 vccd1 _2431_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2362_ _2026_/C _2340_/X _2361_/Y vssd1 vssd1 vccd1 vccd1 _2362_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2293_ _3399_/Q _2268_/X _2292_/Y vssd1 vssd1 vccd1 vccd1 _2293_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2629_ _3164_/Q _2623_/X _1435_/Y vssd1 vssd1 vccd1 vccd1 _2630_/A sky130_fd_sc_hd__o21ai_1
XFILLER_87_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1837__B1 _1836_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input61_A core_dmem_request_put[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2980_ _3103_/A vssd1 vssd1 vccd1 vccd1 _2980_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1931_ _1945_/A _1953_/B _1931_/C vssd1 vssd1 vccd1 vccd1 _1931_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__1786__A _2163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1862_ _1869_/A _1877_/B _1862_/C vssd1 vssd1 vccd1 vccd1 _1862_/Y sky130_fd_sc_hd__nand3_1
Xinput10 EN_ram_dmem_response_put vssd1 vssd1 vccd1 vccd1 _2605_/B sky130_fd_sc_hd__buf_4
Xinput21 core_dmem_request_put[16] vssd1 vssd1 vccd1 vccd1 _1858_/A sky130_fd_sc_hd__clkbuf_1
Xinput32 core_dmem_request_put[26] vssd1 vssd1 vccd1 vccd1 _1897_/A sky130_fd_sc_hd__clkbuf_1
Xinput43 core_dmem_request_put[36] vssd1 vssd1 vccd1 vccd1 _1934_/A sky130_fd_sc_hd__clkbuf_1
Xinput54 core_dmem_request_put[46] vssd1 vssd1 vccd1 vccd1 _1970_/A sky130_fd_sc_hd__buf_2
X_1793_ _1793_/A vssd1 vssd1 vccd1 vccd1 _1794_/C sky130_fd_sc_hd__inv_6
Xinput98 core_dmem_request_put[86] vssd1 vssd1 vccd1 vccd1 _2116_/A sky130_fd_sc_hd__buf_2
Xinput87 core_dmem_request_put[76] vssd1 vssd1 vccd1 vccd1 _2080_/A sky130_fd_sc_hd__buf_2
Xinput65 core_dmem_request_put[56] vssd1 vssd1 vccd1 vccd1 _2007_/A sky130_fd_sc_hd__buf_2
Xinput76 core_dmem_request_put[66] vssd1 vssd1 vccd1 vccd1 _2043_/A sky130_fd_sc_hd__buf_2
XANTENNA__2308__A1 _1960_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3463_ _3473_/CLK _3463_/D vssd1 vssd1 vccd1 vccd1 _3463_/Q sky130_fd_sc_hd__dfxtp_1
X_2414_ _2414_/A vssd1 vssd1 vccd1 vccd1 _2414_/X sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_30_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3432_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3394_ _3394_/CLK _3394_/D vssd1 vssd1 vccd1 vccd1 _3394_/Q sky130_fd_sc_hd__dfxtp_1
X_2345_ _3417_/Q _2326_/X _2344_/Y vssd1 vssd1 vccd1 vccd1 _2345_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2276_ _2269_/X _2270_/X _2271_/X _1920_/C _2262_/X vssd1 vssd1 vccd1 vccd1 _2276_/Y
+ sky130_fd_sc_hd__o311ai_4
XFILLER_69_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_21_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3447_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1862__C _1862_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1770__A2 _1770_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input213_A ram_dmem_response_put[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_CLK clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3388_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2130_ _2130_/A vssd1 vssd1 vccd1 vccd1 _2131_/C sky130_fd_sc_hd__clkinv_2
XFILLER_93_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2061_ _2061_/A vssd1 vssd1 vccd1 vccd1 _2062_/C sky130_fd_sc_hd__clkinv_2
XFILLER_93_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_1_0_0_CLK_A clkbuf_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2963_ _3354_/Q _2779_/X _2959_/X _2143_/Y vssd1 vssd1 vccd1 vccd1 _3354_/D sky130_fd_sc_hd__o211a_1
X_1914_ _3290_/Q _1911_/X _1913_/Y vssd1 vssd1 vccd1 vccd1 _1914_/X sky130_fd_sc_hd__o21a_2
X_2894_ _3317_/Q _2893_/X _2011_/Y vssd1 vssd1 vccd1 vccd1 _2895_/A sky130_fd_sc_hd__o21ai_1
X_1845_ _2408_/A vssd1 vssd1 vccd1 vccd1 _1877_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1776_ _3259_/Q _1776_/B input8/X vssd1 vssd1 vccd1 vccd1 _1777_/A sky130_fd_sc_hd__or3_1
XFILLER_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2140__A _2169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3446_ _3452_/CLK _3446_/D vssd1 vssd1 vccd1 vccd1 _3446_/Q sky130_fd_sc_hd__dfxtp_1
X_3377_ _3461_/CLK _3377_/D vssd1 vssd1 vccd1 vccd1 _3377_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2328_ _2413_/A vssd1 vssd1 vccd1 vccd1 _2328_/X sky130_fd_sc_hd__clkbuf_4
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2701__A1 _1467_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2259_ _3387_/Q _2239_/X _2258_/Y vssd1 vssd1 vccd1 vccd1 _2259_/X sky130_fd_sc_hd__o21a_1
XFILLER_38_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2050__A _2050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input163_A fmc_dmem_response_put[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput211 ram_dmem_response_put[10] vssd1 vssd1 vccd1 vccd1 _2517_/A sky130_fd_sc_hd__buf_2
Xinput200 fmc_imem_response_put[2] vssd1 vssd1 vccd1 vccd1 _1654_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput233 ram_dmem_response_put[30] vssd1 vssd1 vccd1 vccd1 _2598_/A sky130_fd_sc_hd__buf_2
Xinput222 ram_dmem_response_put[20] vssd1 vssd1 vccd1 vccd1 _2560_/A sky130_fd_sc_hd__buf_2
Xinput244 ram_imem_response_put[11] vssd1 vssd1 vccd1 vccd1 _1694_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_75_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput266 ram_imem_response_put[31] vssd1 vssd1 vccd1 vccd1 _1774_/A sky130_fd_sc_hd__clkbuf_4
Xinput255 ram_imem_response_put[21] vssd1 vssd1 vccd1 vccd1 _1737_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input24_A core_dmem_request_put[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2456__B1 _2185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_1_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3244_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2225__A _2225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output382_A _1946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1630_ _3226_/Q _1630_/B vssd1 vssd1 vccd1 vccd1 _1631_/A sky130_fd_sc_hd__or2_1
X_1561_ _3198_/Q _1545_/X _1560_/Y vssd1 vssd1 vccd1 vccd1 _1561_/X sky130_fd_sc_hd__o21a_1
X_3300_ _3432_/CLK _3300_/D vssd1 vssd1 vccd1 vccd1 _3300_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1492_ _1512_/A _1520_/B _1492_/C vssd1 vssd1 vccd1 vccd1 _1492_/Y sky130_fd_sc_hd__nand3_1
XFILLER_86_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _3472_/CLK _3231_/D vssd1 vssd1 vccd1 vccd1 _3231_/Q sky130_fd_sc_hd__dfxtp_1
X_3162_ _3477_/CLK _3162_/D vssd1 vssd1 vccd1 vccd1 _3162_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2113_ _2127_/A _2134_/B _2113_/C vssd1 vssd1 vccd1 vccd1 _2113_/Y sky130_fd_sc_hd__nand3_1
XFILLER_94_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3093_ _3093_/A vssd1 vssd1 vccd1 vccd1 _3093_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2044_ _2072_/A _2044_/B _2044_/C vssd1 vssd1 vccd1 vccd1 _2044_/Y sky130_fd_sc_hd__nand3_1
XFILLER_47_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2998__A1 _1847_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2946_ _3344_/Q _2945_/X _2941_/X _2109_/Y vssd1 vssd1 vccd1 vccd1 _3344_/D sky130_fd_sc_hd__o211a_1
X_2877_ _3309_/Q _2873_/X _1981_/Y vssd1 vssd1 vccd1 vccd1 _2879_/A sky130_fd_sc_hd__o21ai_1
X_1828_ _1828_/A vssd1 vssd1 vccd1 vccd1 _1829_/C sky130_fd_sc_hd__inv_4
X_1759_ _1759_/A _1727_/X vssd1 vssd1 vccd1 vccd1 _1759_/X sky130_fd_sc_hd__or2b_1
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3429_ _3431_/CLK _3429_/D vssd1 vssd1 vccd1 vccd1 _3429_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_1_CLK_A clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2800_ _2959_/A vssd1 vssd1 vccd1 vccd1 _2878_/A sky130_fd_sc_hd__clkbuf_4
X_2731_ input4/X _2975_/B vssd1 vssd1 vccd1 vccd1 _2760_/A sky130_fd_sc_hd__nand2b_4
XFILLER_8_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1794__A _3116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2662_ _3181_/Q _2660_/X _2661_/X _1500_/Y vssd1 vssd1 vccd1 vccd1 _3181_/D sky130_fd_sc_hd__o211a_1
Xoutput526 _2194_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[4] sky130_fd_sc_hd__buf_2
Xoutput515 _2192_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[3] sky130_fd_sc_hd__buf_2
Xoutput504 _2190_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[2] sky130_fd_sc_hd__buf_2
X_1613_ _3216_/Q _1604_/X _1612_/Y vssd1 vssd1 vccd1 vccd1 _1613_/X sky130_fd_sc_hd__o21a_1
X_2593_ _2611_/B vssd1 vssd1 vccd1 vccd1 _2593_/Y sky130_fd_sc_hd__inv_2
Xoutput559 _2202_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[7] sky130_fd_sc_hd__buf_2
Xoutput548 _2200_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[6] sky130_fd_sc_hd__buf_2
Xoutput537 _2198_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[5] sky130_fd_sc_hd__buf_2
X_1544_ _2709_/A vssd1 vssd1 vccd1 vccd1 _1630_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__1707__A2 _1707_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3214_ _3384_/CLK _3214_/D vssd1 vssd1 vccd1 vccd1 _3214_/Q sky130_fd_sc_hd__dfxtp_1
X_1475_ _1475_/A vssd1 vssd1 vccd1 vccd1 _1476_/C sky130_fd_sc_hd__inv_2
XANTENNA__1960__C _1960_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3145_ _3140_/X _3145_/A2 _2548_/X _2549_/X _3141_/X vssd1 vssd1 vccd1 vccd1 _3479_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_27_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3076_ _3429_/Q _3065_/X _2378_/Y _3075_/X vssd1 vssd1 vccd1 vccd1 _3429_/D sky130_fd_sc_hd__o211a_1
XFILLER_82_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1969__A _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2027_ _3321_/Q _2020_/X _2026_/Y vssd1 vssd1 vccd1 vccd1 _2027_/X sky130_fd_sc_hd__o21a_2
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2929_ _2929_/A _2933_/B vssd1 vssd1 vccd1 vccd1 _3335_/D sky130_fd_sc_hd__nand2_1
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input126_A core_imem_request_put[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input91_A core_dmem_request_put[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output512_A _2290_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput8 EN_fmc_imem_response_put vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_4
XANTENNA__2114__A2 _2111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2714_ _3214_/Q _2709_/X _1608_/Y _2710_/X vssd1 vssd1 vccd1 vccd1 _3214_/D sky130_fd_sc_hd__o211a_1
XFILLER_10_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput301 _2575_/X vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[23] sky130_fd_sc_hd__buf_2
X_2645_ _3172_/Q _2644_/X _1467_/Y vssd1 vssd1 vccd1 vccd1 _2646_/A sky130_fd_sc_hd__o21ai_1
Xoutput323 _1708_/Y vssd1 vssd1 vccd1 vccd1 core_imem_response_get[14] sky130_fd_sc_hd__buf_2
Xoutput312 _2493_/Y vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[4] sky130_fd_sc_hd__buf_2
Xoutput334 _1750_/Y vssd1 vssd1 vccd1 vccd1 core_imem_response_get[24] sky130_fd_sc_hd__buf_2
Xoutput378 _1932_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[35] sky130_fd_sc_hd__buf_2
Xoutput367 _1895_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[25] sky130_fd_sc_hd__buf_2
Xoutput345 _1667_/X vssd1 vssd1 vccd1 vccd1 core_imem_response_get[5] sky130_fd_sc_hd__buf_2
X_2576_ _2542_/X _3486_/Q _2543_/X vssd1 vssd1 vccd1 vccd1 _2576_/X sky130_fd_sc_hd__o21ba_1
Xoutput356 _1855_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[15] sky130_fd_sc_hd__buf_2
Xoutput389 _1968_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[45] sky130_fd_sc_hd__buf_2
X_1527_ _1527_/A _1527_/B _1527_/C vssd1 vssd1 vccd1 vccd1 _1527_/Y sky130_fd_sc_hd__nand3_1
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1458_ _1597_/A vssd1 vssd1 vccd1 vccd1 _1488_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_55_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3128_ _3143_/A vssd1 vssd1 vccd1 vccd1 _3128_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3059_ _3417_/Q _3051_/X _2344_/Y _3047_/X vssd1 vssd1 vccd1 vccd1 _3417_/D sky130_fd_sc_hd__o211a_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2026__C _2026_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2323__A _2351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2592__A2 _2592_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3154__A _3154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input243_A ram_imem_response_put[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1751__B1_N _1743_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output462_A _1501_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2430_ _2412_/X _2413_/X _2414_/X _2117_/C _2405_/X vssd1 vssd1 vccd1 vccd1 _2430_/Y
+ sky130_fd_sc_hd__o311ai_4
X_2361_ _2341_/X _2351_/X _3422_/Q vssd1 vssd1 vccd1 vccd1 _2361_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__1543__B1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2292_ _2269_/X _2270_/X _2271_/X _1942_/C _2291_/X vssd1 vssd1 vccd1 vccd1 _2292_/Y
+ sky130_fd_sc_hd__o311ai_2
XANTENNA__2740__C1 _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_41_CLK_A clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2408__A _2408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2628_ _3163_/Q _2619_/X _2621_/X _1432_/Y vssd1 vssd1 vccd1 vccd1 _3163_/D sky130_fd_sc_hd__o211a_1
X_2559_ _2542_/X _3482_/Q _2543_/X vssd1 vssd1 vccd1 vccd1 _2559_/X sky130_fd_sc_hd__o21ba_1
XFILLER_87_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2798__C1 _1829_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input193_A fmc_imem_response_put[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2988__A _3095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input54_A core_dmem_request_put[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2722__C1 _2686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3114__B_N _2682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1930_ _1930_/A vssd1 vssd1 vccd1 vccd1 _1931_/C sky130_fd_sc_hd__inv_2
XFILLER_14_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1861_ _1861_/A vssd1 vssd1 vccd1 vccd1 _1862_/C sky130_fd_sc_hd__clkinv_4
Xinput11 EN_ram_imem_request_get vssd1 vssd1 vccd1 vccd1 _2723_/A sky130_fd_sc_hd__clkbuf_2
Xinput22 core_dmem_request_put[17] vssd1 vssd1 vccd1 vccd1 _1861_/A sky130_fd_sc_hd__clkbuf_1
Xinput33 core_dmem_request_put[27] vssd1 vssd1 vccd1 vccd1 _1900_/A sky130_fd_sc_hd__clkbuf_1
Xinput55 core_dmem_request_put[47] vssd1 vssd1 vccd1 vccd1 _1973_/A sky130_fd_sc_hd__clkbuf_1
Xinput44 core_dmem_request_put[37] vssd1 vssd1 vccd1 vccd1 _1937_/A sky130_fd_sc_hd__clkbuf_1
X_1792_ _2206_/A vssd1 vssd1 vccd1 vccd1 _1821_/B sky130_fd_sc_hd__clkbuf_2
Xinput66 core_dmem_request_put[57] vssd1 vssd1 vccd1 vccd1 _2010_/A sky130_fd_sc_hd__clkbuf_1
Xinput77 core_dmem_request_put[67] vssd1 vssd1 vccd1 vccd1 _2046_/A sky130_fd_sc_hd__clkbuf_1
Xinput88 core_dmem_request_put[77] vssd1 vssd1 vccd1 vccd1 _2083_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__2898__A _2936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput99 core_dmem_request_put[87] vssd1 vssd1 vccd1 vccd1 _2119_/A sky130_fd_sc_hd__clkbuf_2
X_3462_ _3473_/CLK _3462_/D vssd1 vssd1 vccd1 vccd1 _3462_/Q sky130_fd_sc_hd__dfxtp_1
X_3393_ _3397_/CLK _3393_/D vssd1 vssd1 vccd1 vccd1 _3393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2413_ _2413_/A vssd1 vssd1 vccd1 vccd1 _2413_/X sky130_fd_sc_hd__buf_4
XFILLER_69_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2344_ _2327_/X _2328_/X _2329_/X _2008_/C _2320_/X vssd1 vssd1 vccd1 vccd1 _2344_/Y
+ sky130_fd_sc_hd__o311ai_4
X_2275_ _1917_/C _2253_/X _2274_/Y vssd1 vssd1 vccd1 vccd1 _2275_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_52_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2492__A1 _2462_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1977__A _1977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2483__A1 _2462_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input206_A fmc_imem_response_put[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2786__A2 _2779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2171__B1 _2163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2060_ _2097_/A vssd1 vssd1 vccd1 vccd1 _2091_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1797__A _1951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2962_ _2962_/A _2965_/B vssd1 vssd1 vccd1 vccd1 _3353_/D sky130_fd_sc_hd__nand2_1
XFILLER_15_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1913_ _1927_/A _1935_/B _1913_/C vssd1 vssd1 vccd1 vccd1 _1913_/Y sky130_fd_sc_hd__nand3_1
XFILLER_30_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2893_ _2893_/A vssd1 vssd1 vccd1 vccd1 _2893_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1844_ _3272_/Q _1834_/X _1843_/Y vssd1 vssd1 vccd1 vccd1 _1844_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1775_ _1772_/X _2772_/A2 _1773_/X _1774_/X vssd1 vssd1 vccd1 vccd1 _1775_/X sky130_fd_sc_hd__a22o_4
XANTENNA__1963__C _1963_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3445_ _3447_/CLK _3445_/D vssd1 vssd1 vccd1 vccd1 _3445_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2140__B _2967_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3376_ _3384_/CLK _3376_/D vssd1 vssd1 vccd1 vccd1 _3376_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2327_ _2412_/A vssd1 vssd1 vccd1 vccd1 _2327_/X sky130_fd_sc_hd__clkbuf_4
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2258_ _2240_/X _2241_/X _2242_/X _1898_/C _2232_/X vssd1 vssd1 vccd1 vccd1 _2258_/Y
+ sky130_fd_sc_hd__o311ai_2
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2189_ _2176_/X _2178_/X _2180_/X _1804_/C _2152_/A vssd1 vssd1 vccd1 vccd1 _2189_/Y
+ sky130_fd_sc_hd__o311ai_2
XANTENNA__2465__A1 _2464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2217__A1 _1840_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2768__A2 _2768_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1873__C _1873_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput201 fmc_imem_response_put[30] vssd1 vssd1 vccd1 vccd1 _1770_/A2 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input156_A fmc_dmem_response_put[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput234 ram_dmem_response_put[31] vssd1 vssd1 vccd1 vccd1 _2603_/A sky130_fd_sc_hd__clkbuf_4
Xinput223 ram_dmem_response_put[21] vssd1 vssd1 vccd1 vccd1 _2566_/A sky130_fd_sc_hd__clkbuf_4
Xinput212 ram_dmem_response_put[11] vssd1 vssd1 vccd1 vccd1 _2523_/A sky130_fd_sc_hd__clkbuf_4
Xinput245 ram_imem_response_put[12] vssd1 vssd1 vccd1 vccd1 _1697_/A sky130_fd_sc_hd__buf_2
XFILLER_88_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput256 ram_imem_response_put[22] vssd1 vssd1 vccd1 vccd1 _1740_/A sky130_fd_sc_hd__clkbuf_2
Xinput267 ram_imem_response_put[3] vssd1 vssd1 vccd1 vccd1 _1658_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_75_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input17_A core_dmem_request_put[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2456__A1 _2169_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2208__A1 _1832_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2506__A _2506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2759__A2 _2759_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output375_A _1921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1560_ _1546_/X _1547_/X _1548_/X _1438_/C _1527_/A vssd1 vssd1 vccd1 vccd1 _1560_/Y
+ sky130_fd_sc_hd__o311ai_4
X_1491_ _1491_/A vssd1 vssd1 vccd1 vccd1 _1492_/C sky130_fd_sc_hd__inv_2
XFILLER_3_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _3259_/CLK _3230_/D vssd1 vssd1 vccd1 vccd1 _3230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3161_ _3489_/CLK _3161_/D vssd1 vssd1 vccd1 vccd1 _3161_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2112_ _2112_/A vssd1 vssd1 vccd1 vccd1 _2113_/C sky130_fd_sc_hd__clkinv_2
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3092_ _2091_/C _3091_/X _3081_/X _2409_/Y vssd1 vssd1 vccd1 vccd1 _3440_/D sky130_fd_sc_hd__o211ai_1
XFILLER_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2043_ _2043_/A vssd1 vssd1 vccd1 vccd1 _2044_/C sky130_fd_sc_hd__inv_2
XFILLER_22_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2945_ _2945_/A vssd1 vssd1 vccd1 vccd1 _2945_/X sky130_fd_sc_hd__clkbuf_2
X_2876_ _3308_/Q _2868_/X _2864_/X _1978_/Y vssd1 vssd1 vccd1 vccd1 _3308_/D sky130_fd_sc_hd__o211a_1
X_1827_ _2967_/B vssd1 vssd1 vccd1 vccd1 _1859_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_30_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2151__A _2151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1758_ _1735_/X _3254_/Q _1743_/X vssd1 vssd1 vccd1 vccd1 _1758_/X sky130_fd_sc_hd__o21ba_1
X_1689_ _1669_/X _1689_/A2 _1687_/X _1688_/X vssd1 vssd1 vccd1 vccd1 _2748_/B sky130_fd_sc_hd__a22oi_4
X_3428_ _3452_/CLK _3428_/D vssd1 vssd1 vccd1 vccd1 _3428_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_input9_A EN_ram_dmem_request_get vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3359_ _3460_/CLK _3359_/D vssd1 vssd1 vccd1 vccd1 _3359_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input273_A ram_imem_response_put[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2236__A _2351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2730_ _3226_/Q _2681_/X _2684_/X vssd1 vssd1 vccd1 vccd1 _3226_/D sky130_fd_sc_hd__o21a_1
X_2661_ _2677_/B vssd1 vssd1 vccd1 vccd1 _2661_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3067__A _3067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1612_ _1605_/X _1606_/X _1607_/X _1506_/C _1594_/X vssd1 vssd1 vccd1 vccd1 _1612_/Y
+ sky130_fd_sc_hd__o311ai_4
XFILLER_8_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput516 _2302_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[40] sky130_fd_sc_hd__buf_2
Xoutput505 _2273_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[30] sky130_fd_sc_hd__buf_2
Xoutput527 _2331_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[50] sky130_fd_sc_hd__buf_2
X_2592_ _2520_/A _2592_/A2 _2590_/X _2591_/X vssd1 vssd1 vccd1 vccd1 _2611_/B sky130_fd_sc_hd__a22oi_4
Xoutput538 _2360_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[60] sky130_fd_sc_hd__buf_2
Xoutput549 _2388_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[70] sky130_fd_sc_hd__buf_2
X_1543_ _1529_/A _1531_/A _1533_/A input3/X vssd1 vssd1 vccd1 vccd1 _2709_/A sky130_fd_sc_hd__o31a_2
X_1474_ _3174_/Q _1462_/X _1473_/Y vssd1 vssd1 vccd1 vccd1 _1474_/X sky130_fd_sc_hd__o21a_2
X_3213_ _3222_/CLK _3213_/D vssd1 vssd1 vccd1 vccd1 _3213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3144_ _3152_/A _3144_/B vssd1 vssd1 vccd1 vccd1 _3478_/D sky130_fd_sc_hd__nor2_1
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3075_ _3075_/A vssd1 vssd1 vccd1 vccd1 _3075_/X sky130_fd_sc_hd__clkbuf_2
X_2026_ _2054_/A _2026_/B _2026_/C vssd1 vssd1 vccd1 vccd1 _2026_/Y sky130_fd_sc_hd__nand3_1
XFILLER_23_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2146__A _2146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1985__A _1985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2928_ _3335_/Q _2912_/X _2077_/Y vssd1 vssd1 vccd1 vccd1 _2929_/A sky130_fd_sc_hd__o21ai_1
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2859_ _2878_/A vssd1 vssd1 vccd1 vccd1 _2875_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input119_A core_imem_request_put[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3084__A1 _2069_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input84_A core_dmem_request_put[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput9 EN_ram_dmem_request_get vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_2
XFILLER_64_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_0_CLK_A clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2713_ _1496_/C _2707_/X _2712_/X _1602_/Y vssd1 vssd1 vccd1 vccd1 _3213_/D sky130_fd_sc_hd__o211ai_1
X_2644_ _2660_/A vssd1 vssd1 vccd1 vccd1 _2644_/X sky130_fd_sc_hd__clkbuf_2
X_2575_ _2563_/X _3151_/A2 _2573_/X _2574_/X vssd1 vssd1 vccd1 vccd1 _2575_/X sky130_fd_sc_hd__a22o_1
Xoutput335 _1753_/X vssd1 vssd1 vccd1 vccd1 core_imem_response_get[25] sky130_fd_sc_hd__buf_2
Xoutput324 _1711_/X vssd1 vssd1 vccd1 vccd1 core_imem_response_get[15] sky130_fd_sc_hd__buf_2
Xoutput313 _2496_/X vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[5] sky130_fd_sc_hd__buf_2
Xoutput302 _2579_/Y vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[24] sky130_fd_sc_hd__buf_2
XANTENNA__1971__C _1971_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput368 _1899_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[26] sky130_fd_sc_hd__buf_2
Xoutput346 _1675_/Y vssd1 vssd1 vccd1 vccd1 core_imem_response_get[6] sky130_fd_sc_hd__buf_2
X_1526_ _1526_/A vssd1 vssd1 vccd1 vccd1 _1527_/C sky130_fd_sc_hd__inv_2
Xoutput357 _1860_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[16] sky130_fd_sc_hd__buf_2
Xoutput379 _1936_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[36] sky130_fd_sc_hd__buf_2
X_1457_ _3169_/Q _1441_/X _1456_/Y vssd1 vssd1 vccd1 vccd1 _1457_/X sky130_fd_sc_hd__o21a_2
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3127_ _3140_/A vssd1 vssd1 vccd1 vccd1 _3127_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3058_ _2004_/C _3049_/X _3053_/X _2342_/Y vssd1 vssd1 vccd1 vccd1 _3416_/D sky130_fd_sc_hd__o211ai_1
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2009_ _3316_/Q _2002_/X _2008_/Y vssd1 vssd1 vccd1 vccd1 _2009_/X sky130_fd_sc_hd__o21a_1
XFILLER_63_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2041__A2 _2038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1762__B_N _1644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input236_A ram_dmem_response_put[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2514__A _2514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output455_A _1477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2360_ _3421_/Q _2355_/X _2359_/Y vssd1 vssd1 vccd1 vccd1 _2360_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1543__A1 _1529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2291_ _2291_/A vssd1 vssd1 vccd1 vccd1 _2291_/X sky130_fd_sc_hd__buf_2
XFILLER_64_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2023__A2 _2020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2627_ _2627_/A _2636_/B vssd1 vssd1 vccd1 vccd1 _3162_/D sky130_fd_sc_hd__nand2_1
X_2558_ _2520_/X _3147_/A2 _2555_/X _2557_/X vssd1 vssd1 vccd1 vccd1 _2558_/X sky130_fd_sc_hd__a22o_1
X_1509_ _1516_/A _1523_/B _1509_/C vssd1 vssd1 vccd1 vccd1 _1509_/Y sky130_fd_sc_hd__nand3_1
X_2489_ _2464_/X _3466_/Q _2470_/A vssd1 vssd1 vccd1 vccd1 _2489_/X sky130_fd_sc_hd__o21ba_1
XFILLER_87_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input186_A fmc_imem_response_put[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input47_A core_dmem_request_put[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1413__A _1529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2509__A _2509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1860_ _3276_/Q _1852_/X _1859_/Y vssd1 vssd1 vccd1 vccd1 _1860_/X sky130_fd_sc_hd__o21a_1
XFILLER_42_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 EN_ram_imem_response_put vssd1 vssd1 vccd1 vccd1 _1776_/B sky130_fd_sc_hd__buf_4
XANTENNA_output572_A _2443_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1791_ _2104_/A vssd1 vssd1 vccd1 vccd1 _2206_/A sky130_fd_sc_hd__buf_4
XANTENNA__2005__A2 _2002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput34 core_dmem_request_put[28] vssd1 vssd1 vccd1 vccd1 _1905_/A sky130_fd_sc_hd__clkbuf_1
Xinput23 core_dmem_request_put[18] vssd1 vssd1 vccd1 vccd1 _1865_/A sky130_fd_sc_hd__clkbuf_1
Xinput45 core_dmem_request_put[38] vssd1 vssd1 vccd1 vccd1 _1941_/A sky130_fd_sc_hd__clkbuf_1
Xinput89 core_dmem_request_put[78] vssd1 vssd1 vccd1 vccd1 _2087_/A sky130_fd_sc_hd__buf_2
Xinput56 core_dmem_request_put[48] vssd1 vssd1 vccd1 vccd1 _1977_/A sky130_fd_sc_hd__buf_2
Xinput67 core_dmem_request_put[58] vssd1 vssd1 vccd1 vccd1 _2014_/A sky130_fd_sc_hd__buf_2
Xinput78 core_dmem_request_put[68] vssd1 vssd1 vccd1 vccd1 _2050_/A sky130_fd_sc_hd__buf_2
X_3461_ _3461_/CLK _3461_/D vssd1 vssd1 vccd1 vccd1 _3461_/Q sky130_fd_sc_hd__dfxtp_4
X_2412_ _2412_/A vssd1 vssd1 vccd1 vccd1 _2412_/X sky130_fd_sc_hd__buf_4
X_3392_ _3394_/CLK _3392_/D vssd1 vssd1 vccd1 vccd1 _3392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2343_ _2004_/C _2340_/X _2342_/Y vssd1 vssd1 vccd1 vccd1 _2343_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_84_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2274_ _2255_/X _2265_/X _3392_/Q vssd1 vssd1 vccd1 vccd1 _2274_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_37_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2492__A2 _2492_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2154__A _2175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1989_ _1989_/A vssd1 vssd1 vccd1 vccd1 _1990_/C sky130_fd_sc_hd__inv_2
XFILLER_20_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2483__A2 _2483_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input101_A core_dmem_request_put[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1765__B1_N _1743_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2064__A _2064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_40_CLK_A clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1746__A1 _1734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2171__A1 _2175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output418_A _2063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output320_A _1695_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2961_ _3353_/Q _2950_/X _2140_/Y vssd1 vssd1 vccd1 vccd1 _2962_/A sky130_fd_sc_hd__o21ai_1
X_1912_ _1912_/A vssd1 vssd1 vccd1 vccd1 _1913_/C sky130_fd_sc_hd__clkinv_4
X_2892_ _3316_/Q _2888_/X _2884_/X _2008_/Y vssd1 vssd1 vccd1 vccd1 _3316_/D sky130_fd_sc_hd__o211a_1
XFILLER_30_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1843_ _1850_/A _1859_/B _1843_/C vssd1 vssd1 vccd1 vccd1 _1843_/Y sky130_fd_sc_hd__nand3_2
X_1774_ _1774_/A _1635_/X vssd1 vssd1 vccd1 vccd1 _1774_/X sky130_fd_sc_hd__or2b_1
X_3444_ _3448_/CLK _3444_/D vssd1 vssd1 vccd1 vccd1 _3444_/Q sky130_fd_sc_hd__dfxtp_1
X_3375_ _3461_/CLK _3375_/D vssd1 vssd1 vccd1 vccd1 _3375_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2326_ _2326_/A vssd1 vssd1 vccd1 vccd1 _2326_/X sky130_fd_sc_hd__clkbuf_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2149__A _2319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2257_ _1894_/C _2253_/X _2256_/Y vssd1 vssd1 vccd1 vccd1 _2257_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_84_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2188_ _1801_/C _2185_/X _2187_/Y vssd1 vssd1 vccd1 vccd1 _2188_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_65_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2479__B_N _2478_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput202 fmc_imem_response_put[31] vssd1 vssd1 vccd1 vccd1 _2772_/A2 sky130_fd_sc_hd__buf_4
Xinput224 ram_dmem_response_put[22] vssd1 vssd1 vccd1 vccd1 _2569_/A sky130_fd_sc_hd__buf_2
Xinput213 ram_dmem_response_put[12] vssd1 vssd1 vccd1 vccd1 _2526_/A sky130_fd_sc_hd__buf_2
Xinput235 ram_dmem_response_put[3] vssd1 vssd1 vccd1 vccd1 _2487_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input149_A fmc_dmem_response_put[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput257 ram_imem_response_put[23] vssd1 vssd1 vccd1 vccd1 _1745_/A sky130_fd_sc_hd__clkbuf_2
Xinput246 ram_imem_response_put[13] vssd1 vssd1 vccd1 vccd1 _1702_/A sky130_fd_sc_hd__clkbuf_2
Xinput268 ram_imem_response_put[4] vssd1 vssd1 vccd1 vccd1 _1662_/A sky130_fd_sc_hd__buf_2
XFILLER_75_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2613__C1 _3154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output368_A _1899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1490_ _2675_/B vssd1 vssd1 vccd1 vccd1 _1520_/B sky130_fd_sc_hd__clkbuf_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _3466_/CLK _3160_/D vssd1 vssd1 vccd1 vccd1 _3160_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2111_ _2145_/A vssd1 vssd1 vccd1 vccd1 _2111_/X sky130_fd_sc_hd__buf_2
X_3091_ _3091_/A vssd1 vssd1 vccd1 vccd1 _3091_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2042_ _2967_/A vssd1 vssd1 vccd1 vccd1 _2072_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2447__A2 _2426_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2944_ _2944_/A _2952_/B vssd1 vssd1 vccd1 vccd1 _3343_/D sky130_fd_sc_hd__nand2_1
XFILLER_30_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2875_ _2875_/A _2875_/B vssd1 vssd1 vccd1 vccd1 _3307_/D sky130_fd_sc_hd__nand2_1
X_1826_ _2104_/A vssd1 vssd1 vccd1 vccd1 _2967_/B sky130_fd_sc_hd__buf_4
XANTENNA__1974__C _1974_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1757_ _2767_/B vssd1 vssd1 vccd1 vccd1 _1757_/Y sky130_fd_sc_hd__inv_2
X_1688_ _1688_/A _1661_/X vssd1 vssd1 vccd1 vccd1 _1688_/X sky130_fd_sc_hd__or2b_1
X_3427_ _3431_/CLK _3427_/D vssd1 vssd1 vccd1 vccd1 _3427_/Q sky130_fd_sc_hd__dfxtp_1
X_3358_ _3394_/CLK _3358_/D vssd1 vssd1 vccd1 vccd1 _3358_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2309_ _2298_/X _2299_/X _2300_/X _1963_/C _2291_/X vssd1 vssd1 vccd1 vccd1 _2309_/Y
+ sky130_fd_sc_hd__o311ai_4
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3289_ _3486_/CLK _3289_/D vssd1 vssd1 vccd1 vccd1 _3289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2438__A2 _2426_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2607__A _2975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input266_A ram_imem_response_put[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2429__A2 _2426_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2517__A _2517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1421__A _2675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1794__C _1794_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2660_ _2660_/A vssd1 vssd1 vccd1 vccd1 _2660_/X sky130_fd_sc_hd__clkbuf_2
X_1611_ _1503_/C _1590_/X _1610_/Y vssd1 vssd1 vccd1 vccd1 _1611_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_60_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput506 _2275_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[31] sky130_fd_sc_hd__buf_2
Xoutput517 _2304_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[41] sky130_fd_sc_hd__buf_2
X_2591_ _2591_/A _2473_/A vssd1 vssd1 vccd1 vccd1 _2591_/X sky130_fd_sc_hd__or2b_1
Xoutput528 _2333_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[51] sky130_fd_sc_hd__buf_2
Xoutput539 _2362_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[61] sky130_fd_sc_hd__buf_2
X_1542_ _1541_/X _1447_/B _3193_/Q vssd1 vssd1 vccd1 vccd1 _1542_/X sky130_fd_sc_hd__a21o_4
XFILLER_5_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1473_ _1480_/A _1488_/B _1473_/C vssd1 vssd1 vccd1 vccd1 _1473_/Y sky130_fd_sc_hd__nand3_1
XFILLER_86_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3212_ _3222_/CLK _3212_/D vssd1 vssd1 vccd1 vccd1 _3212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3143_ _3143_/A vssd1 vssd1 vccd1 vccd1 _3152_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3074_ _2047_/C _3063_/X _3067_/X _2375_/Y vssd1 vssd1 vccd1 vccd1 _3428_/D sky130_fd_sc_hd__o211ai_1
XFILLER_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2025_ _2025_/A vssd1 vssd1 vccd1 vccd1 _2026_/C sky130_fd_sc_hd__inv_2
XFILLER_35_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2927_ _3334_/Q _2926_/X _2922_/X _2072_/Y vssd1 vssd1 vccd1 vccd1 _3334_/D sky130_fd_sc_hd__o211a_1
XFILLER_10_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2858_ _3299_/Q _2854_/X _1945_/Y vssd1 vssd1 vccd1 vccd1 _2860_/A sky130_fd_sc_hd__o21ai_1
X_1809_ _3263_/Q _1784_/X _1808_/Y vssd1 vssd1 vccd1 vccd1 _1809_/X sky130_fd_sc_hd__o21a_1
X_2789_ _2868_/A vssd1 vssd1 vccd1 vccd1 _2789_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2292__B1 _1942_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2347__A1 _2011_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input77_A core_dmem_request_put[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2800__A _2959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1416__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output400_A _2005_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2807__C1 _1843_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2712_ _2712_/A vssd1 vssd1 vccd1 vccd1 _2712_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2643_ _3171_/Q _2641_/X _2642_/X _1464_/Y vssd1 vssd1 vccd1 vccd1 _3171_/D sky130_fd_sc_hd__o211a_1
X_2574_ _2574_/A _2556_/X vssd1 vssd1 vccd1 vccd1 _2574_/X sky130_fd_sc_hd__or2b_1
Xoutput325 _1718_/Y vssd1 vssd1 vccd1 vccd1 core_imem_response_get[16] sky130_fd_sc_hd__buf_2
Xoutput314 _2504_/Y vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[6] sky130_fd_sc_hd__buf_2
Xoutput303 _2582_/X vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[25] sky130_fd_sc_hd__buf_2
Xoutput369 _1902_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[27] sky130_fd_sc_hd__buf_2
X_1525_ _1597_/A vssd1 vssd1 vccd1 vccd1 _1527_/B sky130_fd_sc_hd__buf_2
Xoutput347 _1678_/X vssd1 vssd1 vccd1 vccd1 core_imem_response_get[7] sky130_fd_sc_hd__buf_2
Xoutput336 _1757_/Y vssd1 vssd1 vccd1 vccd1 core_imem_response_get[26] sky130_fd_sc_hd__buf_2
Xoutput358 _1863_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[17] sky130_fd_sc_hd__buf_2
XFILLER_59_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1456_ _1476_/A _1484_/B _1456_/C vssd1 vssd1 vccd1 vccd1 _1456_/Y sky130_fd_sc_hd__nand3_1
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3126_ _3126_/A _3126_/B vssd1 vssd1 vccd1 vccd1 _3466_/D sky130_fd_sc_hd__nor2_1
XANTENNA__2157__A _2177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3057_ _3415_/Q _3051_/X _2338_/Y _3047_/X vssd1 vssd1 vccd1 vccd1 _3415_/D sky130_fd_sc_hd__o211a_1
XFILLER_82_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2008_ _2036_/A _2008_/B _2008_/C vssd1 vssd1 vccd1 vccd1 _2008_/Y sky130_fd_sc_hd__nand3_1
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2620__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_51_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3258_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input131_A core_imem_request_put[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input229_A ram_dmem_response_put[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_42_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3247_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_output448_A _2168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1543__A2 _1531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2290_ _1938_/C _2283_/X _2289_/Y vssd1 vssd1 vccd1 vccd1 _2290_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2143__C _2143_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2626_ _2658_/A vssd1 vssd1 vccd1 vccd1 _2636_/B sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_33_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3436_/CLK sky130_fd_sc_hd__clkbuf_16
X_2557_ _2557_/A _2556_/X vssd1 vssd1 vccd1 vccd1 _2557_/X sky130_fd_sc_hd__or2b_1
X_2488_ _2471_/X _3125_/A2 _2486_/X _2487_/X vssd1 vssd1 vccd1 vccd1 _2488_/X sky130_fd_sc_hd__a22o_1
X_1508_ _1508_/A vssd1 vssd1 vccd1 vccd1 _1509_/C sky130_fd_sc_hd__inv_2
XFILLER_87_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1439_ _3165_/Q _1415_/X _1438_/Y vssd1 vssd1 vccd1 vccd1 _1439_/X sky130_fd_sc_hd__o21a_2
XFILLER_68_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3109_ _3453_/Q _2174_/A _2444_/Y _3103_/X vssd1 vssd1 vccd1 vccd1 _3453_/D sky130_fd_sc_hd__o211a_1
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2247__B1 _1880_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_CLK clkbuf_2_3_0_CLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_CLK/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_24_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3454_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input179_A fmc_imem_response_put[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1413__B _1531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output398_A _1998_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput13 RST_N vssd1 vssd1 vccd1 vccd1 _2975_/B sky130_fd_sc_hd__buf_6
X_1790_ _2235_/A vssd1 vssd1 vccd1 vccd1 _2104_/A sky130_fd_sc_hd__clkbuf_2
Xinput35 core_dmem_request_put[29] vssd1 vssd1 vccd1 vccd1 _1908_/A sky130_fd_sc_hd__clkbuf_1
Xinput46 core_dmem_request_put[39] vssd1 vssd1 vccd1 vccd1 _1944_/A sky130_fd_sc_hd__clkbuf_1
Xinput24 core_dmem_request_put[19] vssd1 vssd1 vccd1 vccd1 _1868_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_output565_A _2429_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput57 core_dmem_request_put[49] vssd1 vssd1 vccd1 vccd1 _1980_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput68 core_dmem_request_put[59] vssd1 vssd1 vccd1 vccd1 _2017_/A sky130_fd_sc_hd__clkbuf_2
Xinput79 core_dmem_request_put[69] vssd1 vssd1 vccd1 vccd1 _2053_/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_15_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3460_/CLK sky130_fd_sc_hd__clkbuf_16
X_3460_ _3460_/CLK _3460_/D vssd1 vssd1 vccd1 vccd1 _3460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2411_ _2459_/B vssd1 vssd1 vccd1 vccd1 _2411_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3391_ _3397_/CLK _3391_/D vssd1 vssd1 vccd1 vccd1 _3391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2713__A1 _1496_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2342_ _2341_/X _2323_/X _3416_/Q vssd1 vssd1 vccd1 vccd1 _2342_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2273_ _3391_/Q _2268_/X _2272_/Y vssd1 vssd1 vccd1 vccd1 _2273_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1604__A _1630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3091__A _3091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1988_ _2097_/A vssd1 vssd1 vccd1 vccd1 _2018_/A sky130_fd_sc_hd__clkbuf_2
X_2609_ _3143_/A vssd1 vssd1 vccd1 vccd1 _3130_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1746__A2 _2764_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2080__A _2080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2171__A2 _2177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2682__A_N _2723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3120__A1 _3116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_4_CLK clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3197_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2960_ _3352_/Q _2945_/X _2959_/X _2137_/Y vssd1 vssd1 vccd1 vccd1 _3352_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2255__A _2370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1911_ _1965_/A vssd1 vssd1 vccd1 vccd1 _1911_/X sky130_fd_sc_hd__clkbuf_2
X_2891_ _2891_/A _2895_/B vssd1 vssd1 vccd1 vccd1 _3315_/D sky130_fd_sc_hd__nand2_1
XFILLER_8_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1842_ _1842_/A vssd1 vssd1 vccd1 vccd1 _1843_/C sky130_fd_sc_hd__inv_4
XFILLER_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1773_ _1649_/X _3258_/Q _1743_/X vssd1 vssd1 vccd1 vccd1 _1773_/X sky130_fd_sc_hd__o21ba_1
X_3443_ _3447_/CLK _3443_/D vssd1 vssd1 vccd1 vccd1 _3443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _3384_/CLK _3374_/D vssd1 vssd1 vccd1 vccd1 _3374_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2325_ _1981_/C _2311_/X _2324_/Y vssd1 vssd1 vccd1 vccd1 _2325_/Y sky130_fd_sc_hd__o21ai_4
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2256_ _2255_/X _2236_/X _3386_/Q vssd1 vssd1 vccd1 vccd1 _2256_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_38_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2187_ _2165_/X _2186_/X _3362_/Q vssd1 vssd1 vccd1 vccd1 _2187_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_53_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2165__A _2225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1500__C _1500_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2153__A2 _2145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2689__B1 _2686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput225 ram_dmem_response_put[23] vssd1 vssd1 vccd1 vccd1 _2574_/A sky130_fd_sc_hd__clkbuf_4
Xinput214 ram_dmem_response_put[13] vssd1 vssd1 vccd1 vccd1 _2531_/A sky130_fd_sc_hd__clkbuf_4
Xinput236 ram_dmem_response_put[4] vssd1 vssd1 vccd1 vccd1 _2491_/A sky130_fd_sc_hd__buf_2
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput203 fmc_imem_response_put[3] vssd1 vssd1 vccd1 vccd1 _2738_/A2 sky130_fd_sc_hd__buf_4
Xinput269 ram_imem_response_put[5] vssd1 vssd1 vccd1 vccd1 _1666_/A sky130_fd_sc_hd__clkbuf_2
Xinput258 ram_imem_response_put[24] vssd1 vssd1 vccd1 vccd1 _1748_/A sky130_fd_sc_hd__clkbuf_2
Xinput247 ram_imem_response_put[14] vssd1 vssd1 vccd1 vccd1 _1706_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input211_A ram_dmem_response_put[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1419__A _1529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output528_A _2333_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3090_ _3439_/Q _3079_/X _2406_/Y _3089_/X vssd1 vssd1 vccd1 vccd1 _3439_/D sky130_fd_sc_hd__o211a_1
X_2110_ _3344_/Q _2093_/X _2109_/Y vssd1 vssd1 vccd1 vccd1 _2110_/X sky130_fd_sc_hd__o21a_1
XFILLER_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2041_ _3325_/Q _2038_/X _2040_/Y vssd1 vssd1 vccd1 vccd1 _2041_/X sky130_fd_sc_hd__o21a_2
XFILLER_94_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2943_ _3343_/Q _2931_/X _2106_/Y vssd1 vssd1 vccd1 vccd1 _2944_/A sky130_fd_sc_hd__o21ai_1
X_2874_ _3307_/Q _2873_/X _1974_/Y vssd1 vssd1 vccd1 vccd1 _2875_/A sky130_fd_sc_hd__o21ai_1
X_1825_ _3267_/Q _1813_/X _1824_/Y vssd1 vssd1 vccd1 vccd1 _1825_/X sky130_fd_sc_hd__o21a_1
X_1756_ _1691_/A _1756_/A2 _1754_/X _1755_/X vssd1 vssd1 vccd1 vccd1 _2767_/B sky130_fd_sc_hd__a22oi_4
XFILLER_89_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1687_ _1670_/X _3237_/Q _1671_/X vssd1 vssd1 vccd1 vccd1 _1687_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__1990__C _1990_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3426_ _3448_/CLK _3426_/D vssd1 vssd1 vccd1 vccd1 _3426_/Q sky130_fd_sc_hd__dfxtp_1
X_3357_ _3460_/CLK _3357_/D vssd1 vssd1 vccd1 vccd1 _3357_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _1960_/C _2283_/X _2307_/Y vssd1 vssd1 vccd1 vccd1 _2308_/Y sky130_fd_sc_hd__o21ai_2
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1999__A _1999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3288_ _3288_/CLK _3288_/D vssd1 vssd1 vccd1 vccd1 _3288_/Q sky130_fd_sc_hd__dfxtp_1
X_2239_ _2326_/A vssd1 vssd1 vccd1 vccd1 _2239_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2623__A _2660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input259_A ram_imem_response_put[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input161_A fmc_dmem_response_put[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input22_A core_dmem_request_put[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1702__A _1702_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output380_A _1939_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1610_ _1591_/X _1597_/X _3215_/Q vssd1 vssd1 vccd1 vccd1 _1610_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_output478_A _1448_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput507 _2277_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[32] sky130_fd_sc_hd__buf_2
Xoutput518 _2306_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[42] sky130_fd_sc_hd__buf_2
XFILLER_5_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2590_ _2466_/X _3156_/Q _2541_/A vssd1 vssd1 vccd1 vccd1 _2590_/X sky130_fd_sc_hd__o21ba_1
Xoutput529 _2335_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[52] sky130_fd_sc_hd__buf_2
X_1541_ _1541_/A vssd1 vssd1 vccd1 vccd1 _1541_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1472_ _1472_/A vssd1 vssd1 vccd1 vccd1 _1473_/C sky130_fd_sc_hd__inv_2
X_3211_ _3222_/CLK _3211_/D vssd1 vssd1 vccd1 vccd1 _3211_/Q sky130_fd_sc_hd__dfxtp_1
X_3142_ _3140_/X _3142_/A2 _2538_/X _2539_/X _3141_/X vssd1 vssd1 vccd1 vccd1 _3477_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3073_ _3427_/Q _3065_/X _2373_/Y _3061_/X vssd1 vssd1 vccd1 vccd1 _3427_/D sky130_fd_sc_hd__o211a_1
XFILLER_54_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2024_ _2097_/A vssd1 vssd1 vccd1 vccd1 _2054_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2926_ _2945_/A vssd1 vssd1 vccd1 vccd1 _2926_/X sky130_fd_sc_hd__clkbuf_2
X_2857_ _3298_/Q _2849_/X _2845_/X _1942_/Y vssd1 vssd1 vccd1 vccd1 _3298_/D sky130_fd_sc_hd__o211a_1
X_1808_ _1832_/A _1840_/B _1808_/C vssd1 vssd1 vccd1 vccd1 _1808_/Y sky130_fd_sc_hd__nand3_1
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2788_ _2794_/A vssd1 vssd1 vccd1 vccd1 _2868_/A sky130_fd_sc_hd__buf_2
XFILLER_2_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1739_ _1713_/X _3249_/Q _1714_/X vssd1 vssd1 vccd1 vccd1 _1739_/X sky130_fd_sc_hd__o21ba_1
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3409_ _3457_/CLK _3409_/D vssd1 vssd1 vccd1 vccd1 _3409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1432__A _2725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2711_ _3212_/Q _2709_/X _1600_/Y _2710_/X vssd1 vssd1 vccd1 vccd1 _3212_/D sky130_fd_sc_hd__o211a_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2616__A_N _3130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2642_ _2677_/B vssd1 vssd1 vccd1 vccd1 _2642_/X sky130_fd_sc_hd__clkbuf_2
X_2573_ _2564_/X _3485_/Q _2572_/X vssd1 vssd1 vccd1 vccd1 _2573_/X sky130_fd_sc_hd__o21ba_1
Xoutput315 _2507_/X vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[7] sky130_fd_sc_hd__buf_2
Xoutput326 _1721_/X vssd1 vssd1 vccd1 vccd1 core_imem_response_get[17] sky130_fd_sc_hd__buf_2
Xoutput304 _2586_/Y vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[26] sky130_fd_sc_hd__buf_2
X_1524_ _3188_/Q _1514_/X _1523_/Y vssd1 vssd1 vccd1 vccd1 _1524_/X sky130_fd_sc_hd__o21a_2
Xoutput348 _1682_/Y vssd1 vssd1 vccd1 vccd1 core_imem_response_get[8] sky130_fd_sc_hd__buf_2
Xoutput337 _1760_/X vssd1 vssd1 vccd1 vccd1 core_imem_response_get[27] sky130_fd_sc_hd__buf_2
Xoutput359 _1867_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[18] sky130_fd_sc_hd__buf_2
X_1455_ _1455_/A vssd1 vssd1 vccd1 vccd1 _1456_/C sky130_fd_sc_hd__inv_2
XFILLER_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3125_ _2601_/X _3125_/A2 _2486_/X _2487_/X _3154_/A vssd1 vssd1 vccd1 vccd1 _3465_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2510__A2 _2510_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3056_ _1997_/C _3049_/X _3053_/X _2336_/Y vssd1 vssd1 vccd1 vccd1 _3414_/D sky130_fd_sc_hd__o211ai_1
XFILLER_55_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2007_ _2007_/A vssd1 vssd1 vccd1 vccd1 _2008_/C sky130_fd_sc_hd__inv_2
XFILLER_23_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2909_ _3325_/Q _2893_/X _2040_/Y vssd1 vssd1 vccd1 vccd1 _2910_/A sky130_fd_sc_hd__o21ai_1
XFILLER_86_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input124_A core_imem_request_put[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_CLK CLK vssd1 vssd1 vccd1 vccd1 clkbuf_0_CLK/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__1543__A3 _1533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2740__A2 _2740_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output510_A _2286_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3089__A _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2625_ _2677_/B vssd1 vssd1 vccd1 vccd1 _2658_/A sky130_fd_sc_hd__clkbuf_2
X_2556_ _2564_/A vssd1 vssd1 vccd1 vccd1 _2556_/X sky130_fd_sc_hd__clkbuf_1
X_1507_ _3183_/Q _1498_/X _1506_/Y vssd1 vssd1 vccd1 vccd1 _1507_/X sky130_fd_sc_hd__o21a_2
X_2487_ _2487_/A _2478_/X vssd1 vssd1 vccd1 vccd1 _2487_/X sky130_fd_sc_hd__or2b_1
X_1438_ _2725_/A _1447_/B _1438_/C vssd1 vssd1 vccd1 vccd1 _1438_/Y sky130_fd_sc_hd__nand3_2
XFILLER_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3108_ _2134_/C _3105_/X _3003_/A _2442_/Y vssd1 vssd1 vccd1 vccd1 _3452_/D sky130_fd_sc_hd__o211ai_1
XANTENNA__1503__C _1503_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3039_ _3067_/A vssd1 vssd1 vccd1 vccd1 _3039_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2183__B1 _2163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2722__A2 _1630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input241_A ram_dmem_response_put[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1413__C _1533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2238__A1 _1869_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2806__A _2864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1710__A _1710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput36 core_dmem_request_put[2] vssd1 vssd1 vccd1 vccd1 _1803_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput25 core_dmem_request_put[1] vssd1 vssd1 vccd1 vccd1 _1800_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput14 core_dmem_request_put[0] vssd1 vssd1 vccd1 vccd1 _1793_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2410__A1 _2091_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2961__A2 _2950_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput69 core_dmem_request_put[5] vssd1 vssd1 vccd1 vccd1 _1814_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput47 core_dmem_request_put[3] vssd1 vssd1 vccd1 vccd1 _1807_/A sky130_fd_sc_hd__clkbuf_1
Xinput58 core_dmem_request_put[4] vssd1 vssd1 vccd1 vccd1 _1810_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_output460_A _1497_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output558_A _2410_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2410_ _2091_/C _2397_/X _2409_/Y vssd1 vssd1 vccd1 vccd1 _2410_/Y sky130_fd_sc_hd__o21ai_4
X_3390_ _3394_/CLK _3390_/D vssd1 vssd1 vccd1 vccd1 _3390_/Q sky130_fd_sc_hd__dfxtp_1
X_2341_ _2370_/A vssd1 vssd1 vccd1 vccd1 _2341_/X sky130_fd_sc_hd__clkbuf_2
X_2272_ _2269_/X _2270_/X _2271_/X _1913_/C _2262_/X vssd1 vssd1 vccd1 vccd1 _2272_/Y
+ sky130_fd_sc_hd__o311ai_4
XFILLER_69_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3123__C1 _3154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1987_ _3310_/Q _1984_/X _1986_/Y vssd1 vssd1 vccd1 vccd1 _1987_/X sky130_fd_sc_hd__o21a_1
XFILLER_20_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2451__A _3091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2608_ input2/X _2682_/B vssd1 vssd1 vccd1 vccd1 _3143_/A sky130_fd_sc_hd__nand2b_2
X_2539_ _2539_/A _2513_/X vssd1 vssd1 vccd1 vccd1 _2539_/X sky130_fd_sc_hd__or2b_1
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2468__A1 _2462_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input191_A fmc_imem_response_put[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input52_A core_dmem_request_put[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2171__A3 _2179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1910_ _3289_/Q _1892_/X _1909_/Y vssd1 vssd1 vccd1 vccd1 _1910_/X sky130_fd_sc_hd__o21a_2
XFILLER_30_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2890_ _3315_/Q _2873_/X _2004_/Y vssd1 vssd1 vccd1 vccd1 _2891_/A sky130_fd_sc_hd__o21ai_1
X_1841_ _3271_/Q _1834_/X _1840_/Y vssd1 vssd1 vccd1 vccd1 _1841_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1772_ _2757_/A vssd1 vssd1 vccd1 vccd1 _1772_/X sky130_fd_sc_hd__clkbuf_2
X_3442_ _3448_/CLK _3442_/D vssd1 vssd1 vccd1 vccd1 _3442_/Q sky130_fd_sc_hd__dfxtp_1
X_3373_ _3461_/CLK _3373_/D vssd1 vssd1 vccd1 vccd1 _3373_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2324_ _2312_/X _2323_/X _3410_/Q vssd1 vssd1 vccd1 vccd1 _2324_/Y sky130_fd_sc_hd__o21ai_2
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2255_ _2370_/A vssd1 vssd1 vccd1 vccd1 _2255_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3111__A2 _2174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2186_ _2206_/A vssd1 vssd1 vccd1 vccd1 _2186_/X sky130_fd_sc_hd__buf_2
XFILLER_38_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_CLK clkbuf_2_3_0_CLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_0_CLK/X sky130_fd_sc_hd__clkbuf_2
XFILLER_25_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2689__A1 _1435_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput226 ram_dmem_response_put[24] vssd1 vssd1 vccd1 vccd1 _2577_/A sky130_fd_sc_hd__buf_2
Xinput215 ram_dmem_response_put[14] vssd1 vssd1 vccd1 vccd1 _2535_/A sky130_fd_sc_hd__buf_2
XFILLER_88_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput204 fmc_imem_response_put[4] vssd1 vssd1 vccd1 vccd1 _1663_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput237 ram_dmem_response_put[5] vssd1 vssd1 vccd1 vccd1 _2495_/A sky130_fd_sc_hd__buf_2
Xinput259 ram_imem_response_put[25] vssd1 vssd1 vccd1 vccd1 _1752_/A sky130_fd_sc_hd__clkbuf_2
Xinput248 ram_imem_response_put[15] vssd1 vssd1 vccd1 vccd1 _1710_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1898__C _1898_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input204_A fmc_imem_response_put[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2613__A1 _2601_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1419__B _1531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1435__A _1443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2040_ _2054_/A _2062_/B _2040_/C vssd1 vssd1 vccd1 vccd1 _2040_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__2301__B1 _1949_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2942_ _3342_/Q _2926_/X _2941_/X _2102_/Y vssd1 vssd1 vccd1 vccd1 _3342_/D sky130_fd_sc_hd__o211a_1
XFILLER_62_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2604__A1 _2601_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2873_ _2893_/A vssd1 vssd1 vccd1 vccd1 _2873_/X sky130_fd_sc_hd__clkbuf_2
X_1824_ _1832_/A _1840_/B _1824_/C vssd1 vssd1 vccd1 vccd1 _1824_/Y sky130_fd_sc_hd__nand3_1
X_1755_ _1755_/A _1644_/A vssd1 vssd1 vccd1 vccd1 _1755_/X sky130_fd_sc_hd__or2b_1
X_1686_ _1642_/X _2746_/A2 _1683_/X _1685_/X vssd1 vssd1 vccd1 vccd1 _1686_/X sky130_fd_sc_hd__a22o_1
X_3425_ _3449_/CLK _3425_/D vssd1 vssd1 vccd1 vccd1 _3425_/Q sky130_fd_sc_hd__dfxtp_1
X_3356_ _3356_/CLK _3356_/D vssd1 vssd1 vccd1 vccd1 _3356_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2307_ _2284_/X _2294_/X _3404_/Q vssd1 vssd1 vccd1 vccd1 _2307_/Y sky130_fd_sc_hd__o21ai_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _3288_/CLK _3287_/D vssd1 vssd1 vccd1 vccd1 _3287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2238_ _1869_/C _2224_/X _2237_/Y vssd1 vssd1 vccd1 vccd1 _2238_/Y sky130_fd_sc_hd__o21ai_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3096__A1 _2099_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2169_ _2169_/A vssd1 vssd1 vccd1 vccd1 _2169_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_26_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input154_A fmc_dmem_response_put[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input15_A core_dmem_request_put[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2086__A _2206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3011__A1 _1877_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output373_A _1914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput508 _2279_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[33] sky130_fd_sc_hd__buf_2
X_1540_ _1530_/X _2725_/B _1534_/X _1537_/X _3192_/Q vssd1 vssd1 vccd1 vccd1 _1540_/X
+ sky130_fd_sc_hd__o41a_4
Xoutput519 _2308_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[43] sky130_fd_sc_hd__buf_2
XFILLER_5_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1471_ _3173_/Q _1462_/X _1470_/Y vssd1 vssd1 vccd1 vccd1 _1471_/X sky130_fd_sc_hd__o21a_2
XFILLER_79_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3210_ _3222_/CLK _3210_/D vssd1 vssd1 vccd1 vccd1 _3210_/Q sky130_fd_sc_hd__dfxtp_1
X_3141_ _3143_/A vssd1 vssd1 vccd1 vccd1 _3141_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_79_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1638__B_N _1637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3078__A1 _2054_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3072_ _2040_/C _3063_/X _3067_/X _2371_/Y vssd1 vssd1 vccd1 vccd1 _3426_/D sky130_fd_sc_hd__o211ai_1
X_2023_ _3320_/Q _2020_/X _2022_/Y vssd1 vssd1 vccd1 vccd1 _2023_/X sky130_fd_sc_hd__o21a_1
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2925_ _2925_/A _2933_/B vssd1 vssd1 vccd1 vccd1 _3333_/D sky130_fd_sc_hd__nand2_1
X_2856_ _2856_/A _2856_/B vssd1 vssd1 vccd1 vccd1 _3297_/D sky130_fd_sc_hd__nand2_1
XANTENNA__3002__A1 _1862_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1807_ _1807_/A vssd1 vssd1 vccd1 vccd1 _1808_/C sky130_fd_sc_hd__inv_4
X_2787_ _2787_/A _2797_/B vssd1 vssd1 vccd1 vccd1 _3263_/D sky130_fd_sc_hd__nand2_1
X_1738_ _1734_/X _2762_/A2 _1736_/X _1737_/X vssd1 vssd1 vccd1 vccd1 _1738_/X sky130_fd_sc_hd__a22o_2
X_1669_ _1712_/A vssd1 vssd1 vccd1 vccd1 _1669_/X sky130_fd_sc_hd__buf_4
X_3408_ _3410_/CLK _3408_/D vssd1 vssd1 vccd1 vccd1 _3408_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1506__C _1506_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input7_A EN_fmc_imem_request_get vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _3440_/CLK _3339_/D vssd1 vssd1 vccd1 vccd1 _3339_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input271_A ram_imem_response_put[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1555__A1 _1429_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2710_ _2712_/A vssd1 vssd1 vccd1 vccd1 _2710_/X sky130_fd_sc_hd__clkbuf_2
X_2641_ _2660_/A vssd1 vssd1 vccd1 vccd1 _2641_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2572_ _2572_/A vssd1 vssd1 vccd1 vccd1 _2572_/X sky130_fd_sc_hd__clkbuf_2
Xoutput316 _2511_/Y vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[8] sky130_fd_sc_hd__buf_2
Xoutput305 _2589_/X vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[27] sky130_fd_sc_hd__buf_2
Xoutput349 _1686_/X vssd1 vssd1 vccd1 vccd1 core_imem_response_get[9] sky130_fd_sc_hd__buf_2
Xoutput338 _1764_/Y vssd1 vssd1 vccd1 vccd1 core_imem_response_get[28] sky130_fd_sc_hd__buf_2
Xoutput327 _1725_/Y vssd1 vssd1 vccd1 vccd1 core_imem_response_get[18] sky130_fd_sc_hd__buf_2
X_1523_ _1541_/A _1523_/B _1523_/C vssd1 vssd1 vccd1 vccd1 _1523_/Y sky130_fd_sc_hd__nand3_1
X_1454_ _2675_/B vssd1 vssd1 vccd1 vccd1 _1484_/B sky130_fd_sc_hd__clkbuf_2
X_3124_ _3126_/A _3124_/B vssd1 vssd1 vccd1 vccd1 _3464_/D sky130_fd_sc_hd__nor2_1
X_3055_ _3413_/Q _3051_/X _2334_/Y _3047_/X vssd1 vssd1 vccd1 vccd1 _3413_/D sky130_fd_sc_hd__o211a_1
XFILLER_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2006_ _2006_/A vssd1 vssd1 vccd1 vccd1 _2036_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2908_ _3324_/Q _2907_/X _2903_/X _2036_/Y vssd1 vssd1 vccd1 vccd1 _3324_/D sky130_fd_sc_hd__o211a_1
X_2839_ _3289_/Q _2835_/X _1909_/Y vssd1 vssd1 vccd1 vccd1 _2841_/A sky130_fd_sc_hd__o21ai_1
XFILLER_2_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1533__A _1533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input117_A core_imem_request_put[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input82_A core_dmem_request_put[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2539__A _2539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1443__A _1443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output503_A _2267_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1767__A1 _1734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2624_ _3162_/Q _2623_/X _1429_/Y vssd1 vssd1 vccd1 vccd1 _2627_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__2192__A1 _1808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2555_ _2521_/X _3481_/Q _2529_/X vssd1 vssd1 vccd1 vccd1 _2555_/X sky130_fd_sc_hd__o21ba_1
X_1506_ _1512_/A _1520_/B _1506_/C vssd1 vssd1 vccd1 vccd1 _1506_/Y sky130_fd_sc_hd__nand3_1
X_2486_ _2473_/X _3465_/Q _2485_/X vssd1 vssd1 vccd1 vccd1 _2486_/X sky130_fd_sc_hd__o21ba_1
XFILLER_68_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1437_ _1437_/A vssd1 vssd1 vccd1 vccd1 _1438_/C sky130_fd_sc_hd__clkinv_4
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3107_ _3451_/Q _2174_/A _2440_/Y _3103_/X vssd1 vssd1 vccd1 vccd1 _3451_/D sky130_fd_sc_hd__o211a_1
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3038_ _3401_/Q _3037_/X _2301_/Y _3033_/X vssd1 vssd1 vccd1 vccd1 _3401_/D sky130_fd_sc_hd__o211a_1
XFILLER_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2912__A _2950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2183__A1 _2175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input234_A ram_dmem_response_put[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2094__A _2094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput37 core_dmem_request_put[30] vssd1 vssd1 vccd1 vccd1 _1912_/A sky130_fd_sc_hd__clkbuf_1
Xinput15 core_dmem_request_put[10] vssd1 vssd1 vccd1 vccd1 _1835_/A sky130_fd_sc_hd__clkbuf_1
Xinput26 core_dmem_request_put[20] vssd1 vssd1 vccd1 vccd1 _1872_/A sky130_fd_sc_hd__clkbuf_1
Xinput48 core_dmem_request_put[40] vssd1 vssd1 vccd1 vccd1 _1948_/A sky130_fd_sc_hd__clkbuf_1
Xinput59 core_dmem_request_put[50] vssd1 vssd1 vccd1 vccd1 _1985_/A sky130_fd_sc_hd__buf_2
XANTENNA__1438__A _2725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output453_A _1471_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2340_ _2397_/A vssd1 vssd1 vccd1 vccd1 _2340_/X sky130_fd_sc_hd__buf_2
X_2271_ _2300_/A vssd1 vssd1 vccd1 vccd1 _2271_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_77_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1986_ _2000_/A _2008_/B _1986_/C vssd1 vssd1 vccd1 vccd1 _1986_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__2732__A _2760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2607_ _2975_/B vssd1 vssd1 vccd1 vccd1 _2682_/B sky130_fd_sc_hd__buf_4
XANTENNA__2968__B1_N _2959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2538_ _2521_/X _3477_/Q _2529_/X vssd1 vssd1 vccd1 vccd1 _2538_/X sky130_fd_sc_hd__o21ba_1
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2179__A _2179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2469_ _3122_/B vssd1 vssd1 vccd1 vccd1 _2469_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2468__A2 _2468_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2907__A _2945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1811__A _3116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2642__A _2677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1600__B1 _1492_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input184_A fmc_imem_response_put[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input45_A core_dmem_request_put[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1840_ _1869_/A _1840_/B _1840_/C vssd1 vssd1 vccd1 vccd1 _1840_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__2552__A _2552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1771_ _2771_/B vssd1 vssd1 vccd1 vccd1 _1771_/Y sky130_fd_sc_hd__inv_2
X_3441_ _3447_/CLK _3441_/D vssd1 vssd1 vccd1 vccd1 _3441_/Q sky130_fd_sc_hd__dfxtp_1
X_3372_ _3372_/CLK _3372_/D vssd1 vssd1 vccd1 vccd1 _3372_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2323_ _2351_/A vssd1 vssd1 vccd1 vccd1 _2323_/X sky130_fd_sc_hd__clkbuf_2
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2254_ _2427_/A vssd1 vssd1 vccd1 vccd1 _2370_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2185_ _2253_/A vssd1 vssd1 vccd1 vccd1 _2185_/X sky130_fd_sc_hd__buf_2
XFILLER_65_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1830__B1 _1829_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1969_ _2006_/A vssd1 vssd1 vccd1 vccd1 _2000_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1509__C _1509_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1806__A _2408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput227 ram_dmem_response_put[25] vssd1 vssd1 vccd1 vccd1 _2581_/A sky130_fd_sc_hd__clkbuf_4
Xinput216 ram_dmem_response_put[15] vssd1 vssd1 vccd1 vccd1 _2539_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput205 fmc_imem_response_put[5] vssd1 vssd1 vccd1 vccd1 _2740_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput238 ram_dmem_response_put[6] vssd1 vssd1 vccd1 vccd1 _2502_/A sky130_fd_sc_hd__buf_2
Xinput249 ram_imem_response_put[16] vssd1 vssd1 vccd1 vccd1 _1716_/A sky130_fd_sc_hd__buf_2
XFILLER_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2613__A2 _2613_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1419__C _1533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1716__A _1716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1435__B _1452_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2941_ _2969_/B vssd1 vssd1 vccd1 vccd1 _2941_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2604__A2 _2615_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2872_ _3306_/Q _2868_/X _2864_/X _1971_/Y vssd1 vssd1 vccd1 vccd1 _3306_/D sky130_fd_sc_hd__o211a_1
XFILLER_30_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1823_ _1823_/A vssd1 vssd1 vccd1 vccd1 _1824_/C sky130_fd_sc_hd__inv_4
X_1754_ _1637_/X _3253_/Q _1712_/A vssd1 vssd1 vccd1 vccd1 _1754_/X sky130_fd_sc_hd__o21ba_1
XFILLER_7_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3424_ _3452_/CLK _3424_/D vssd1 vssd1 vccd1 vccd1 _3424_/Q sky130_fd_sc_hd__dfxtp_1
X_1685_ _1685_/A _1684_/X vssd1 vssd1 vccd1 vccd1 _1685_/X sky130_fd_sc_hd__or2b_1
X_3355_ _3454_/CLK _3355_/D vssd1 vssd1 vccd1 vccd1 _3355_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ _3403_/Q _2297_/X _2305_/Y vssd1 vssd1 vccd1 vccd1 _2306_/X sky130_fd_sc_hd__o21a_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _3486_/CLK _3286_/D vssd1 vssd1 vccd1 vccd1 _3286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2237_ _2225_/X _2236_/X _3380_/Q vssd1 vssd1 vccd1 vccd1 _2237_/Y sky130_fd_sc_hd__o21ai_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2168_ _2156_/X _3116_/B _2162_/X _2165_/X _3359_/Q vssd1 vssd1 vccd1 vccd1 _2168_/X
+ sky130_fd_sc_hd__o41a_2
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2099_ _2127_/A _2099_/B _2099_/C vssd1 vssd1 vccd1 vccd1 _2099_/Y sky130_fd_sc_hd__nand3_1
XFILLER_80_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input147_A fmc_dmem_response_put[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2830__A _2868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput509 _2281_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[34] sky130_fd_sc_hd__buf_2
XFILLER_8_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_CLK clkbuf_2_1_0_CLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_CLK/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_output366_A _1889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1470_ _1476_/A _1484_/B _1470_/C vssd1 vssd1 vccd1 vccd1 _1470_/Y sky130_fd_sc_hd__nand3_1
XFILLER_67_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3140_ _3140_/A vssd1 vssd1 vccd1 vccd1 _3140_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3071_ _3425_/Q _3065_/X _2367_/Y _3061_/X vssd1 vssd1 vccd1 vccd1 _3425_/D sky130_fd_sc_hd__o211a_1
X_2022_ _2036_/A _2044_/B _2022_/C vssd1 vssd1 vccd1 vccd1 _2022_/Y sky130_fd_sc_hd__nand3_1
XFILLER_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2924_ _3333_/Q _2912_/X _2069_/Y vssd1 vssd1 vccd1 vccd1 _2925_/A sky130_fd_sc_hd__o21ai_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2855_ _3297_/Q _2854_/X _1938_/Y vssd1 vssd1 vccd1 vccd1 _2856_/A sky130_fd_sc_hd__o21ai_1
X_1806_ _2408_/A vssd1 vssd1 vccd1 vccd1 _1840_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_2786_ _3263_/Q _2779_/X _1808_/Y vssd1 vssd1 vccd1 vccd1 _2787_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__1564__A2 _1527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1737_ _1737_/A _1727_/X vssd1 vssd1 vccd1 vccd1 _1737_/X sky130_fd_sc_hd__or2b_1
X_1668_ input8/X vssd1 vssd1 vccd1 vccd1 _1712_/A sky130_fd_sc_hd__clkbuf_2
X_3407_ _3457_/CLK _3407_/D vssd1 vssd1 vccd1 vccd1 _3407_/Q sky130_fd_sc_hd__dfxtp_1
X_3338_ _3447_/CLK _3338_/D vssd1 vssd1 vccd1 vccd1 _3338_/Q sky130_fd_sc_hd__dfxtp_1
X_1599_ _1488_/C _1590_/X _1598_/Y vssd1 vssd1 vccd1 vccd1 _1599_/Y sky130_fd_sc_hd__o21ai_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3269_ _3360_/CLK _3269_/D vssd1 vssd1 vccd1 vccd1 _3269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input264_A ram_imem_response_put[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1432__C _1432_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2440__B1 _2131_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2640_ _2640_/A _2655_/B vssd1 vssd1 vccd1 vccd1 _3170_/D sky130_fd_sc_hd__nand2_1
XANTENNA__2560__A _2560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_45_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3477_/CLK sky130_fd_sc_hd__clkbuf_16
X_2571_ _3150_/B vssd1 vssd1 vccd1 vccd1 _2571_/Y sky130_fd_sc_hd__inv_2
Xoutput317 _2515_/X vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[9] sky130_fd_sc_hd__buf_2
Xoutput306 _2593_/Y vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[28] sky130_fd_sc_hd__buf_2
Xoutput339 _1767_/X vssd1 vssd1 vccd1 vccd1 core_imem_response_get[29] sky130_fd_sc_hd__buf_2
Xoutput328 _1729_/X vssd1 vssd1 vccd1 vccd1 core_imem_response_get[19] sky130_fd_sc_hd__buf_2
X_1522_ _1522_/A vssd1 vssd1 vccd1 vccd1 _1523_/C sky130_fd_sc_hd__clkinv_4
X_1453_ _3168_/Q _1441_/X _1452_/Y vssd1 vssd1 vccd1 vccd1 _1453_/X sky130_fd_sc_hd__o21a_2
XANTENNA__1904__A _2049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3123_ _2601_/X _3123_/A2 _2476_/X _2479_/X _3154_/A vssd1 vssd1 vccd1 vccd1 _3463_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1755__B_N _1644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3054_ _1990_/C _3049_/X _3053_/X _2332_/Y vssd1 vssd1 vccd1 vccd1 _3412_/D sky130_fd_sc_hd__o211ai_1
XFILLER_82_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2735__A _2760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2005_ _3315_/Q _2002_/X _2004_/Y vssd1 vssd1 vccd1 vccd1 _2005_/X sky130_fd_sc_hd__o21a_2
XFILLER_63_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2907_ _2945_/A vssd1 vssd1 vccd1 vccd1 _2907_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_36_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3360_/CLK sky130_fd_sc_hd__clkbuf_16
X_2838_ _3288_/Q _2830_/X _2826_/X _1906_/Y vssd1 vssd1 vccd1 vccd1 _3288_/D sky130_fd_sc_hd__o211a_1
X_2769_ _2769_/A _2769_/B vssd1 vssd1 vccd1 vccd1 _3255_/D sky130_fd_sc_hd__nor2_1
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2380__A _2408_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3456_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_input75_A core_dmem_request_put[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1528__A2 _1514_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output329_A _1651_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1443__B _1452_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1767__A2 _2770_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3413_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2623_ _2660_/A vssd1 vssd1 vccd1 vccd1 _2623_/X sky130_fd_sc_hd__clkbuf_2
X_2554_ _3146_/B vssd1 vssd1 vccd1 vccd1 _2554_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2192__A2 _2185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1505_ _1505_/A vssd1 vssd1 vccd1 vccd1 _1506_/C sky130_fd_sc_hd__inv_2
X_2485_ _2572_/A vssd1 vssd1 vccd1 vccd1 _2485_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1634__A _1776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1436_ _3164_/Q _1415_/X _1435_/Y vssd1 vssd1 vccd1 vccd1 _1436_/X sky130_fd_sc_hd__o21a_2
XFILLER_68_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3106_ _2127_/C _3105_/X _3095_/X _2437_/Y vssd1 vssd1 vccd1 vccd1 _3450_/D sky130_fd_sc_hd__o211ai_1
XFILLER_28_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3037_ _3037_/A vssd1 vssd1 vccd1 vccd1 _3037_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2183__A2 _2177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1544__A _2709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input227_A ram_dmem_response_put[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput16 core_dmem_request_put[11] vssd1 vssd1 vccd1 vccd1 _1839_/A sky130_fd_sc_hd__clkbuf_1
Xinput27 core_dmem_request_put[21] vssd1 vssd1 vccd1 vccd1 _1876_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__1749__A2 _1749_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput49 core_dmem_request_put[41] vssd1 vssd1 vccd1 vccd1 _1952_/A sky130_fd_sc_hd__clkbuf_1
Xinput38 core_dmem_request_put[31] vssd1 vssd1 vccd1 vccd1 _1916_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_output279_A _3490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output446_A _2166_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1454__A _2675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2270_ _2299_/A vssd1 vssd1 vccd1 vccd1 _2270_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3123__A1 _2601_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_7_CLK clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3372_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_65_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1985_ _1985_/A vssd1 vssd1 vccd1 vccd1 _1986_/C sky130_fd_sc_hd__inv_2
XFILLER_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2606_ _2606_/A vssd1 vssd1 vccd1 vccd1 _2616_/B sky130_fd_sc_hd__clkbuf_1
X_2537_ _3139_/B vssd1 vssd1 vccd1 vccd1 _2537_/Y sky130_fd_sc_hd__inv_2
X_2468_ _2462_/X _2468_/A2 _2465_/X _2467_/X vssd1 vssd1 vccd1 vccd1 _3122_/B sky130_fd_sc_hd__a22oi_2
X_1419_ _1529_/A _1531_/A _1533_/A vssd1 vssd1 vccd1 vccd1 _1426_/A sky130_fd_sc_hd__nor3_1
X_2399_ _2398_/X _2380_/X _3436_/Q vssd1 vssd1 vccd1 vccd1 _2399_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input177_A fmc_dmem_response_put[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input38_A core_dmem_request_put[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output396_A _1991_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1770_ _1691_/A _1770_/A2 _1768_/X _1769_/X vssd1 vssd1 vccd1 vccd1 _2771_/B sky130_fd_sc_hd__a22oi_4
XANTENNA_output563_A _2422_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3440_ _3440_/CLK _3440_/D vssd1 vssd1 vccd1 vccd1 _3440_/Q sky130_fd_sc_hd__dfxtp_1
X_3371_ _3397_/CLK _3371_/D vssd1 vssd1 vccd1 vccd1 _3371_/Q sky130_fd_sc_hd__dfxtp_1
X_2322_ _3409_/Q _2297_/X _2321_/Y vssd1 vssd1 vccd1 vccd1 _2322_/X sky130_fd_sc_hd__o21a_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2253_ _2253_/A vssd1 vssd1 vccd1 vccd1 _2253_/X sky130_fd_sc_hd__buf_2
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2184_ _3105_/A vssd1 vssd1 vccd1 vccd1 _2253_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1968_ _3305_/Q _1965_/X _1967_/Y vssd1 vssd1 vccd1 vccd1 _1968_/X sky130_fd_sc_hd__o21a_2
X_1899_ _3286_/Q _1892_/X _1898_/Y vssd1 vssd1 vccd1 vccd1 _1899_/X sky130_fd_sc_hd__o21a_2
XFILLER_88_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput217 ram_dmem_response_put[16] vssd1 vssd1 vccd1 vccd1 _2545_/A sky130_fd_sc_hd__buf_2
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput206 fmc_imem_response_put[6] vssd1 vssd1 vccd1 vccd1 _1674_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput228 ram_dmem_response_put[26] vssd1 vssd1 vccd1 vccd1 _2584_/A sky130_fd_sc_hd__buf_2
Xinput239 ram_dmem_response_put[7] vssd1 vssd1 vccd1 vccd1 _2506_/A sky130_fd_sc_hd__buf_2
XFILLER_75_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2091__C _2091_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1435__C _1435_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output409_A _2034_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2940_ _2940_/A _2952_/B vssd1 vssd1 vccd1 vccd1 _3341_/D sky130_fd_sc_hd__nand2_1
X_2871_ _2871_/A _2875_/B vssd1 vssd1 vccd1 vccd1 _3305_/D sky130_fd_sc_hd__nand2_1
XFILLER_15_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1822_ _3266_/Q _1813_/X _1821_/Y vssd1 vssd1 vccd1 vccd1 _1822_/X sky130_fd_sc_hd__o21a_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1753_ _1734_/X _2766_/A2 _1751_/X _1752_/X vssd1 vssd1 vccd1 vccd1 _1753_/X sky130_fd_sc_hd__a22o_1
X_1684_ _1735_/A vssd1 vssd1 vccd1 vccd1 _1684_/X sky130_fd_sc_hd__clkbuf_1
X_3423_ _3449_/CLK _3423_/D vssd1 vssd1 vccd1 vccd1 _3423_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _3356_/CLK _3354_/D vssd1 vssd1 vccd1 vccd1 _3354_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _2298_/X _2299_/X _2300_/X _1956_/C _2291_/X vssd1 vssd1 vccd1 vccd1 _2305_/Y
+ sky130_fd_sc_hd__o311ai_2
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2540__A2 _3142_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3285_ _3288_/CLK _3285_/D vssd1 vssd1 vccd1 vccd1 _3285_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1642__A _1691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2236_ _2351_/A vssd1 vssd1 vccd1 vccd1 _2236_/X sky130_fd_sc_hd__clkbuf_2
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2167_ _2156_/X _3116_/B _2162_/X _2165_/X _3358_/Q vssd1 vssd1 vccd1 vccd1 _2167_/X
+ sky130_fd_sc_hd__o41a_2
XFILLER_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2098_ _2098_/A vssd1 vssd1 vccd1 vccd1 _2099_/C sky130_fd_sc_hd__inv_2
XANTENNA__2473__A _2473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1567__B1 _1447_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1817__A _2163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2383__A _2459_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2770__A2 _2770_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3070_ _2033_/C _3063_/X _3067_/X _2365_/Y vssd1 vssd1 vccd1 vccd1 _3424_/D sky130_fd_sc_hd__o211ai_1
XFILLER_94_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2021_ _2021_/A vssd1 vssd1 vccd1 vccd1 _2022_/C sky130_fd_sc_hd__clkinv_2
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2286__A1 _1931_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2589__A2 _3155_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2923_ _3332_/Q _2907_/X _2922_/X _2065_/Y vssd1 vssd1 vccd1 vccd1 _3332_/D sky130_fd_sc_hd__o211a_1
X_2854_ _2893_/A vssd1 vssd1 vccd1 vccd1 _2854_/X sky130_fd_sc_hd__clkbuf_2
X_1805_ _3262_/Q _1784_/X _1804_/Y vssd1 vssd1 vccd1 vccd1 _1805_/X sky130_fd_sc_hd__o21a_1
X_2785_ _3262_/Q _2145_/X _2784_/X _1804_/Y vssd1 vssd1 vccd1 vccd1 _3262_/D sky130_fd_sc_hd__o211a_1
XANTENNA__1549__B1 _1423_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1637__A _1776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1736_ _1735_/X _3248_/Q _1700_/X vssd1 vssd1 vccd1 vccd1 _1736_/X sky130_fd_sc_hd__o21ba_1
XFILLER_7_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1667_ _1642_/X _2740_/A2 _1665_/X _1666_/X vssd1 vssd1 vccd1 vccd1 _1667_/X sky130_fd_sc_hd__a22o_1
X_1598_ _1591_/X _1597_/X _3211_/Q vssd1 vssd1 vccd1 vccd1 _1598_/Y sky130_fd_sc_hd__o21ai_1
X_3406_ _3410_/CLK _3406_/D vssd1 vssd1 vccd1 vccd1 _3406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3337_ _3337_/CLK _3337_/D vssd1 vssd1 vccd1 vccd1 _3337_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _3337_/CLK _3268_/D vssd1 vssd1 vccd1 vccd1 _3268_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2219_ _3373_/Q _2210_/X _2218_/Y vssd1 vssd1 vccd1 vccd1 _2219_/X sky130_fd_sc_hd__o21a_1
XFILLER_66_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3199_ _3226_/CLK _3199_/D vssd1 vssd1 vccd1 vccd1 _3199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2931__A _2950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input257_A ram_imem_response_put[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input20_A core_dmem_request_put[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output476_A _1439_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput307 _2596_/X vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[29] sky130_fd_sc_hd__buf_2
X_2570_ _2541_/X _2570_/A2 _2568_/X _2569_/X vssd1 vssd1 vccd1 vccd1 _3150_/B sky130_fd_sc_hd__a22oi_4
X_1521_ _3187_/Q _1514_/X _1520_/Y vssd1 vssd1 vccd1 vccd1 _1521_/X sky130_fd_sc_hd__o21a_2
Xoutput318 _1640_/Y vssd1 vssd1 vccd1 vccd1 core_imem_response_get[0] sky130_fd_sc_hd__buf_2
Xoutput329 _1651_/X vssd1 vssd1 vccd1 vccd1 core_imem_response_get[1] sky130_fd_sc_hd__buf_2
XFILLER_4_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1452_ _1480_/A _1452_/B _1452_/C vssd1 vssd1 vccd1 vccd1 _1452_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__3153__C1 _3130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3122_ _3126_/A _3122_/B vssd1 vssd1 vccd1 vccd1 _3462_/D sky130_fd_sc_hd__nor2_1
XFILLER_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3053_ _3067_/A vssd1 vssd1 vccd1 vccd1 _3053_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2482__B_N _2466_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2004_ _2018_/A _2026_/B _2004_/C vssd1 vssd1 vccd1 vccd1 _2004_/Y sky130_fd_sc_hd__nand3_1
XFILLER_50_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2906_ _2906_/A _2914_/B vssd1 vssd1 vccd1 vccd1 _3323_/D sky130_fd_sc_hd__nand2_1
X_2837_ _2837_/A _2837_/B vssd1 vssd1 vccd1 vccd1 _3287_/D sky130_fd_sc_hd__nand2_1
X_2768_ _2757_/X _2768_/A2 _1758_/X _1759_/X _2758_/X vssd1 vssd1 vccd1 vccd1 _3254_/D
+ sky130_fd_sc_hd__a221o_1
X_2699_ _1460_/C _2693_/X _2698_/X _1574_/Y vssd1 vssd1 vccd1 vccd1 _3203_/D sky130_fd_sc_hd__o211ai_1
XFILLER_2_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1719_ _1692_/X _3244_/Q _1700_/X vssd1 vssd1 vccd1 vccd1 _1719_/X sky130_fd_sc_hd__o21ba_1
XFILLER_76_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2926__A _2945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_2_0_0_CLK clkbuf_2_1_0_CLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_0_CLK/X sky130_fd_sc_hd__clkbuf_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2661__A _2677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input68_A core_dmem_request_put[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2489__A1 _2464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1443__C _1443_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1740__A _1740_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output593_A _1555_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2964__A2 _2950_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1621__C1 _1443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2622_ _3161_/Q _2619_/X _2621_/X _1423_/Y vssd1 vssd1 vccd1 vccd1 _3161_/D sky130_fd_sc_hd__o211a_1
X_2553_ _2541_/X _2553_/A2 _2551_/X _2552_/X vssd1 vssd1 vccd1 vccd1 _3146_/B sky130_fd_sc_hd__a22oi_4
XANTENNA__1915__A _1951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1504_ _3182_/Q _1498_/X _1503_/Y vssd1 vssd1 vccd1 vccd1 _1504_/X sky130_fd_sc_hd__o21a_2
X_2484_ _3124_/B vssd1 vssd1 vccd1 vccd1 _2484_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1435_ _1443_/A _1452_/B _1435_/C vssd1 vssd1 vccd1 vccd1 _1435_/Y sky130_fd_sc_hd__nand3_1
XFILLER_95_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3105_ _3105_/A vssd1 vssd1 vccd1 vccd1 _3105_/X sky130_fd_sc_hd__buf_2
XFILLER_55_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3036_ _1945_/C _3035_/X _3025_/X _2295_/Y vssd1 vssd1 vccd1 vccd1 _3400_/D sky130_fd_sc_hd__o211ai_1
XANTENNA__1650__A _1650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2183__A3 _2179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3132__A2 _3132_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input122_A core_imem_request_put[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput17 core_dmem_request_put[12] vssd1 vssd1 vccd1 vccd1 _1842_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput28 core_dmem_request_put[22] vssd1 vssd1 vccd1 vccd1 _1879_/A sky130_fd_sc_hd__clkbuf_1
Xinput39 core_dmem_request_put[32] vssd1 vssd1 vccd1 vccd1 _1919_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__1438__C _1438_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3123__A2 _3123_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2566__A _2566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output606_A _1629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1901__C _1901_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1984_ _2056_/A vssd1 vssd1 vccd1 vccd1 _1984_/X sky130_fd_sc_hd__buf_2
XFILLER_9_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2605_ _3160_/Q _2605_/B input6/X vssd1 vssd1 vccd1 vccd1 _2606_/A sky130_fd_sc_hd__or3_1
XANTENNA__1645__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2536_ _2498_/X _2536_/A2 _2533_/X _2535_/X vssd1 vssd1 vccd1 vccd1 _3139_/B sky130_fd_sc_hd__a22oi_4
X_2467_ _2467_/A _2466_/X vssd1 vssd1 vccd1 vccd1 _2467_/X sky130_fd_sc_hd__or2b_1
X_1418_ _1541_/A vssd1 vssd1 vccd1 vccd1 _2725_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2398_ _2427_/A vssd1 vssd1 vccd1 vccd1 _2398_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1811__C _1811_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3019_ _3075_/A vssd1 vssd1 vccd1 vccd1 _3019_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3050__A1 _1981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1781__D_N input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput490 _2231_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[17] sky130_fd_sc_hd__buf_2
XFILLER_93_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1667__A2 _2740_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2092__A2 _2075_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3010__A _3067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output389_A _1968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output556_A _2404_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3370_ _3372_/CLK _3370_/D vssd1 vssd1 vccd1 vccd1 _3370_/Q sky130_fd_sc_hd__dfxtp_1
X_2321_ _2298_/X _2299_/X _2300_/X _1978_/C _2320_/X vssd1 vssd1 vccd1 vccd1 _2321_/Y
+ sky130_fd_sc_hd__o311ai_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2252_ _3385_/Q _2239_/X _2251_/Y vssd1 vssd1 vccd1 vccd1 _2252_/X sky130_fd_sc_hd__o21a_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2183_ _2175_/A _2177_/A _2179_/A _2163_/A vssd1 vssd1 vccd1 vccd1 _3105_/A sky130_fd_sc_hd__o31ai_4
XFILLER_38_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3032__A1 _1938_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1967_ _1981_/A _1990_/B _1967_/C vssd1 vssd1 vccd1 vccd1 _1967_/Y sky130_fd_sc_hd__nand3_1
X_1898_ _1927_/A _1898_/B _1898_/C vssd1 vssd1 vccd1 vccd1 _1898_/Y sky130_fd_sc_hd__nand3_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2519_ _3135_/B vssd1 vssd1 vccd1 vccd1 _2519_/Y sky130_fd_sc_hd__inv_2
Xinput218 ram_dmem_response_put[17] vssd1 vssd1 vccd1 vccd1 _2549_/A sky130_fd_sc_hd__clkbuf_4
Xinput207 fmc_imem_response_put[7] vssd1 vssd1 vccd1 vccd1 _2742_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput229 ram_dmem_response_put[27] vssd1 vssd1 vccd1 vccd1 _2588_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_75_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_51_CLK_A clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input50_A core_dmem_request_put[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_19_CLK_A clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3005__A _3035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2870_ _3305_/Q _2854_/X _1967_/Y vssd1 vssd1 vccd1 vccd1 _2871_/A sky130_fd_sc_hd__o21ai_1
XFILLER_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1821_ _1850_/A _1821_/B _1821_/C vssd1 vssd1 vccd1 vccd1 _1821_/Y sky130_fd_sc_hd__nand3_2
XFILLER_90_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1752_ _1752_/A _1727_/X vssd1 vssd1 vccd1 vccd1 _1752_/X sky130_fd_sc_hd__or2b_1
X_1683_ _1644_/X _3236_/Q _1656_/X vssd1 vssd1 vccd1 vccd1 _1683_/X sky130_fd_sc_hd__o21ba_1
X_3422_ _3452_/CLK _3422_/D vssd1 vssd1 vccd1 vccd1 _3422_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _3454_/CLK _3353_/D vssd1 vssd1 vccd1 vccd1 _3353_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ _1953_/C _2283_/X _2303_/Y vssd1 vssd1 vccd1 vccd1 _2304_/Y sky130_fd_sc_hd__o21ai_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _3288_/CLK _3284_/D vssd1 vssd1 vccd1 vccd1 _3284_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2235_ _2235_/A vssd1 vssd1 vccd1 vccd1 _2351_/A sky130_fd_sc_hd__buf_2
X_2166_ _2156_/X _3116_/B _2162_/X _2165_/X _3357_/Q vssd1 vssd1 vccd1 vccd1 _2166_/X
+ sky130_fd_sc_hd__o41a_2
XFILLER_38_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2097_ _2097_/A vssd1 vssd1 vccd1 vccd1 _2127_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2999_ _3375_/Q _2993_/X _2222_/Y _2989_/X vssd1 vssd1 vccd1 vccd1 _3375_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input202_A fmc_imem_response_put[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input98_A core_dmem_request_put[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output519_A _2308_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2020_ _2056_/A vssd1 vssd1 vccd1 vccd1 _2020_/X sky130_fd_sc_hd__buf_2
XFILLER_10_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2574__A _2574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2922_ _2969_/B vssd1 vssd1 vccd1 vccd1 _2922_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2853_ _3296_/Q _2849_/X _2845_/X _1935_/Y vssd1 vssd1 vccd1 vccd1 _3296_/D sky130_fd_sc_hd__o211a_1
X_1804_ _3116_/A _1821_/B _1804_/C vssd1 vssd1 vccd1 vccd1 _1804_/Y sky130_fd_sc_hd__nand3_2
X_2784_ _2864_/A vssd1 vssd1 vccd1 vccd1 _2784_/X sky130_fd_sc_hd__clkbuf_2
X_1735_ _1735_/A vssd1 vssd1 vccd1 vccd1 _1735_/X sky130_fd_sc_hd__buf_2
X_1666_ _1666_/A _1649_/X vssd1 vssd1 vccd1 vccd1 _1666_/X sky130_fd_sc_hd__or2b_1
X_3405_ _3457_/CLK _3405_/D vssd1 vssd1 vccd1 vccd1 _3405_/Q sky130_fd_sc_hd__dfxtp_1
X_1597_ _1597_/A vssd1 vssd1 vccd1 vccd1 _1597_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1653__A _1653_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3336_ _3447_/CLK _3336_/D vssd1 vssd1 vccd1 vccd1 _3336_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _3360_/CLK _3267_/D vssd1 vssd1 vccd1 vccd1 _3267_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2218_ _2211_/X _2212_/X _2213_/X _1843_/C _2203_/X vssd1 vssd1 vccd1 vccd1 _2218_/Y
+ sky130_fd_sc_hd__o311ai_2
X_3198_ _3226_/CLK _3198_/D vssd1 vssd1 vccd1 vccd1 _3198_/Q sky130_fd_sc_hd__dfxtp_1
X_2149_ _2319_/A vssd1 vssd1 vccd1 vccd1 _2291_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2201__A2 _2186_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input152_A fmc_dmem_response_put[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input13_A RST_N vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output371_A _1910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output469_A _1524_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput308 _2484_/Y vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[2] sky130_fd_sc_hd__buf_2
X_1520_ _1527_/A _1520_/B _1520_/C vssd1 vssd1 vccd1 vccd1 _1520_/Y sky130_fd_sc_hd__nand3_1
Xoutput319 _1690_/Y vssd1 vssd1 vccd1 vccd1 core_imem_response_get[10] sky130_fd_sc_hd__buf_2
X_1451_ _1451_/A vssd1 vssd1 vccd1 vccd1 _1452_/C sky130_fd_sc_hd__clkinv_4
XANTENNA__2569__A _2569_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1473__A _1480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3121_ _3461_/Q _2439_/X _2978_/X vssd1 vssd1 vccd1 vccd1 _3461_/D sky130_fd_sc_hd__o21a_1
X_3052_ _3411_/Q _3051_/X _2330_/Y _3047_/X vssd1 vssd1 vccd1 vccd1 _3411_/D sky130_fd_sc_hd__o211a_1
XFILLER_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2003_ _2003_/A vssd1 vssd1 vccd1 vccd1 _2004_/C sky130_fd_sc_hd__inv_2
XFILLER_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2905_ _3323_/Q _2893_/X _2033_/Y vssd1 vssd1 vccd1 vccd1 _2906_/A sky130_fd_sc_hd__o21ai_1
X_2836_ _3287_/Q _2835_/X _1901_/Y vssd1 vssd1 vccd1 vccd1 _2837_/A sky130_fd_sc_hd__o21ai_1
XFILLER_31_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1648__A _1776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2767_ _2769_/A _2767_/B vssd1 vssd1 vccd1 vccd1 _3253_/D sky130_fd_sc_hd__nor2_1
X_2698_ _2712_/A vssd1 vssd1 vccd1 vccd1 _2698_/X sky130_fd_sc_hd__clkbuf_2
X_1718_ _2754_/B vssd1 vssd1 vccd1 vccd1 _1718_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2479__A _2479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1649_ _1735_/A vssd1 vssd1 vccd1 vccd1 _1649_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input5_A EN_fmc_dmem_request_get vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ _3432_/CLK _3319_/D vssd1 vssd1 vccd1 vccd1 _3319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3103__A _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1621__B1 _1520_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2621_ _2677_/B vssd1 vssd1 vccd1 vccd1 _2621_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2552_ _2552_/A _2534_/X vssd1 vssd1 vccd1 vccd1 _2552_/X sky130_fd_sc_hd__or2b_1
X_1503_ _1516_/A _1523_/B _1503_/C vssd1 vssd1 vccd1 vccd1 _1503_/Y sky130_fd_sc_hd__nand3_1
X_2483_ _2462_/X _2483_/A2 _2481_/X _2482_/X vssd1 vssd1 vccd1 vccd1 _3124_/B sky130_fd_sc_hd__a22oi_2
XFILLER_87_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1434_ _1434_/A vssd1 vssd1 vccd1 vccd1 _1435_/C sky130_fd_sc_hd__clkinv_4
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3104_ _3449_/Q _3093_/X _2435_/Y _3103_/X vssd1 vssd1 vccd1 vccd1 _3449_/D sky130_fd_sc_hd__o211a_1
X_3035_ _3035_/A vssd1 vssd1 vccd1 vccd1 _3035_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1612__B1 _1506_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2819_ _3278_/Q _2810_/X _2806_/X _1866_/Y vssd1 vssd1 vccd1 vccd1 _3278_/D sky130_fd_sc_hd__o211a_1
XFILLER_11_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input115_A core_imem_request_put[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput18 core_dmem_request_put[13] vssd1 vssd1 vccd1 vccd1 _1846_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input80_A core_dmem_request_put[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput29 core_dmem_request_put[23] vssd1 vssd1 vccd1 vccd1 _1884_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__3108__B1 _3003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1983_ _2794_/A vssd1 vssd1 vccd1 vccd1 _2056_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2604_ _2601_/X _2615_/A2 _2602_/X _2603_/X vssd1 vssd1 vccd1 vccd1 _2604_/X sky130_fd_sc_hd__a22o_1
X_2535_ _2535_/A _2534_/X vssd1 vssd1 vccd1 vccd1 _2535_/X sky130_fd_sc_hd__or2b_1
XFILLER_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2466_ _2605_/B vssd1 vssd1 vccd1 vccd1 _2466_/X sky130_fd_sc_hd__buf_2
X_1417_ _1486_/A vssd1 vssd1 vccd1 vccd1 _1541_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2397_ _2397_/A vssd1 vssd1 vccd1 vccd1 _2397_/X sky130_fd_sc_hd__buf_4
XFILLER_83_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3018_ _3095_/A vssd1 vssd1 vccd1 vccd1 _3075_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2495__B_N _2478_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput480 _1457_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[8] sky130_fd_sc_hd__buf_2
Xoutput491 _2234_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[18] sky130_fd_sc_hd__buf_2
XANTENNA_input232_A ram_dmem_response_put[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output451_A _1465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2320_ _2434_/A vssd1 vssd1 vccd1 vccd1 _2320_/X sky130_fd_sc_hd__clkbuf_4
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2251_ _2240_/X _2241_/X _2242_/X _1888_/C _2232_/X vssd1 vssd1 vccd1 vccd1 _2251_/Y
+ sky130_fd_sc_hd__o311ai_2
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2577__A _2577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2304__A1 _1953_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2182_ _3361_/Q _2174_/X _2181_/Y vssd1 vssd1 vccd1 vccd1 _2182_/X sky130_fd_sc_hd__o21a_1
XFILLER_77_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1966_ _1966_/A vssd1 vssd1 vccd1 vccd1 _1967_/C sky130_fd_sc_hd__inv_2
X_1897_ _1897_/A vssd1 vssd1 vccd1 vccd1 _1898_/C sky130_fd_sc_hd__clkinv_4
X_2518_ _2498_/X _2518_/A2 _2516_/X _2517_/X vssd1 vssd1 vccd1 vccd1 _3135_/B sky130_fd_sc_hd__a22oi_4
XFILLER_0_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2487__A _2487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput208 fmc_imem_response_put[8] vssd1 vssd1 vccd1 vccd1 _1681_/A2 sky130_fd_sc_hd__clkbuf_4
X_2449_ _3455_/Q _2439_/X _2448_/Y vssd1 vssd1 vccd1 vccd1 _2449_/X sky130_fd_sc_hd__o21a_1
Xinput219 ram_dmem_response_put[18] vssd1 vssd1 vccd1 vccd1 _2552_/A sky130_fd_sc_hd__buf_2
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2950__A _2950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input182_A fmc_imem_response_put[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input43_A core_dmem_request_put[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2397__A _2397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3021__A _3035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1820_ _1820_/A vssd1 vssd1 vccd1 vccd1 _1821_/C sky130_fd_sc_hd__inv_6
XFILLER_30_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2222__B1 _1850_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1751_ _1735_/X _3252_/Q _1743_/X vssd1 vssd1 vccd1 vccd1 _1751_/X sky130_fd_sc_hd__o21ba_1
X_1682_ _2743_/B vssd1 vssd1 vccd1 vccd1 _1682_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3421_ _3457_/CLK _3421_/D vssd1 vssd1 vccd1 vccd1 _3421_/Q sky130_fd_sc_hd__dfxtp_1
X_3352_ _3454_/CLK _3352_/D vssd1 vssd1 vccd1 vccd1 _3352_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ _2284_/X _2294_/X _3402_/Q vssd1 vssd1 vccd1 vccd1 _2303_/Y sky130_fd_sc_hd__o21ai_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _3288_/CLK _3283_/D vssd1 vssd1 vccd1 vccd1 _3283_/Q sky130_fd_sc_hd__dfxtp_1
X_2234_ _3379_/Q _2210_/X _2233_/Y vssd1 vssd1 vccd1 vccd1 _2234_/X sky130_fd_sc_hd__o21a_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2165_ _2225_/A vssd1 vssd1 vccd1 vccd1 _2165_/X sky130_fd_sc_hd__buf_2
XFILLER_26_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2096_ _3340_/Q _2093_/X _2095_/Y vssd1 vssd1 vccd1 vccd1 _2096_/X sky130_fd_sc_hd__o21a_1
XFILLER_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2998_ _1847_/C _2991_/X _2995_/X _2220_/Y vssd1 vssd1 vccd1 vccd1 _3374_/D sky130_fd_sc_hd__o211ai_1
X_1949_ _1963_/A _1971_/B _1949_/C vssd1 vssd1 vccd1 vccd1 _1949_/Y sky130_fd_sc_hd__nand3_1
XFILLER_88_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2945__A _2945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2204__B1 _1829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1558__A2 _1527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2691__B1 _2686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2921_ _2921_/A _2933_/B vssd1 vssd1 vccd1 vccd1 _3331_/D sky130_fd_sc_hd__nand2_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_48_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3466_/CLK sky130_fd_sc_hd__clkbuf_16
X_2852_ _2852_/A _2856_/B vssd1 vssd1 vccd1 vccd1 _3295_/D sky130_fd_sc_hd__nand2_1
X_1803_ _1803_/A vssd1 vssd1 vccd1 vccd1 _1804_/C sky130_fd_sc_hd__inv_6
X_2783_ _2959_/A vssd1 vssd1 vccd1 vccd1 _2864_/A sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_50_CLK_A clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1734_ _2757_/A vssd1 vssd1 vccd1 vccd1 _1734_/X sky130_fd_sc_hd__buf_2
X_3404_ _3404_/CLK _3404_/D vssd1 vssd1 vccd1 vccd1 _3404_/Q sky130_fd_sc_hd__dfxtp_1
X_1665_ _1644_/X _3232_/Q _1656_/X vssd1 vssd1 vccd1 vccd1 _1665_/X sky130_fd_sc_hd__o21ba_1
X_1596_ _3210_/Q _1576_/X _1595_/Y vssd1 vssd1 vccd1 vccd1 _1596_/X sky130_fd_sc_hd__o21a_1
X_3335_ _3337_/CLK _3335_/D vssd1 vssd1 vccd1 vccd1 _3335_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3266_ _3337_/CLK _3266_/D vssd1 vssd1 vccd1 vccd1 _3266_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1721__A2 _2755_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2217_ _1840_/C _2195_/X _2216_/Y vssd1 vssd1 vccd1 vccd1 _2217_/Y sky130_fd_sc_hd__o21ai_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3197_ _3197_/CLK _3197_/D vssd1 vssd1 vccd1 vccd1 _3197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2148_ _3355_/Q _2145_/X _2147_/Y vssd1 vssd1 vccd1 vccd1 _2148_/X sky130_fd_sc_hd__o21a_1
XFILLER_26_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2079_ _2967_/A vssd1 vssd1 vccd1 vccd1 _2109_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2985__A1 _1815_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3486_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_18_CLK_A clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input145_A core_imem_request_put[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2189__C1 _2152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput309 _2600_/Y vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[30] sky130_fd_sc_hd__buf_2
XANTENNA_output364_A _1881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1450_ _2675_/A vssd1 vssd1 vccd1 vccd1 _1480_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__3153__A1 _2462_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3120_ _3116_/A _2156_/X _2253_/A _3460_/Q _3114_/X vssd1 vssd1 vccd1 vccd1 _3460_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1703__A2 _2751_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3051_ _3093_/A vssd1 vssd1 vccd1 vccd1 _3051_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2002_ _2056_/A vssd1 vssd1 vccd1 vccd1 _2002_/X sky130_fd_sc_hd__buf_2
XANTENNA__1920__C _1920_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2904_ _3322_/Q _2888_/X _2903_/X _2029_/Y vssd1 vssd1 vccd1 vccd1 _3322_/D sky130_fd_sc_hd__o211a_1
X_2835_ _2893_/A vssd1 vssd1 vccd1 vccd1 _2835_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2719__A1 _1516_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2766_ _2757_/X _2766_/A2 _1751_/X _1752_/X _2758_/X vssd1 vssd1 vccd1 vccd1 _3252_/D
+ sky130_fd_sc_hd__a221o_1
X_2697_ _3202_/Q _2695_/X _1572_/Y _2696_/X vssd1 vssd1 vccd1 vccd1 _3202_/D sky130_fd_sc_hd__o211a_1
X_1717_ _1712_/X _1717_/A2 _1715_/X _1716_/X vssd1 vssd1 vccd1 vccd1 _2754_/B sky130_fd_sc_hd__a22oi_4
XFILLER_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1648_ _1776_/B vssd1 vssd1 vccd1 vccd1 _1735_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3318_ _3431_/CLK _3318_/D vssd1 vssd1 vccd1 vccd1 _3318_/Q sky130_fd_sc_hd__dfxtp_1
X_1579_ _1607_/A vssd1 vssd1 vccd1 vccd1 _1579_/X sky130_fd_sc_hd__buf_4
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2495__A _2495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3249_ _3297_/CLK _3249_/D vssd1 vssd1 vccd1 vccd1 _3249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input262_A ram_imem_response_put[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2110__A2 _2093_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output481_A _1461_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2620_ input7/X _2682_/B vssd1 vssd1 vccd1 vccd1 _2677_/B sky130_fd_sc_hd__nor2b_4
X_2551_ _2542_/X _3480_/Q _2543_/X vssd1 vssd1 vccd1 vccd1 _2551_/X sky130_fd_sc_hd__o21ba_1
X_2482_ _2482_/A _2466_/X vssd1 vssd1 vccd1 vccd1 _2482_/X sky130_fd_sc_hd__or2b_1
X_1502_ _1502_/A vssd1 vssd1 vccd1 vccd1 _1503_/C sky130_fd_sc_hd__inv_2
XFILLER_87_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1433_ _3163_/Q _1415_/X _1432_/Y vssd1 vssd1 vccd1 vccd1 _1433_/X sky130_fd_sc_hd__o21a_2
XFILLER_68_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3103_ _3103_/A vssd1 vssd1 vccd1 vccd1 _3103_/X sky130_fd_sc_hd__clkbuf_2
X_3034_ _3399_/Q _3023_/X _2292_/Y _3033_/X vssd1 vssd1 vccd1 vccd1 _3399_/D sky130_fd_sc_hd__o211a_1
XFILLER_55_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2818_ _2818_/A _2818_/B vssd1 vssd1 vccd1 vccd1 _3277_/D sky130_fd_sc_hd__nand2_1
XFILLER_11_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2749_ _2744_/X _2749_/A2 _1693_/X _1694_/X _2745_/X vssd1 vssd1 vccd1 vccd1 _3238_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2876__B1 _2864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3114__A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input108_A core_dmem_request_put[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1569__A _2675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1603__A1 _1496_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput19 core_dmem_request_put[14] vssd1 vssd1 vccd1 vccd1 _1849_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input73_A core_dmem_request_put[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_2_0_CLK_A clkbuf_2_3_0_CLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1470__C _1470_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1982_ _3309_/Q _1965_/X _1981_/Y vssd1 vssd1 vccd1 vccd1 _1982_/X sky130_fd_sc_hd__o21a_2
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2603_ _2603_/A _2464_/X vssd1 vssd1 vccd1 vccd1 _2603_/X sky130_fd_sc_hd__or2b_1
X_2534_ _2542_/A vssd1 vssd1 vccd1 vccd1 _2534_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2465_ _2464_/X _3462_/Q _2470_/A vssd1 vssd1 vccd1 vccd1 _2465_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__2570__A2 _2570_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2396_ _3435_/Q _2383_/X _2395_/Y vssd1 vssd1 vccd1 vccd1 _2396_/X sky130_fd_sc_hd__o21a_1
X_1416_ input3/X vssd1 vssd1 vccd1 vccd1 _1486_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3017_ _1901_/C _3005_/X _3010_/X _2260_/Y vssd1 vssd1 vccd1 vccd1 _3388_/D sky130_fd_sc_hd__o211ai_1
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2013__A _2049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput470 _1528_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[28] sky130_fd_sc_hd__buf_2
XANTENNA__2561__A2 _2561_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput492 _2238_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[19] sky130_fd_sc_hd__buf_2
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput481 _1461_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[9] sky130_fd_sc_hd__buf_2
XFILLER_86_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input225_A ram_dmem_response_put[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1588__B1 _1476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output444_A _2148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2250_ _1885_/C _2224_/X _2249_/Y vssd1 vssd1 vccd1 vccd1 _2250_/Y sky130_fd_sc_hd__o21ai_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1762__A _1762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2181_ _2176_/X _2178_/X _2180_/X _1794_/C _2152_/A vssd1 vssd1 vccd1 vccd1 _2181_/Y
+ sky130_fd_sc_hd__o311ai_4
XFILLER_65_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1965_ _1965_/A vssd1 vssd1 vccd1 vccd1 _1965_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2791__A2 _2779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1896_ _2006_/A vssd1 vssd1 vccd1 vccd1 _1927_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2517_ _2517_/A _2490_/X vssd1 vssd1 vccd1 vccd1 _2517_/X sky130_fd_sc_hd__or2b_1
X_2448_ _2156_/A _2159_/A _2162_/A _2143_/C _2434_/X vssd1 vssd1 vccd1 vccd1 _2448_/Y
+ sky130_fd_sc_hd__o311ai_4
Xinput209 fmc_imem_response_put[9] vssd1 vssd1 vccd1 vccd1 _2746_/A2 sky130_fd_sc_hd__clkbuf_4
X_2379_ _3429_/Q _2355_/X _2378_/Y vssd1 vssd1 vccd1 vccd1 _2379_/X sky130_fd_sc_hd__o21a_1
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2231__A1 _1862_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input175_A fmc_dmem_response_put[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input36_A core_dmem_request_put[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1750_ _2765_/B vssd1 vssd1 vccd1 vccd1 _1750_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output561_A _2418_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1681_ _1669_/X _1681_/A2 _1679_/X _1680_/X vssd1 vssd1 vccd1 vccd1 _2743_/B sky130_fd_sc_hd__a22oi_4
X_3420_ _3420_/CLK _3420_/D vssd1 vssd1 vccd1 vccd1 _3420_/Q sky130_fd_sc_hd__dfxtp_1
X_3351_ _3452_/CLK _3351_/D vssd1 vssd1 vccd1 vccd1 _3351_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2588__A _2588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2302_ _3401_/Q _2297_/X _2301_/Y vssd1 vssd1 vccd1 vccd1 _2302_/X sky130_fd_sc_hd__o21a_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _3288_/CLK _3282_/D vssd1 vssd1 vccd1 vccd1 _3282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2233_ _2211_/X _2212_/X _2213_/X _1866_/C _2232_/X vssd1 vssd1 vccd1 vccd1 _2233_/Y
+ sky130_fd_sc_hd__o311ai_4
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2164_ _2427_/A vssd1 vssd1 vccd1 vccd1 _2225_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_38_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2095_ _2109_/A _2117_/B _2095_/C vssd1 vssd1 vccd1 vccd1 _2095_/Y sky130_fd_sc_hd__nand3_1
XFILLER_65_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2997_ _3373_/Q _2993_/X _2218_/Y _2989_/X vssd1 vssd1 vccd1 vccd1 _3373_/D sky130_fd_sc_hd__o211a_1
X_1948_ _1948_/A vssd1 vssd1 vccd1 vccd1 _1949_/C sky130_fd_sc_hd__clkinv_4
XFILLER_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1879_ _1879_/A vssd1 vssd1 vccd1 vccd1 _1880_/C sky130_fd_sc_hd__inv_4
XANTENNA__2764__A2 _2764_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3122__A _3126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2452__A1 _2225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2755__A2 _2755_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2507__A2 _3132_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output407_A _2027_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2691__A1 _1443_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2920_ _3331_/Q _2912_/X _2062_/Y vssd1 vssd1 vccd1 vccd1 _2921_/A sky130_fd_sc_hd__o21ai_1
XFILLER_31_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2851_ _3295_/Q _2835_/X _1931_/Y vssd1 vssd1 vccd1 vccd1 _2852_/A sky130_fd_sc_hd__o21ai_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2782_ _2782_/A _2797_/B vssd1 vssd1 vccd1 vccd1 _3261_/D sky130_fd_sc_hd__nand2_1
X_1802_ _3261_/Q _1784_/X _1801_/Y vssd1 vssd1 vccd1 vccd1 _1802_/X sky130_fd_sc_hd__o21a_1
X_1733_ _2761_/B vssd1 vssd1 vccd1 vccd1 _1733_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2746__A2 _2746_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3403_ _3459_/CLK _3403_/D vssd1 vssd1 vccd1 vccd1 _3403_/Q sky130_fd_sc_hd__dfxtp_1
X_1664_ _2739_/B vssd1 vssd1 vccd1 vccd1 _1664_/Y sky130_fd_sc_hd__inv_2
X_1595_ _1577_/X _1578_/X _1579_/X _1484_/C _1594_/X vssd1 vssd1 vccd1 vccd1 _1595_/Y
+ sky130_fd_sc_hd__o311ai_4
X_3334_ _3454_/CLK _3334_/D vssd1 vssd1 vccd1 vccd1 _3334_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3265_ _3360_/CLK _3265_/D vssd1 vssd1 vccd1 vccd1 _3265_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ _2196_/X _2206_/X _3372_/Q vssd1 vssd1 vccd1 vccd1 _2216_/Y sky130_fd_sc_hd__o21ai_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ _3226_/CLK _3196_/D vssd1 vssd1 vccd1 vccd1 _3196_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2765__B _2765_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2147_ _2169_/A _2967_/B _2147_/C vssd1 vssd1 vccd1 vccd1 _2147_/Y sky130_fd_sc_hd__nand3_1
XFILLER_53_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2078_ _3335_/Q _2075_/X _2077_/Y vssd1 vssd1 vccd1 vccd1 _2078_/X sky130_fd_sc_hd__o21a_2
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2781__A _2936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2985__A2 _2451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2021__A _2021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2675__B _2675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input138_A core_imem_request_put[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1748__B_N _1644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2189__B1 _1804_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3153__A2 _3153_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1473__C _1473_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3050_ _1981_/C _3049_/X _3039_/X _2324_/Y vssd1 vssd1 vccd1 vccd1 _3410_/D sky130_fd_sc_hd__o211ai_1
X_2001_ _3314_/Q _1984_/X _2000_/Y vssd1 vssd1 vccd1 vccd1 _2001_/X sky130_fd_sc_hd__o21a_1
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2903_ _2969_/B vssd1 vssd1 vccd1 vccd1 _2903_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2834_ _3286_/Q _2830_/X _2826_/X _1898_/Y vssd1 vssd1 vccd1 vccd1 _3286_/D sky130_fd_sc_hd__o211a_1
X_2765_ _2769_/A _2765_/B vssd1 vssd1 vccd1 vccd1 _3251_/D sky130_fd_sc_hd__nor2_1
X_2696_ _2712_/A vssd1 vssd1 vccd1 vccd1 _2696_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1716_ _1716_/A _1705_/X vssd1 vssd1 vccd1 vccd1 _1716_/X sky130_fd_sc_hd__or2b_1
X_1647_ _1644_/X _3228_/Q _2757_/A vssd1 vssd1 vccd1 vccd1 _1647_/X sky130_fd_sc_hd__o21ba_1
X_1578_ _1606_/A vssd1 vssd1 vccd1 vccd1 _1578_/X sky130_fd_sc_hd__buf_4
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2776__A _2959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3317_ _3432_/CLK _3317_/D vssd1 vssd1 vccd1 vccd1 _3317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1680__A _1680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _3252_/CLK _3248_/D vssd1 vssd1 vccd1 vccd1 _3248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3179_ _3244_/CLK _3179_/D vssd1 vssd1 vccd1 vccd1 _3179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input255_A ram_imem_response_put[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output474_A _1540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2550_ _2520_/X _3145_/A2 _2548_/X _2549_/X vssd1 vssd1 vccd1 vccd1 _2550_/X sky130_fd_sc_hd__a22o_1
X_2481_ _2464_/X _3464_/Q _2470_/A vssd1 vssd1 vccd1 vccd1 _2481_/X sky130_fd_sc_hd__o21ba_1
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1501_ _3181_/Q _1498_/X _1500_/Y vssd1 vssd1 vccd1 vccd1 _1501_/X sky130_fd_sc_hd__o21a_2
X_1432_ _2725_/A _1447_/B _1432_/C vssd1 vssd1 vccd1 vccd1 _1432_/Y sky130_fd_sc_hd__nand3_1
XANTENNA_clkbuf_leaf_17_CLK_A clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1931__C _1931_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3102_ _2120_/C _3091_/X _3095_/X _2432_/Y vssd1 vssd1 vccd1 vccd1 _3448_/D sky130_fd_sc_hd__o211ai_1
XFILLER_95_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3033_ _3075_/A vssd1 vssd1 vccd1 vccd1 _3033_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2817_ _3277_/Q _2816_/X _1862_/Y vssd1 vssd1 vccd1 vccd1 _2818_/A sky130_fd_sc_hd__o21ai_1
X_2748_ _2756_/A _2748_/B vssd1 vssd1 vccd1 vccd1 _3237_/D sky130_fd_sc_hd__nor2_1
XFILLER_11_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2679_ _2677_/A _3192_/Q _2658_/A vssd1 vssd1 vccd1 vccd1 _3192_/D sky130_fd_sc_hd__a21bo_1
XFILLER_59_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3130__A _3130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input66_A core_dmem_request_put[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3108__A2 _3105_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3044__A1 _1967_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1981_ _1981_/A _1990_/B _1981_/C vssd1 vssd1 vccd1 vccd1 _1981_/Y sky130_fd_sc_hd__nand3_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2602_ _2478_/X _3159_/Q _2572_/X vssd1 vssd1 vccd1 vccd1 _2602_/X sky130_fd_sc_hd__o21ba_1
X_2533_ _2499_/X _3476_/Q _2500_/X vssd1 vssd1 vccd1 vccd1 _2533_/X sky130_fd_sc_hd__o21ba_1
X_2464_ _2542_/A vssd1 vssd1 vccd1 vccd1 _2464_/X sky130_fd_sc_hd__clkbuf_4
X_2395_ _2384_/X _2385_/X _2386_/X _2072_/C _2377_/X vssd1 vssd1 vccd1 vccd1 _2395_/Y
+ sky130_fd_sc_hd__o311ai_4
X_1415_ _1415_/A vssd1 vssd1 vccd1 vccd1 _1415_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3016_ _3387_/Q _3007_/X _2258_/Y _3003_/X vssd1 vssd1 vccd1 vccd1 _3387_/D sky130_fd_sc_hd__o211a_1
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1836__C _1836_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput471 _1538_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[29] sky130_fd_sc_hd__buf_2
Xoutput460 _1497_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[19] sky130_fd_sc_hd__buf_2
Xoutput493 _2188_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[1] sky130_fd_sc_hd__buf_2
Xoutput482 _2182_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[0] sky130_fd_sc_hd__buf_2
XFILLER_59_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input218_A ram_dmem_response_put[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input120_A core_imem_request_put[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3026__A1 _1917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output437_A _2128_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1760__A1 _1734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2180_ _2300_/A vssd1 vssd1 vccd1 vccd1 _2180_/X sky130_fd_sc_hd__buf_2
XANTENNA__3035__A _3035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3017__A1 _1901_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1964_ _3304_/Q _1947_/X _1963_/Y vssd1 vssd1 vccd1 vccd1 _1964_/X sky130_fd_sc_hd__o21a_2
X_1895_ _3285_/Q _1892_/X _1894_/Y vssd1 vssd1 vccd1 vccd1 _1895_/X sky130_fd_sc_hd__o21a_2
X_2516_ _2499_/X _3472_/Q _2500_/X vssd1 vssd1 vccd1 vccd1 _2516_/X sky130_fd_sc_hd__o21ba_1
X_2447_ _2140_/C _2426_/X _2446_/Y vssd1 vssd1 vccd1 vccd1 _2447_/Y sky130_fd_sc_hd__o21ai_2
X_2378_ _2356_/X _2357_/X _2358_/X _2051_/C _2377_/X vssd1 vssd1 vccd1 vccd1 _2378_/Y
+ sky130_fd_sc_hd__o311ai_2
XANTENNA__2784__A _2864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2059__A2 _2056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2959__A _2959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input168_A fmc_dmem_response_put[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput290 _2532_/X vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[13] sky130_fd_sc_hd__buf_2
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input29_A core_dmem_request_put[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output387_A _1961_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1476__C _1476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1680_ _1680_/A _1661_/X vssd1 vssd1 vccd1 vccd1 _1680_/X sky130_fd_sc_hd__or2b_1
XANTENNA_output554_A _2400_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3350_ _3454_/CLK _3350_/D vssd1 vssd1 vccd1 vccd1 _3350_/Q sky130_fd_sc_hd__dfxtp_1
X_2301_ _2298_/X _2299_/X _2300_/X _1949_/C _2291_/X vssd1 vssd1 vccd1 vccd1 _2301_/Y
+ sky130_fd_sc_hd__o311ai_2
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _3288_/CLK _3281_/D vssd1 vssd1 vccd1 vccd1 _3281_/Q sky130_fd_sc_hd__dfxtp_1
X_2232_ _2291_/A vssd1 vssd1 vccd1 vccd1 _2232_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_78_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2163_ _2163_/A vssd1 vssd1 vccd1 vccd1 _2427_/A sky130_fd_sc_hd__inv_2
XFILLER_38_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2094_ _2094_/A vssd1 vssd1 vccd1 vccd1 _2095_/C sky130_fd_sc_hd__inv_2
XFILLER_0_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2996_ _1840_/C _2991_/X _2995_/X _2216_/Y vssd1 vssd1 vccd1 vccd1 _3372_/D sky130_fd_sc_hd__o211ai_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1947_ _1965_/A vssd1 vssd1 vccd1 vccd1 _1947_/X sky130_fd_sc_hd__clkbuf_2
X_1878_ _3281_/Q _1871_/X _1877_/Y vssd1 vssd1 vccd1 vccd1 _1878_/X sky130_fd_sc_hd__o21a_2
XANTENNA__2779__A _2950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3479_ _3485_/CLK _3479_/D vssd1 vssd1 vccd1 vccd1 _3479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2452__A2 _1801_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2443__A2 _2426_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2850_ _3294_/Q _2849_/X _2845_/X _1927_/Y vssd1 vssd1 vccd1 vccd1 _3294_/D sky130_fd_sc_hd__o211a_1
XFILLER_31_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1801_ _1832_/A _1801_/B _1801_/C vssd1 vssd1 vccd1 vccd1 _1801_/Y sky130_fd_sc_hd__nand3_1
X_2781_ _2936_/A vssd1 vssd1 vccd1 vccd1 _2797_/B sky130_fd_sc_hd__clkbuf_2
X_1732_ _1712_/X _1732_/A2 _1730_/X _1731_/X vssd1 vssd1 vccd1 vccd1 _2761_/B sky130_fd_sc_hd__a22oi_4
XFILLER_7_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1663_ _1633_/X _1663_/A2 _1660_/X _1662_/X vssd1 vssd1 vccd1 vccd1 _2739_/B sky130_fd_sc_hd__a22oi_2
X_3402_ _3404_/CLK _3402_/D vssd1 vssd1 vccd1 vccd1 _3402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1594_ _2675_/A vssd1 vssd1 vccd1 vccd1 _1594_/X sky130_fd_sc_hd__buf_4
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _3337_/CLK _3333_/D vssd1 vssd1 vccd1 vccd1 _3333_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3264_ _3271_/CLK _3264_/D vssd1 vssd1 vccd1 vccd1 _3264_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2215_ _3371_/Q _2210_/X _2214_/Y vssd1 vssd1 vccd1 vccd1 _2215_/X sky130_fd_sc_hd__o21a_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _3226_/CLK _3195_/D vssd1 vssd1 vccd1 vccd1 _3195_/Q sky130_fd_sc_hd__dfxtp_1
X_2146_ _2146_/A vssd1 vssd1 vccd1 vccd1 _2147_/C sky130_fd_sc_hd__clkinv_2
XFILLER_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2077_ _2091_/A _2099_/B _2077_/C vssd1 vssd1 vccd1 vccd1 _2077_/Y sky130_fd_sc_hd__nand3_1
XFILLER_26_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2979_ _3361_/Q _2974_/X _2181_/Y _2978_/X vssd1 vssd1 vccd1 vccd1 _3361_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2198__A1 _1815_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1413__D_N input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input200_A fmc_imem_response_put[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input96_A core_dmem_request_put[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output517_A _2304_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2000_ _2000_/A _2008_/B _2000_/C vssd1 vssd1 vccd1 vccd1 _2000_/Y sky130_fd_sc_hd__nand3_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2902_ _2902_/A _2914_/B vssd1 vssd1 vccd1 vccd1 _3321_/D sky130_fd_sc_hd__nand2_1
X_2833_ _2833_/A _2837_/B vssd1 vssd1 vccd1 vccd1 _3285_/D sky130_fd_sc_hd__nand2_1
XFILLER_31_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2764_ _2757_/X _2764_/A2 _1744_/X _1745_/X _2758_/X vssd1 vssd1 vccd1 vccd1 _3250_/D
+ sky130_fd_sc_hd__a221o_1
X_1715_ _1713_/X _3243_/Q _1714_/X vssd1 vssd1 vccd1 vccd1 _1715_/X sky130_fd_sc_hd__o21ba_1
X_2695_ _2709_/A vssd1 vssd1 vccd1 vccd1 _2695_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2122__A _2206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1646_ _1743_/A vssd1 vssd1 vccd1 vccd1 _2757_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1577_ _1605_/A vssd1 vssd1 vccd1 vccd1 _1577_/X sky130_fd_sc_hd__buf_4
X_3316_ _3431_/CLK _3316_/D vssd1 vssd1 vccd1 vccd1 _3316_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ _3247_/CLK _3247_/D vssd1 vssd1 vccd1 vccd1 _3247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3178_ _3241_/CLK _3178_/D vssd1 vssd1 vccd1 vccd1 _3178_/Q sky130_fd_sc_hd__dfxtp_1
X_2129_ _2145_/A vssd1 vssd1 vccd1 vccd1 _2129_/X sky130_fd_sc_hd__clkbuf_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2343__A1 _2004_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input150_A fmc_dmem_response_put[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input248_A ram_imem_response_put[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input11_A EN_ram_imem_request_get vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2803__C1 _1836_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output467_A _1517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2480_ _2471_/X _3123_/A2 _2476_/X _2479_/X vssd1 vssd1 vccd1 vccd1 _2480_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1484__C _1484_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1500_ _1512_/A _1520_/B _1500_/C vssd1 vssd1 vccd1 vccd1 _1500_/Y sky130_fd_sc_hd__nand3_1
X_1431_ _1431_/A vssd1 vssd1 vccd1 vccd1 _1432_/C sky130_fd_sc_hd__inv_2
XANTENNA__1781__A _2175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3101_ _3447_/Q _3093_/X _2430_/Y _3089_/X vssd1 vssd1 vccd1 vccd1 _3447_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2885__A2 _2868_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3032_ _1938_/C _3021_/X _3025_/X _2289_/Y vssd1 vssd1 vccd1 vccd1 _3398_/D sky130_fd_sc_hd__o211ai_1
XFILLER_36_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput190 fmc_imem_response_put[20] vssd1 vssd1 vccd1 vccd1 _1732_/A2 sky130_fd_sc_hd__buf_2
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2816_ _2893_/A vssd1 vssd1 vccd1 vccd1 _2816_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2168__A4 _2165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2747_ _2747_/A vssd1 vssd1 vccd1 vccd1 _2756_/A sky130_fd_sc_hd__clkbuf_2
X_2678_ _2678_/A vssd1 vssd1 vccd1 vccd1 _3191_/D sky130_fd_sc_hd__clkbuf_1
X_1629_ _1541_/X _1530_/X _1553_/X _3225_/Q vssd1 vssd1 vccd1 vccd1 _1629_/X sky130_fd_sc_hd__a22o_2
XANTENNA__2325__A1 _1981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1691__A _1691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2876__A2 _2868_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input3_A EN_core_imem_request_put vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input198_A fmc_imem_response_put[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input59_A core_dmem_request_put[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1980_ _1980_/A vssd1 vssd1 vccd1 vccd1 _1981_/C sky130_fd_sc_hd__inv_2
XFILLER_26_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2601_ _3140_/A vssd1 vssd1 vccd1 vccd1 _2601_/X sky130_fd_sc_hd__buf_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2532_ _2520_/X _3138_/A2 _2530_/X _2531_/X vssd1 vssd1 vccd1 vccd1 _2532_/X sky130_fd_sc_hd__a22o_1
X_2463_ _2605_/B vssd1 vssd1 vccd1 vccd1 _2542_/A sky130_fd_sc_hd__buf_2
XFILLER_68_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1414_ _2618_/A vssd1 vssd1 vccd1 vccd1 _1415_/A sky130_fd_sc_hd__buf_2
X_2394_ _2069_/C _2369_/X _2393_/Y vssd1 vssd1 vccd1 vccd1 _2394_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__1942__C _1942_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3015_ _1894_/C _3005_/X _3010_/X _2256_/Y vssd1 vssd1 vccd1 vccd1 _3386_/D sky130_fd_sc_hd__o211ai_1
XFILLER_64_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1773__B1_N _1743_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2243__B1 _1873_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput461 _1430_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[1] sky130_fd_sc_hd__buf_2
Xoutput450 _1424_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[0] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_20_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3449_/CLK sky130_fd_sc_hd__clkbuf_16
Xoutput483 _2215_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[10] sky130_fd_sc_hd__buf_2
Xoutput494 _2244_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[20] sky130_fd_sc_hd__buf_2
Xoutput472 _1433_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[2] sky130_fd_sc_hd__buf_2
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1521__A2 _1514_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input113_A core_dmem_request_put[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2980__A _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_16_CLK_A clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_11_CLK clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3222_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1760__A2 _2768_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1963_ _1963_/A _1971_/B _1963_/C vssd1 vssd1 vccd1 vccd1 _1963_/Y sky130_fd_sc_hd__nand3_1
X_1894_ _1909_/A _1917_/B _1894_/C vssd1 vssd1 vccd1 vccd1 _1894_/Y sky130_fd_sc_hd__nand3_1
X_2515_ _2471_/X _3134_/A2 _2512_/X _2514_/X vssd1 vssd1 vccd1 vccd1 _2515_/X sky130_fd_sc_hd__a22o_1
XANTENNA__2130__A _2130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2446_ _2427_/X _1801_/B _3454_/Q vssd1 vssd1 vccd1 vccd1 _2446_/Y sky130_fd_sc_hd__o21ai_1
X_2377_ _2434_/A vssd1 vssd1 vccd1 vccd1 _2377_/X sky130_fd_sc_hd__buf_2
XFILLER_68_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1847__C _1847_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput280 _1542_/X vssd1 vssd1 vccd1 vccd1 RDY_fmc_imem_request_get sky130_fd_sc_hd__buf_2
Xoutput291 _2537_/Y vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[14] sky130_fd_sc_hd__buf_2
XANTENNA_input230_A ram_dmem_response_put[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3241_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output547_A _2382_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2300_ _2300_/A vssd1 vssd1 vccd1 vccd1 _2300_/X sky130_fd_sc_hd__buf_2
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3280_ _3360_/CLK _3280_/D vssd1 vssd1 vccd1 vccd1 _3280_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1492__C _1492_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2231_ _1862_/C _2224_/X _2230_/Y vssd1 vssd1 vccd1 vccd1 _2231_/Y sky130_fd_sc_hd__o21ai_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2162_ _2162_/A vssd1 vssd1 vccd1 vccd1 _2162_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2694__B1 _2686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2093_ _2145_/A vssd1 vssd1 vccd1 vccd1 _2093_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2995_ _3103_/A vssd1 vssd1 vccd1 vccd1 _2995_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1946_ _3299_/Q _1929_/X _1945_/Y vssd1 vssd1 vccd1 vccd1 _1946_/X sky130_fd_sc_hd__o21a_2
X_1877_ _1909_/A _1877_/B _1877_/C vssd1 vssd1 vccd1 vccd1 _1877_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__1724__A2 _1724_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3478_ _3482_/CLK _3478_/D vssd1 vssd1 vccd1 vccd1 _3478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2429_ _2113_/C _2426_/X _2428_/Y vssd1 vssd1 vccd1 vccd1 _2429_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__2795__A _2945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2035__A _2035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input180_A fmc_imem_response_put[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input41_A core_dmem_request_put[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1800_ _1800_/A vssd1 vssd1 vccd1 vccd1 _1801_/C sky130_fd_sc_hd__inv_6
XFILLER_31_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2780_ _3261_/Q _2779_/X _1801_/Y vssd1 vssd1 vccd1 vccd1 _2782_/A sky130_fd_sc_hd__o21ai_1
X_1731_ _1731_/A _1705_/X vssd1 vssd1 vccd1 vccd1 _1731_/X sky130_fd_sc_hd__or2b_1
XFILLER_7_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1662_ _1662_/A _1661_/X vssd1 vssd1 vccd1 vccd1 _1662_/X sky130_fd_sc_hd__or2b_1
X_3401_ _3459_/CLK _3401_/D vssd1 vssd1 vccd1 vccd1 _3401_/Q sky130_fd_sc_hd__dfxtp_1
X_3332_ _3454_/CLK _3332_/D vssd1 vssd1 vccd1 vccd1 _3332_/Q sky130_fd_sc_hd__dfxtp_1
X_1593_ _1480_/C _1590_/X _1592_/Y vssd1 vssd1 vccd1 vccd1 _1593_/Y sky130_fd_sc_hd__o21ai_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _3271_/CLK _3263_/D vssd1 vssd1 vccd1 vccd1 _3263_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _2211_/X _2212_/X _2213_/X _1836_/C _2203_/X vssd1 vssd1 vccd1 vccd1 _2214_/Y
+ sky130_fd_sc_hd__o311ai_2
X_3194_ _3226_/CLK _3194_/D vssd1 vssd1 vccd1 vccd1 _3194_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2145_ _2145_/A vssd1 vssd1 vccd1 vccd1 _2145_/X sky130_fd_sc_hd__buf_4
XFILLER_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2076_ _2076_/A vssd1 vssd1 vccd1 vccd1 _2077_/C sky130_fd_sc_hd__clkinv_2
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2978_ _3103_/A vssd1 vssd1 vccd1 vccd1 _2978_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1929_ _1965_/A vssd1 vssd1 vccd1 vccd1 _1929_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1694__A _1694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input89_A core_dmem_request_put[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1624__A1 _1523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2901_ _3321_/Q _2893_/X _2026_/Y vssd1 vssd1 vccd1 vccd1 _2902_/A sky130_fd_sc_hd__o21ai_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2832_ _3285_/Q _2816_/X _1894_/Y vssd1 vssd1 vccd1 vccd1 _2833_/A sky130_fd_sc_hd__o21ai_1
X_2763_ _2769_/A _2763_/B vssd1 vssd1 vccd1 vccd1 _3249_/D sky130_fd_sc_hd__nor2_1
X_1714_ input8/X vssd1 vssd1 vccd1 vccd1 _1714_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1945__C _1945_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2694_ _1452_/C _2693_/X _2686_/X _1570_/Y vssd1 vssd1 vccd1 vccd1 _3201_/D sky130_fd_sc_hd__o211ai_1
XFILLER_6_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1645_ input8/X vssd1 vssd1 vccd1 vccd1 _1743_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1576_ _1630_/B vssd1 vssd1 vccd1 vccd1 _1576_/X sky130_fd_sc_hd__clkbuf_2
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3315_ _3432_/CLK _3315_/D vssd1 vssd1 vccd1 vccd1 _3315_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__1560__B1 _1438_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ _3252_/CLK _3246_/D vssd1 vssd1 vccd1 vccd1 _3246_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3177_ _3247_/CLK _3177_/D vssd1 vssd1 vccd1 vccd1 _3177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2128_ _3349_/Q _2111_/X _2127_/Y vssd1 vssd1 vccd1 vccd1 _2128_/X sky130_fd_sc_hd__o21a_2
X_2059_ _3330_/Q _2056_/X _2058_/Y vssd1 vssd1 vccd1 vccd1 _2059_/X sky130_fd_sc_hd__o21a_1
XFILLER_54_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1615__A1 _1509_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2967__B _2967_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input143_A core_imem_request_put[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2582__A2 _3153_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output362_A _1874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1430_ _3162_/Q _1415_/X _1429_/Y vssd1 vssd1 vccd1 vccd1 _1430_/X sky130_fd_sc_hd__o21a_2
XANTENNA__1781__B _2177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3100_ _2113_/C _3091_/X _3095_/X _2428_/Y vssd1 vssd1 vccd1 vccd1 _3446_/D sky130_fd_sc_hd__o211ai_1
X_3031_ _3397_/Q _3023_/X _2287_/Y _3019_/X vssd1 vssd1 vccd1 vccd1 _3397_/D sky130_fd_sc_hd__o211a_1
Xinput180 fmc_imem_response_put[11] vssd1 vssd1 vccd1 vccd1 _2749_/A2 sky130_fd_sc_hd__clkbuf_4
XANTENNA__2893__A _2893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput191 fmc_imem_response_put[21] vssd1 vssd1 vccd1 vccd1 _2762_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2815_ _2815_/A vssd1 vssd1 vccd1 vccd1 _2893_/A sky130_fd_sc_hd__buf_2
XANTENNA__2133__A _2133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2746_ _2744_/X _2746_/A2 _1683_/X _1685_/X _2745_/X vssd1 vssd1 vccd1 vccd1 _3236_/D
+ sky130_fd_sc_hd__a221o_1
Xoutput610 _1568_/X vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[6] sky130_fd_sc_hd__buf_2
X_2677_ _2677_/A _2677_/B _3191_/Q vssd1 vssd1 vccd1 vccd1 _2678_/A sky130_fd_sc_hd__and3_1
X_1628_ _1541_/X _2725_/B _1553_/X _3224_/Q vssd1 vssd1 vccd1 vccd1 _1628_/X sky130_fd_sc_hd__a22o_2
X_1559_ _1435_/C _1553_/X _1558_/Y vssd1 vssd1 vccd1 vccd1 _1559_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_86_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3229_ _3466_/CLK _3229_/D vssd1 vssd1 vccd1 vccd1 _3229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2261__A1 _1901_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2043__A _2043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2978__A _3103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input260_A ram_imem_response_put[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1776__B _1776_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3049__A _3091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2600_ _2614_/B vssd1 vssd1 vccd1 vccd1 _2600_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2888__A _2945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2531_ _2531_/A _2513_/X vssd1 vssd1 vccd1 vccd1 _2531_/X sky130_fd_sc_hd__or2b_1
XFILLER_5_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1792__A _2206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2462_ _2470_/A vssd1 vssd1 vccd1 vccd1 _2462_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1413_ _1529_/A _1531_/A _1533_/A input3/X vssd1 vssd1 vccd1 vccd1 _2618_/A sky130_fd_sc_hd__nor4b_1
X_2393_ _2370_/X _2380_/X _3434_/Q vssd1 vssd1 vccd1 vccd1 _2393_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_68_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3014_ _3385_/Q _3007_/X _2251_/Y _3003_/X vssd1 vssd1 vccd1 vccd1 _3385_/D sky130_fd_sc_hd__o211a_1
XFILLER_36_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2729_ _2725_/A _1530_/X _1562_/A _3225_/Q _2723_/X vssd1 vssd1 vccd1 vccd1 _3225_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_3_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2546__A2 _2546_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput440 _2135_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[91] sky130_fd_sc_hd__buf_2
Xoutput451 _1465_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[10] sky130_fd_sc_hd__buf_2
Xoutput462 _1501_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[20] sky130_fd_sc_hd__buf_2
Xoutput484 _2217_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[11] sky130_fd_sc_hd__buf_2
Xoutput495 _2246_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[21] sky130_fd_sc_hd__buf_2
Xoutput473 _1539_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[30] sky130_fd_sc_hd__buf_2
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input106_A core_dmem_request_put[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2785__A2 _2145_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input71_A core_dmem_request_put[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2170__B1 _3360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1787__A _2319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1962_ _1962_/A vssd1 vssd1 vccd1 vccd1 _1963_/C sky130_fd_sc_hd__clkinv_4
X_1893_ _1893_/A vssd1 vssd1 vccd1 vccd1 _1894_/C sky130_fd_sc_hd__clkinv_4
XANTENNA__2411__A _2459_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2514_ _2514_/A _2513_/X vssd1 vssd1 vccd1 vccd1 _2514_/X sky130_fd_sc_hd__or2b_1
XANTENNA__1953__C _1953_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2445_ _3453_/Q _2439_/X _2444_/Y vssd1 vssd1 vccd1 vccd1 _2445_/X sky130_fd_sc_hd__o21a_1
XFILLER_88_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2376_ _2047_/C _2369_/X _2375_/Y vssd1 vssd1 vccd1 vccd1 _2376_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1697__A _1697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput281 _3491_/A vssd1 vssd1 vccd1 vccd1 RDY_fmc_imem_response_put sky130_fd_sc_hd__buf_2
Xoutput292 _2540_/X vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[15] sky130_fd_sc_hd__buf_2
XFILLER_87_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2975__B _2975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input223_A ram_dmem_response_put[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2991__A _3035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output442_A _2141_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _2225_/X _2206_/X _3378_/Q vssd1 vssd1 vccd1 vccd1 _2230_/Y sky130_fd_sc_hd__o21ai_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2161_ _2414_/A vssd1 vssd1 vccd1 vccd1 _2162_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_65_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2694__A1 _1452_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2092_ _3339_/Q _2075_/X _2091_/Y vssd1 vssd1 vccd1 vccd1 _2092_/X sky130_fd_sc_hd__o21a_2
XFILLER_65_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2994_ _3371_/Q _2993_/X _2214_/Y _2989_/X vssd1 vssd1 vccd1 vccd1 _3371_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1945_ _1945_/A _1953_/B _1945_/C vssd1 vssd1 vccd1 vccd1 _1945_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__2749__A2 _2749_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1876_ _1876_/A vssd1 vssd1 vccd1 vccd1 _1877_/C sky130_fd_sc_hd__clkinv_4
XFILLER_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3477_ _3477_/CLK _3477_/D vssd1 vssd1 vccd1 vccd1 _3477_/Q sky130_fd_sc_hd__dfxtp_1
X_2428_ _2427_/X _2408_/X _3446_/Q vssd1 vssd1 vccd1 vccd1 _2428_/Y sky130_fd_sc_hd__o21ai_2
X_2359_ _2356_/X _2357_/X _2358_/X _2022_/C _2348_/X vssd1 vssd1 vccd1 vccd1 _2359_/Y
+ sky130_fd_sc_hd__o311ai_4
XFILLER_69_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_15_CLK_A clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input173_A fmc_dmem_response_put[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input34_A core_dmem_request_put[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1651__A2 _2736_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1730_ _1713_/X _3247_/Q _1714_/X vssd1 vssd1 vccd1 vccd1 _1730_/X sky130_fd_sc_hd__o21ba_1
X_1661_ _1713_/A vssd1 vssd1 vccd1 vccd1 _1661_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3400_ _3404_/CLK _3400_/D vssd1 vssd1 vccd1 vccd1 _3400_/Q sky130_fd_sc_hd__dfxtp_1
X_1592_ _1591_/X _1569_/X _3209_/Q vssd1 vssd1 vccd1 vccd1 _1592_/Y sky130_fd_sc_hd__o21ai_1
X_3331_ _3337_/CLK _3331_/D vssd1 vssd1 vccd1 vccd1 _3331_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3271_/CLK _3262_/D vssd1 vssd1 vccd1 vccd1 _3262_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ _2300_/A vssd1 vssd1 vccd1 vccd1 _2213_/X sky130_fd_sc_hd__clkbuf_4
X_3193_ _3241_/CLK _3193_/D vssd1 vssd1 vccd1 vccd1 _3193_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2144_ _3354_/Q _2129_/X _2143_/Y vssd1 vssd1 vccd1 vccd1 _2144_/X sky130_fd_sc_hd__o21a_1
XFILLER_66_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2075_ _2145_/A vssd1 vssd1 vccd1 vccd1 _2075_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_19_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3092__A1 _2091_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2136__A _2136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2977_ _3095_/A vssd1 vssd1 vccd1 vccd1 _3103_/A sky130_fd_sc_hd__clkbuf_4
X_1928_ _3294_/Q _1911_/X _1927_/Y vssd1 vssd1 vccd1 vccd1 _1928_/X sky130_fd_sc_hd__o21a_2
X_1859_ _1888_/A _1859_/B _1859_/C vssd1 vssd1 vccd1 vccd1 _1859_/Y sky130_fd_sc_hd__nand3_2
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3147__A2 _3147_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3138__A2 _3138_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3074__A1 _2047_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2900_ _3320_/Q _2888_/X _2884_/X _2022_/Y vssd1 vssd1 vccd1 vccd1 _3320_/D sky130_fd_sc_hd__o211a_1
XFILLER_91_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2831_ _3284_/Q _2830_/X _2826_/X _1888_/Y vssd1 vssd1 vccd1 vccd1 _3284_/D sky130_fd_sc_hd__o211a_1
XFILLER_31_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2762_ _2757_/X _2762_/A2 _1736_/X _1737_/X _2758_/X vssd1 vssd1 vccd1 vccd1 _3248_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_8_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1713_ _1713_/A vssd1 vssd1 vccd1 vccd1 _1713_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2693_ _2707_/A vssd1 vssd1 vccd1 vccd1 _2693_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__3129__A2 _3129_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1644_ _1644_/A vssd1 vssd1 vccd1 vccd1 _1644_/X sky130_fd_sc_hd__clkbuf_2
X_1575_ _1460_/C _1562_/X _1574_/Y vssd1 vssd1 vccd1 vccd1 _1575_/Y sky130_fd_sc_hd__o21ai_2
X_3314_ _3460_/CLK _3314_/D vssd1 vssd1 vccd1 vccd1 _3314_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _3247_/CLK _3245_/D vssd1 vssd1 vccd1 vccd1 _3245_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3176_ _3241_/CLK _3176_/D vssd1 vssd1 vccd1 vccd1 _3176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2127_ _2127_/A _2134_/B _2127_/C vssd1 vssd1 vccd1 vccd1 _2127_/Y sky130_fd_sc_hd__nand3_1
X_2058_ _2072_/A _2081_/B _2058_/C vssd1 vssd1 vccd1 vccd1 _2058_/Y sky130_fd_sc_hd__nand3_1
XFILLER_54_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input136_A core_imem_request_put[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__3056__A1 _1997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1781__C _2179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput170 fmc_dmem_response_put[31] vssd1 vssd1 vccd1 vccd1 _2615_/A2 sky130_fd_sc_hd__clkbuf_4
X_3030_ _1931_/C _3021_/X _3025_/X _2285_/Y vssd1 vssd1 vccd1 vccd1 _3396_/D sky130_fd_sc_hd__o211ai_1
XFILLER_48_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput181 fmc_imem_response_put[12] vssd1 vssd1 vccd1 vccd1 _1698_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput192 fmc_imem_response_put[22] vssd1 vssd1 vccd1 vccd1 _1741_/A2 sky130_fd_sc_hd__buf_2
XFILLER_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2814_ _3276_/Q _2810_/X _2806_/X _1859_/Y vssd1 vssd1 vccd1 vccd1 _3276_/D sky130_fd_sc_hd__o211a_1
XFILLER_31_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1956__C _1956_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2745_ _2760_/A vssd1 vssd1 vccd1 vccd1 _2745_/X sky130_fd_sc_hd__clkbuf_2
Xoutput611 _1571_/Y vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[7] sky130_fd_sc_hd__buf_2
Xoutput600 _1622_/X vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[26] sky130_fd_sc_hd__buf_2
X_2676_ _2677_/A _3190_/Q _2658_/A vssd1 vssd1 vccd1 vccd1 _3190_/D sky130_fd_sc_hd__a21bo_1
X_1627_ _1541_/X _1534_/X _1553_/X _3223_/Q vssd1 vssd1 vccd1 vccd1 _1627_/X sky130_fd_sc_hd__a22o_2
XFILLER_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1558_ _1537_/X _1527_/B _3197_/Q vssd1 vssd1 vccd1 vccd1 _1558_/Y sky130_fd_sc_hd__o21ai_1
X_1489_ _3178_/Q _1478_/X _1488_/Y vssd1 vssd1 vccd1 vccd1 _1489_/X sky130_fd_sc_hd__o21a_2
XANTENNA__2089__A2 _2075_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3228_ _3259_/CLK _3228_/D vssd1 vssd1 vccd1 vccd1 _3228_/Q sky130_fd_sc_hd__dfxtp_1
X_3159_ _3489_/CLK _3159_/D vssd1 vssd1 vccd1 vccd1 _3159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1866__C _1866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input253_A ram_imem_response_put[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1776__C input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output472_A _1433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2530_ _2521_/X _3475_/Q _2529_/X vssd1 vssd1 vccd1 vccd1 _2530_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__2960__B1 _2959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2461_ input6/X vssd1 vssd1 vccd1 vccd1 _2470_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1763__A1 _1691_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1412_ _3461_/Q _3360_/Q vssd1 vssd1 vccd1 vccd1 _1412_/Y sky130_fd_sc_hd__nor2_1
X_2392_ _3433_/Q _2383_/X _2391_/Y vssd1 vssd1 vccd1 vccd1 _2392_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3013_ _1885_/C _3005_/X _3010_/X _2249_/Y vssd1 vssd1 vccd1 vccd1 _3384_/D sky130_fd_sc_hd__o211ai_1
XFILLER_36_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1983__A _2794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2728_ _2725_/Y _2727_/Y _2723_/X vssd1 vssd1 vccd1 vccd1 _3224_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__1754__A1 _1637_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput430 _2103_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[82] sky130_fd_sc_hd__buf_2
Xoutput441 _2138_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[92] sky130_fd_sc_hd__buf_2
Xoutput452 _1468_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[11] sky130_fd_sc_hd__buf_2
X_2659_ _2659_/A _2673_/B vssd1 vssd1 vccd1 vccd1 _3180_/D sky130_fd_sc_hd__nand2_1
Xoutput485 _2219_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[12] sky130_fd_sc_hd__buf_2
Xoutput496 _2248_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[22] sky130_fd_sc_hd__buf_2
Xoutput474 _1540_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[31] sky130_fd_sc_hd__buf_2
Xoutput463 _1504_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[21] sky130_fd_sc_hd__buf_2
XFILLER_86_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2319__A _2319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2989__A _3003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input64_A core_dmem_request_put[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2170__A1 _2169_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1961_ _3303_/Q _1947_/X _1960_/Y vssd1 vssd1 vccd1 vccd1 _1961_/X sky130_fd_sc_hd__o21a_2
XFILLER_14_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1892_ _1965_/A vssd1 vssd1 vccd1 vccd1 _1892_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2513_ _2564_/A vssd1 vssd1 vccd1 vccd1 _2513_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2444_ _2156_/A _2159_/A _2162_/A _2137_/C _2434_/X vssd1 vssd1 vccd1 vccd1 _2444_/Y
+ sky130_fd_sc_hd__o311ai_4
X_2375_ _2370_/X _2351_/X _3428_/Q vssd1 vssd1 vccd1 vccd1 _2375_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_68_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2139__A _2139_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3110__B1 _3003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2040__C _2040_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput282 _2460_/X vssd1 vssd1 vccd1 vccd1 RDY_ram_dmem_request_get sky130_fd_sc_hd__buf_2
Xoutput293 _2547_/Y vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[16] sky130_fd_sc_hd__buf_2
XFILLER_87_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2049__A _2049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2455__A2 _2439_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input216_A ram_dmem_response_put[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output435_A _2121_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2160_ _2179_/A vssd1 vssd1 vccd1 vccd1 _2414_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output602_A _1626_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2091_ _2091_/A _2099_/B _2091_/C vssd1 vssd1 vccd1 vccd1 _2091_/Y sky130_fd_sc_hd__nand3_1
XFILLER_93_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2446__A2 _1801_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2993_ _3037_/A vssd1 vssd1 vccd1 vccd1 _2993_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1944_ _1944_/A vssd1 vssd1 vccd1 vccd1 _1945_/C sky130_fd_sc_hd__inv_2
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1875_ _1951_/A vssd1 vssd1 vccd1 vccd1 _1909_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3476_ _3476_/CLK _3476_/D vssd1 vssd1 vccd1 vccd1 _3476_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2382__A1 _2054_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2427_ _2427_/A vssd1 vssd1 vccd1 vccd1 _2427_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2358_ _2414_/A vssd1 vssd1 vccd1 vccd1 _2358_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2289_ _2284_/X _2265_/X _3398_/Q vssd1 vssd1 vccd1 vccd1 _2289_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2437__A2 _1801_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2620__B_N _2682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input166_A fmc_dmem_response_put[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input27_A core_dmem_request_put[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1411__A _3226_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output385_A _1954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1660_ _1635_/X _3231_/Q _1641_/A vssd1 vssd1 vccd1 vccd1 _1660_/X sky130_fd_sc_hd__o21ba_1
XANTENNA_output552_A _2394_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1591_ _1591_/A vssd1 vssd1 vccd1 vccd1 _1591_/X sky130_fd_sc_hd__clkbuf_2
X_3330_ _3330_/CLK _3330_/D vssd1 vssd1 vccd1 vccd1 _3330_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3261_ _3271_/CLK _3261_/D vssd1 vssd1 vccd1 vccd1 _3261_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ _2299_/A vssd1 vssd1 vccd1 vccd1 _2212_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3192_ _3258_/CLK _3192_/D vssd1 vssd1 vccd1 vccd1 _3192_/Q sky130_fd_sc_hd__dfxtp_1
X_2143_ _2143_/A _2152_/B _2143_/C vssd1 vssd1 vccd1 vccd1 _2143_/Y sky130_fd_sc_hd__nand3_1
XFILLER_66_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2074_ _2794_/A vssd1 vssd1 vccd1 vccd1 _2145_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2976_ _3009_/A vssd1 vssd1 vccd1 vccd1 _3095_/A sky130_fd_sc_hd__clkbuf_4
X_1927_ _1927_/A _1935_/B _1927_/C vssd1 vssd1 vccd1 vccd1 _1927_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__2152__A _2152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1858_ _1858_/A vssd1 vssd1 vccd1 vccd1 _1859_/C sky130_fd_sc_hd__inv_4
X_1789_ _1789_/A _1789_/B _1789_/C vssd1 vssd1 vccd1 vccd1 _2235_/A sky130_fd_sc_hd__nor3_2
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3459_ _3459_/CLK _3459_/D vssd1 vssd1 vccd1 vccd1 _3459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1869__C _1869_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2830_ _2868_/A vssd1 vssd1 vccd1 vccd1 _2830_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2761_ _2769_/A _2761_/B vssd1 vssd1 vccd1 vccd1 _3247_/D sky130_fd_sc_hd__nor2_1
XFILLER_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2692_ _3200_/Q _2681_/X _1567_/Y _2684_/X vssd1 vssd1 vccd1 vccd1 _3200_/D sky130_fd_sc_hd__o211a_1
XANTENNA__2585__A1 _2520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1712_ _1712_/A vssd1 vssd1 vccd1 vccd1 _1712_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_14_CLK_A clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1643_ _1776_/B vssd1 vssd1 vccd1 vccd1 _1644_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2337__A1 _1997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1574_ _1563_/X _1569_/X _3203_/Q vssd1 vssd1 vccd1 vccd1 _1574_/Y sky130_fd_sc_hd__o21ai_1
X_3313_ _3420_/CLK _3313_/D vssd1 vssd1 vccd1 vccd1 _3313_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_29_CLK_A clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3244_ _3244_/CLK _3244_/D vssd1 vssd1 vccd1 vccd1 _3244_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3175_ _3247_/CLK _3175_/D vssd1 vssd1 vccd1 vccd1 _3175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2126_ _2126_/A vssd1 vssd1 vccd1 vccd1 _2127_/C sky130_fd_sc_hd__inv_2
XANTENNA__2147__A _2169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2057_ _2057_/A vssd1 vssd1 vccd1 vccd1 _2058_/C sky130_fd_sc_hd__inv_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2959_ _2959_/A vssd1 vssd1 vccd1 vccd1 _2959_/X sky130_fd_sc_hd__buf_2
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2610__A _3130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3259_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input129_A core_imem_request_put[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2057__A _2057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1896__A _2006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input94_A core_dmem_request_put[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2520__A _2520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_41_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3252_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput171 fmc_dmem_response_put[3] vssd1 vssd1 vccd1 vccd1 _3125_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput160 fmc_dmem_response_put[22] vssd1 vssd1 vccd1 vccd1 _2570_/A2 sky130_fd_sc_hd__buf_2
Xinput193 fmc_imem_response_put[23] vssd1 vssd1 vccd1 vccd1 _2764_/A2 sky130_fd_sc_hd__buf_2
XFILLER_48_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput182 fmc_imem_response_put[13] vssd1 vssd1 vccd1 vccd1 _2751_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_63_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2813_ _2813_/A _2818_/B vssd1 vssd1 vccd1 vccd1 _3275_/D sky130_fd_sc_hd__nand2_1
XFILLER_31_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2744_ _2757_/A vssd1 vssd1 vccd1 vccd1 _2744_/X sky130_fd_sc_hd__clkbuf_2
Xoutput601 _1624_/Y vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[27] sky130_fd_sc_hd__buf_2
X_2675_ _2675_/A _2675_/B vssd1 vssd1 vccd1 vccd1 _2677_/A sky130_fd_sc_hd__nand2_1
Xoutput612 _1573_/X vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[8] sky130_fd_sc_hd__buf_2
X_1626_ _3222_/Q _1604_/X _1625_/Y vssd1 vssd1 vccd1 vccd1 _1626_/X sky130_fd_sc_hd__o21a_2
Xclkbuf_leaf_32_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3440_/CLK sky130_fd_sc_hd__clkbuf_16
X_1557_ _3196_/Q _1545_/X _1556_/Y vssd1 vssd1 vccd1 vccd1 _1557_/X sky130_fd_sc_hd__o21a_1
XFILLER_86_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2730__A1 _3226_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1488_ _1516_/A _1488_/B _1488_/C vssd1 vssd1 vccd1 vccd1 _1488_/Y sky130_fd_sc_hd__nand3_1
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3227_ _3472_/CLK _3227_/D vssd1 vssd1 vccd1 vccd1 _3227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3158_ _3489_/CLK _3158_/D vssd1 vssd1 vccd1 vccd1 _3158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2109_ _2109_/A _2117_/B _2109_/C vssd1 vssd1 vccd1 vccd1 _2109_/Y sky130_fd_sc_hd__nand3_1
XFILLER_54_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3089_ _3103_/A vssd1 vssd1 vccd1 vccd1 _3089_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_23_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3330_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2340__A _2397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2721__A1 _1523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1524__A2 _1514_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input246_A ram_imem_response_put[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output465_A _1510_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2460_ _2460_/A vssd1 vssd1 vccd1 vccd1 _2460_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_14_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3394_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__1763__A2 _1763_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1411_ _3226_/Q _3193_/Q vssd1 vssd1 vccd1 vccd1 _1411_/Y sky130_fd_sc_hd__nor2_2
X_2391_ _2384_/X _2385_/X _2386_/X _2065_/C _2377_/X vssd1 vssd1 vccd1 vccd1 _2391_/Y
+ sky130_fd_sc_hd__o311ai_2
XFILLER_3_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3081__A _3095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3012_ _3383_/Q _3007_/X _2247_/Y _3003_/X vssd1 vssd1 vccd1 vccd1 _3383_/D sky130_fd_sc_hd__o211a_1
XFILLER_83_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2228__B1 _1859_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1967__C _1967_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2727_ _1563_/A _1527_/B _2726_/Y vssd1 vssd1 vccd1 vccd1 _2727_/Y sky130_fd_sc_hd__o21bai_1
Xoutput420 _2070_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[73] sky130_fd_sc_hd__buf_2
XANTENNA__2160__A _2179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput442 _2141_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[93] sky130_fd_sc_hd__buf_2
Xoutput431 _2107_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[83] sky130_fd_sc_hd__buf_2
Xoutput453 _1471_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[12] sky130_fd_sc_hd__buf_2
X_2658_ _2658_/A vssd1 vssd1 vccd1 vccd1 _2673_/B sky130_fd_sc_hd__clkbuf_2
Xoutput486 _2221_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[13] sky130_fd_sc_hd__buf_2
X_1609_ _3214_/Q _1604_/X _1608_/Y vssd1 vssd1 vccd1 vccd1 _1609_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2703__A1 _1473_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput475 _1436_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[3] sky130_fd_sc_hd__buf_2
X_2589_ _2563_/X _3155_/A2 _2587_/X _2588_/X vssd1 vssd1 vccd1 vccd1 _2589_/X sky130_fd_sc_hd__a22o_1
Xoutput464 _1507_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[22] sky130_fd_sc_hd__buf_2
Xoutput497 _2250_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[23] sky130_fd_sc_hd__buf_2
XFILLER_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input1_A EN_core_dmem_request_put vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1877__C _1877_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input196_A fmc_imem_response_put[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input57_A core_dmem_request_put[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2458__B1 _2185_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_CLK clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3225_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1960_ _1981_/A _1990_/B _1960_/C vssd1 vssd1 vccd1 vccd1 _1960_/Y sky130_fd_sc_hd__nand3_1
X_1891_ _2794_/A vssd1 vssd1 vccd1 vccd1 _1965_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2512_ _2473_/X _3471_/Q _2485_/X vssd1 vssd1 vccd1 vccd1 _2512_/X sky130_fd_sc_hd__o21ba_1
X_2443_ _2134_/C _2426_/X _2442_/Y vssd1 vssd1 vccd1 vccd1 _2443_/Y sky130_fd_sc_hd__o21ai_2
X_2374_ _3427_/Q _2355_/X _2373_/Y vssd1 vssd1 vccd1 vccd1 _2374_/X sky130_fd_sc_hd__o21a_1
XFILLER_68_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput283 _3490_/X vssd1 vssd1 vccd1 vccd1 RDY_ram_dmem_response_put sky130_fd_sc_hd__buf_2
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput294 _2550_/X vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[17] sky130_fd_sc_hd__buf_2
XFILLER_59_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input111_A core_dmem_request_put[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input209_A fmc_imem_response_put[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2090_ _2090_/A vssd1 vssd1 vccd1 vccd1 _2091_/C sky130_fd_sc_hd__clkinv_2
XFILLER_19_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2992_ _1832_/C _2991_/X _2980_/X _2207_/Y vssd1 vssd1 vccd1 vccd1 _3370_/D sky130_fd_sc_hd__o211ai_1
XFILLER_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1943_ _3298_/Q _1929_/X _1942_/Y vssd1 vssd1 vccd1 vccd1 _1943_/X sky130_fd_sc_hd__o21a_2
X_1874_ _3280_/Q _1871_/X _1873_/Y vssd1 vssd1 vccd1 vccd1 _1874_/X sky130_fd_sc_hd__o21a_1
X_3475_ _3477_/CLK _3475_/D vssd1 vssd1 vccd1 vccd1 _3475_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2426_ _3035_/A vssd1 vssd1 vccd1 vccd1 _2426_/X sky130_fd_sc_hd__buf_4
XFILLER_84_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2357_ _2413_/A vssd1 vssd1 vccd1 vccd1 _2357_/X sky130_fd_sc_hd__clkbuf_4
X_2288_ _3397_/Q _2268_/X _2287_/Y vssd1 vssd1 vccd1 vccd1 _2288_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2125__A2 _2111_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input159_A fmc_dmem_response_put[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2595__B_N _2464_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2523__A _2523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output378_A _1932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output280_A _1542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1590_ _2707_/A vssd1 vssd1 vccd1 vccd1 _1590_/X sky130_fd_sc_hd__buf_2
XANTENNA__1572__B1 _1456_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _3271_/CLK _3260_/D vssd1 vssd1 vccd1 vccd1 _3260_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2211_ _2298_/A vssd1 vssd1 vccd1 vccd1 _2211_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ _3197_/CLK _3191_/D vssd1 vssd1 vccd1 vccd1 _3191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2142_ _2142_/A vssd1 vssd1 vccd1 vccd1 _2143_/C sky130_fd_sc_hd__clkinv_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2073_ _3334_/Q _2056_/X _2072_/Y vssd1 vssd1 vccd1 vccd1 _2073_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2975_ input9/X _2975_/B vssd1 vssd1 vccd1 vccd1 _3009_/A sky130_fd_sc_hd__and2b_1
X_1926_ _1926_/A vssd1 vssd1 vccd1 vccd1 _1927_/C sky130_fd_sc_hd__clkinv_4
X_1857_ _2006_/A vssd1 vssd1 vccd1 vccd1 _1888_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1788_ _2967_/A vssd1 vssd1 vccd1 vccd1 _3116_/A sky130_fd_sc_hd__buf_4
XFILLER_89_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3458_ _3460_/CLK _3458_/D vssd1 vssd1 vccd1 vccd1 _3458_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2107__A2 _2093_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3389_ _3397_/CLK _3389_/D vssd1 vssd1 vccd1 vccd1 _3389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2409_ _2398_/X _2408_/X _3440_/Q vssd1 vssd1 vccd1 vccd1 _2409_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_84_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1885__C _1885_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_CLK clkbuf_0_CLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_CLK/A sky130_fd_sc_hd__clkbuf_2
X_2760_ _2760_/A vssd1 vssd1 vccd1 vccd1 _2769_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2691_ _1443_/C _1618_/X _2686_/X _1564_/Y vssd1 vssd1 vccd1 vccd1 _3199_/D sky130_fd_sc_hd__o211ai_1
XFILLER_8_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2585__A2 _2585_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1711_ _1691_/X _2753_/A2 _1709_/X _1710_/X vssd1 vssd1 vccd1 vccd1 _1711_/X sky130_fd_sc_hd__a22o_1
XFILLER_6_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1642_ _1691_/A vssd1 vssd1 vccd1 vccd1 _1642_/X sky130_fd_sc_hd__clkbuf_2
X_1573_ _3202_/Q _1545_/X _1572_/Y vssd1 vssd1 vccd1 vccd1 _1573_/X sky130_fd_sc_hd__o21a_1
XANTENNA__2742__C1 _2771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3312_ _3460_/CLK _3312_/D vssd1 vssd1 vccd1 vccd1 _3312_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _3247_/CLK _3243_/D vssd1 vssd1 vccd1 vccd1 _3243_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3174_ _3247_/CLK _3174_/D vssd1 vssd1 vccd1 vccd1 _3174_/Q sky130_fd_sc_hd__dfxtp_1
X_2125_ _3348_/Q _2111_/X _2124_/Y vssd1 vssd1 vccd1 vccd1 _2125_/X sky130_fd_sc_hd__o21a_1
XFILLER_54_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2147__B _2967_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2056_ _2056_/A vssd1 vssd1 vccd1 vccd1 _2056_/X sky130_fd_sc_hd__clkbuf_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2163__A _2163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2958_ _2958_/A _2965_/B vssd1 vssd1 vccd1 vccd1 _3351_/D sky130_fd_sc_hd__nand2_1
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1909_ _1909_/A _1917_/B _1909_/C vssd1 vssd1 vccd1 vccd1 _1909_/Y sky130_fd_sc_hd__nand3_1
X_2889_ _3314_/Q _2888_/X _2884_/X _2000_/Y vssd1 vssd1 vccd1 vccd1 _3314_/D sky130_fd_sc_hd__o211a_1
XFILLER_77_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2567__A2 _3149_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input87_A core_dmem_request_put[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2801__A _2878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput161 fmc_dmem_response_put[23] vssd1 vssd1 vccd1 vccd1 _3151_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput172 fmc_dmem_response_put[4] vssd1 vssd1 vccd1 vccd1 _2492_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput150 fmc_dmem_response_put[13] vssd1 vssd1 vccd1 vccd1 _3138_/A2 sky130_fd_sc_hd__clkbuf_4
XANTENNA_output508_A _2279_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput194 fmc_imem_response_put[24] vssd1 vssd1 vccd1 vccd1 _1749_/A2 sky130_fd_sc_hd__buf_2
Xinput183 fmc_imem_response_put[14] vssd1 vssd1 vccd1 vccd1 _1707_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_63_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2812_ _3275_/Q _2795_/X _1854_/Y vssd1 vssd1 vccd1 vccd1 _2813_/A sky130_fd_sc_hd__o21ai_1
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2558__A2 _3147_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2743_ _2743_/A _2743_/B vssd1 vssd1 vccd1 vccd1 _3235_/D sky130_fd_sc_hd__nor2_1
XFILLER_8_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput602 _1626_/X vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[28] sky130_fd_sc_hd__buf_2
X_2674_ _3189_/Q _2660_/X _2661_/X _1527_/Y vssd1 vssd1 vccd1 vccd1 _3189_/D sky130_fd_sc_hd__o211a_1
Xoutput613 _1575_/Y vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[9] sky130_fd_sc_hd__buf_2
X_1625_ _1605_/X _1606_/X _1607_/X _1527_/C _1443_/A vssd1 vssd1 vccd1 vccd1 _1625_/Y
+ sky130_fd_sc_hd__o311ai_4
X_1556_ _1546_/X _1547_/X _1548_/X _1432_/C _1527_/A vssd1 vssd1 vccd1 vccd1 _1556_/Y
+ sky130_fd_sc_hd__o311ai_4
X_1487_ _1487_/A vssd1 vssd1 vccd1 vccd1 _1488_/C sky130_fd_sc_hd__inv_2
X_3226_ _3226_/CLK _3226_/D vssd1 vssd1 vccd1 vccd1 _3226_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3157_ _3489_/CLK _3157_/D vssd1 vssd1 vccd1 vccd1 _3157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2108_ _2108_/A vssd1 vssd1 vccd1 vccd1 _2109_/C sky130_fd_sc_hd__inv_2
XFILLER_82_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2506__B_N _2478_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3088_ _2084_/C _3077_/X _3081_/X _2403_/Y vssd1 vssd1 vccd1 vccd1 _3438_/D sky130_fd_sc_hd__o211ai_1
XANTENNA__2246__A1 _1877_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2039_ _2039_/A vssd1 vssd1 vccd1 vccd1 _2040_/C sky130_fd_sc_hd__inv_2
XFILLER_35_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2605__B _2605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2621__A _2677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input239_A ram_dmem_response_put[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input141_A core_imem_request_put[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_13_CLK_A clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_28_CLK_A clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2531__A _2531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output360_A _1870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1410_ _3160_/Q vssd1 vssd1 vccd1 vccd1 _3490_/A sky130_fd_sc_hd__inv_6
XFILLER_5_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output458_A _1489_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2390_ _2062_/C _2369_/X _2389_/Y vssd1 vssd1 vccd1 vccd1 _2390_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_95_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3011_ _1877_/C _3005_/X _3010_/X _2245_/Y vssd1 vssd1 vccd1 vccd1 _3382_/D sky130_fd_sc_hd__o211ai_1
XFILLER_64_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2726_ _3224_/Q vssd1 vssd1 vccd1 vccd1 _2726_/Y sky130_fd_sc_hd__inv_2
XANTENNA__2400__A1 _2077_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput410 _2037_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[64] sky130_fd_sc_hd__buf_2
X_2657_ _3180_/Q _2644_/X _1496_/Y vssd1 vssd1 vccd1 vccd1 _2659_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__2951__A2 _2950_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput443 _2144_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[94] sky130_fd_sc_hd__buf_2
Xoutput432 _2110_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[84] sky130_fd_sc_hd__buf_2
Xoutput421 _2073_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[74] sky130_fd_sc_hd__buf_2
X_1608_ _1605_/X _1606_/X _1607_/X _1500_/C _1594_/X vssd1 vssd1 vccd1 vccd1 _1608_/Y
+ sky130_fd_sc_hd__o311ai_4
Xoutput487 _2223_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[14] sky130_fd_sc_hd__buf_2
X_2588_ _2588_/A _2556_/X vssd1 vssd1 vccd1 vccd1 _2588_/X sky130_fd_sc_hd__or2b_1
Xoutput476 _1439_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[4] sky130_fd_sc_hd__buf_2
Xoutput454 _1474_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[13] sky130_fd_sc_hd__buf_2
Xoutput465 _1510_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[23] sky130_fd_sc_hd__buf_2
Xoutput498 _2252_/X vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[24] sky130_fd_sc_hd__buf_2
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1539_ _1530_/X _2725_/B _1534_/X _1537_/X _3191_/Q vssd1 vssd1 vccd1 vccd1 _1539_/X
+ sky130_fd_sc_hd__o41a_4
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3209_ _3225_/CLK _3209_/D vssd1 vssd1 vccd1 vccd1 _3209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2054__C _2054_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2351__A _2351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input189_A fmc_imem_response_put[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2458__A1 _2169_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2526__A _2526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1681__A2 _1681_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1890_ _2815_/A vssd1 vssd1 vccd1 vccd1 _2794_/A sky130_fd_sc_hd__buf_2
XFILLER_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2511_ _3133_/B vssd1 vssd1 vccd1 vccd1 _2511_/Y sky130_fd_sc_hd__inv_2
X_3491_ _3491_/A vssd1 vssd1 vccd1 vccd1 _3491_/X sky130_fd_sc_hd__clkbuf_1
X_2442_ _2427_/X _1801_/B _3452_/Q vssd1 vssd1 vccd1 vccd1 _2442_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2373_ _2356_/X _2357_/X _2358_/X _2044_/C _2348_/X vssd1 vssd1 vccd1 vccd1 _2373_/Y
+ sky130_fd_sc_hd__o311ai_2
XFILLER_68_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3110__A2 _3105_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2709_ _2709_/A vssd1 vssd1 vccd1 vccd1 _2709_/X sky130_fd_sc_hd__clkbuf_2
Xoutput284 _1631_/X vssd1 vssd1 vccd1 vccd1 RDY_ram_imem_request_get sky130_fd_sc_hd__buf_2
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput295 _2554_/Y vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[18] sky130_fd_sc_hd__buf_2
XFILLER_87_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1663__A2 _1663_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1888__C _1888_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input104_A core_dmem_request_put[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1654__A2 _1654_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2991_ _3035_/A vssd1 vssd1 vccd1 vccd1 _2991_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1942_ _1963_/A _1971_/B _1942_/C vssd1 vssd1 vccd1 vccd1 _1942_/Y sky130_fd_sc_hd__nand3_1
XFILLER_9_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1873_ _1888_/A _1898_/B _1873_/C vssd1 vssd1 vccd1 vccd1 _1873_/Y sky130_fd_sc_hd__nand3_2
XFILLER_6_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3474_ _3476_/CLK _3474_/D vssd1 vssd1 vccd1 vccd1 _3474_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2425_ _3105_/A vssd1 vssd1 vccd1 vccd1 _3035_/A sky130_fd_sc_hd__buf_2
X_2356_ _2412_/A vssd1 vssd1 vccd1 vccd1 _2356_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2287_ _2269_/X _2270_/X _2271_/X _1935_/C _2262_/X vssd1 vssd1 vccd1 vccd1 _2287_/Y
+ sky130_fd_sc_hd__o311ai_2
XFILLER_56_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2070__A2 _2056_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input221_A ram_dmem_response_put[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3086__A1 _2077_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output440_A _2135_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _2326_/A vssd1 vssd1 vccd1 vccd1 _2210_/X sky130_fd_sc_hd__clkbuf_2
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _3197_/CLK _3190_/D vssd1 vssd1 vccd1 vccd1 _3190_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2141_ _3353_/Q _2129_/X _2140_/Y vssd1 vssd1 vccd1 vccd1 _2141_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2072_ _2072_/A _2081_/B _2072_/C vssd1 vssd1 vccd1 vccd1 _2072_/Y sky130_fd_sc_hd__nand3_1
XFILLER_81_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2974_ _3037_/A vssd1 vssd1 vccd1 vccd1 _2974_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1925_ _3293_/Q _1911_/X _1924_/Y vssd1 vssd1 vccd1 vccd1 _1925_/X sky130_fd_sc_hd__o21a_2
XANTENNA__2052__A2 _2038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1856_ _2319_/A vssd1 vssd1 vccd1 vccd1 _2006_/A sky130_fd_sc_hd__clkbuf_4
X_1787_ _2319_/A vssd1 vssd1 vccd1 vccd1 _2967_/A sky130_fd_sc_hd__clkbuf_2
X_3457_ _3457_/CLK _3457_/D vssd1 vssd1 vccd1 vccd1 _3457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3388_ _3388_/CLK _3388_/D vssd1 vssd1 vccd1 vccd1 _3388_/Q sky130_fd_sc_hd__dfxtp_1
X_2408_ _2408_/A vssd1 vssd1 vccd1 vccd1 _2408_/X sky130_fd_sc_hd__buf_2
X_2339_ _3415_/Q _2326_/X _2338_/Y vssd1 vssd1 vccd1 vccd1 _2339_/X sky130_fd_sc_hd__o21a_1
XFILLER_57_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3068__A1 _2026_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2608__B _2682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2062__C _2062_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input171_A fmc_dmem_response_put[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input269_A ram_imem_response_put[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input32_A core_dmem_request_put[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output390_A _1972_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2034__A2 _2020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2690_ _3198_/Q _2681_/X _1560_/Y _2684_/X vssd1 vssd1 vccd1 vccd1 _3198_/D sky130_fd_sc_hd__o211a_1
X_1710_ _1710_/A _1684_/X vssd1 vssd1 vccd1 vccd1 _1710_/X sky130_fd_sc_hd__or2b_1
XFILLER_6_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1641_ _1641_/A vssd1 vssd1 vccd1 vccd1 _1691_/A sky130_fd_sc_hd__buf_4
X_1572_ _1546_/X _1547_/X _1548_/X _1456_/C _1566_/X vssd1 vssd1 vccd1 vccd1 _1572_/Y
+ sky130_fd_sc_hd__o311ai_4
X_3311_ _3410_/CLK _3311_/D vssd1 vssd1 vccd1 vccd1 _3311_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ _3244_/CLK _3242_/D vssd1 vssd1 vccd1 vccd1 _3242_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__2709__A _2709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ _3482_/CLK _3173_/D vssd1 vssd1 vccd1 vccd1 _3173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2124_ _2143_/A _2152_/B _2124_/C vssd1 vssd1 vccd1 vccd1 _2124_/Y sky130_fd_sc_hd__nand3_1
XFILLER_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2055_ _3329_/Q _2038_/X _2054_/Y vssd1 vssd1 vccd1 vccd1 _2055_/X sky130_fd_sc_hd__o21a_2
XFILLER_26_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2957_ _3351_/Q _2950_/X _2134_/Y vssd1 vssd1 vccd1 vccd1 _2958_/A sky130_fd_sc_hd__o21ai_1
X_2888_ _2945_/A vssd1 vssd1 vccd1 vccd1 _2888_/X sky130_fd_sc_hd__clkbuf_2
X_1908_ _1908_/A vssd1 vssd1 vccd1 vccd1 _1909_/C sky130_fd_sc_hd__inv_2
X_1839_ _1839_/A vssd1 vssd1 vccd1 vccd1 _1840_/C sky130_fd_sc_hd__inv_4
XFILLER_89_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2619__A _2660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2016__A2 _2002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput162 fmc_dmem_response_put[24] vssd1 vssd1 vccd1 vccd1 _2578_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput140 core_imem_request_put[4] vssd1 vssd1 vccd1 vccd1 _1437_/A sky130_fd_sc_hd__clkbuf_1
Xinput151 fmc_dmem_response_put[14] vssd1 vssd1 vccd1 vccd1 _2536_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput195 fmc_imem_response_put[25] vssd1 vssd1 vccd1 vccd1 _2766_/A2 sky130_fd_sc_hd__buf_2
Xinput173 fmc_dmem_response_put[5] vssd1 vssd1 vccd1 vccd1 _3129_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput184 fmc_imem_response_put[15] vssd1 vssd1 vccd1 vccd1 _2753_/A2 sky130_fd_sc_hd__buf_2
XFILLER_91_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2811_ _3274_/Q _2810_/X _2806_/X _1850_/Y vssd1 vssd1 vccd1 vccd1 _3274_/D sky130_fd_sc_hd__o211a_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2742_ _1772_/X _2742_/A2 _1676_/X _1677_/X _2771_/A vssd1 vssd1 vccd1 vccd1 _3234_/D
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2963__B1 _2959_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2673_ _2673_/A _2673_/B vssd1 vssd1 vccd1 vccd1 _3188_/D sky130_fd_sc_hd__nand2_1
XANTENNA__3095__A _3095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput603 _1627_/X vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[29] sky130_fd_sc_hd__buf_2
X_1624_ _1523_/C _1618_/X _1623_/Y vssd1 vssd1 vccd1 vccd1 _1624_/Y sky130_fd_sc_hd__o21ai_4
X_1555_ _1429_/C _1553_/X _1554_/Y vssd1 vssd1 vccd1 vccd1 _1555_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__2191__A1 _2165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3225_ _3225_/CLK _3225_/D vssd1 vssd1 vccd1 vccd1 _3225_/Q sky130_fd_sc_hd__dfxtp_1
X_1486_ _1486_/A vssd1 vssd1 vccd1 vccd1 _1516_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2439__A _2459_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3156_ _3489_/CLK _3156_/D vssd1 vssd1 vccd1 vccd1 _3156_/Q sky130_fd_sc_hd__dfxtp_1
X_3087_ _3437_/Q _3079_/X _2401_/Y _3075_/X vssd1 vssd1 vccd1 vccd1 _3437_/D sky130_fd_sc_hd__o211a_1
XFILLER_27_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2107_ _3343_/Q _2093_/X _2106_/Y vssd1 vssd1 vccd1 vccd1 _2107_/X sky130_fd_sc_hd__o21a_2
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2038_ _2056_/A vssd1 vssd1 vccd1 vccd1 _2038_/X sky130_fd_sc_hd__buf_2
XANTENNA__2174__A _2174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2605__C input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_CLK clkbuf_0_CLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_CLK/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input134_A core_imem_request_put[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3010_ _3067_/A vssd1 vssd1 vccd1 vccd1 _3010_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2725_ _2725_/A _2725_/B vssd1 vssd1 vccd1 vccd1 _2725_/Y sky130_fd_sc_hd__nand2_1
Xoutput411 _2041_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[65] sky130_fd_sc_hd__buf_2
Xoutput400 _2005_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[55] sky130_fd_sc_hd__buf_2
X_2656_ _3179_/Q _2641_/X _2642_/X _1492_/Y vssd1 vssd1 vccd1 vccd1 _3179_/D sky130_fd_sc_hd__o211a_1
Xoutput433 _2114_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[85] sky130_fd_sc_hd__buf_2
Xoutput444 _2148_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[95] sky130_fd_sc_hd__buf_2
Xoutput422 _2078_/X vssd1 vssd1 vccd1 vccd1 fmc_dmem_request_get[75] sky130_fd_sc_hd__buf_2
X_1607_ _1607_/A vssd1 vssd1 vccd1 vccd1 _1607_/X sky130_fd_sc_hd__buf_4
Xoutput466 _1513_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[24] sky130_fd_sc_hd__buf_2
X_2587_ _2564_/X _3489_/Q _2572_/X vssd1 vssd1 vccd1 vccd1 _2587_/X sky130_fd_sc_hd__o21ba_1
Xoutput477 _1444_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[5] sky130_fd_sc_hd__buf_2
Xoutput455 _1477_/X vssd1 vssd1 vccd1 vccd1 fmc_imem_request_get[14] sky130_fd_sc_hd__buf_2
Xoutput499 _2257_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[25] sky130_fd_sc_hd__buf_2
Xoutput488 _2227_/Y vssd1 vssd1 vccd1 vccd1 ram_dmem_request_get[15] sky130_fd_sc_hd__buf_2
XFILLER_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1538_ _1530_/X _2725_/B _1534_/X _1537_/X _3190_/Q vssd1 vssd1 vccd1 vccd1 _1538_/X
+ sky130_fd_sc_hd__o41a_4
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1469_ _1469_/A vssd1 vssd1 vccd1 vccd1 _1470_/C sky130_fd_sc_hd__inv_2
XANTENNA__2169__A _2169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3208_ _3222_/CLK _3208_/D vssd1 vssd1 vccd1 vccd1 _3208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3139_ _3139_/A _3139_/B vssd1 vssd1 vccd1 vccd1 _3476_/D sky130_fd_sc_hd__nor2_1
XFILLER_94_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input251_A ram_imem_response_put[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2615__C1 _3154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output470_A _1528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3490_ _3490_/A vssd1 vssd1 vccd1 vccd1 _3490_/X sky130_fd_sc_hd__clkbuf_1
X_2510_ _2498_/X _2510_/A2 _2508_/X _2509_/X vssd1 vssd1 vccd1 vccd1 _3133_/B sky130_fd_sc_hd__a22oi_4
XANTENNA__2394__A1 _2069_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2441_ _3451_/Q _2439_/X _2440_/Y vssd1 vssd1 vccd1 vccd1 _2441_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2372_ _2040_/C _2369_/X _2371_/Y vssd1 vssd1 vccd1 vccd1 _2372_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2449__A2 _2439_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2708_ _1488_/C _2707_/X _2698_/X _1598_/Y vssd1 vssd1 vccd1 vccd1 _3211_/D sky130_fd_sc_hd__o211ai_1
XANTENNA_clkbuf_leaf_12_CLK_A clkbuf_2_2_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2639_ _2658_/A vssd1 vssd1 vccd1 vccd1 _2655_/B sky130_fd_sc_hd__clkbuf_2
Xoutput285 _3491_/X vssd1 vssd1 vccd1 vccd1 RDY_ram_imem_response_put sky130_fd_sc_hd__buf_2
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput274 _1412_/Y vssd1 vssd1 vccd1 vccd1 RDY_core_dmem_request_put sky130_fd_sc_hd__buf_2
XFILLER_59_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput296 _2558_/X vssd1 vssd1 vccd1 vccd1 core_dmem_response_get[19] sky130_fd_sc_hd__buf_2
XFILLER_87_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_27_CLK_A clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1531__A _1531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2376__A1 _2047_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input62_A core_dmem_request_put[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1706__A _1706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2990_ _3369_/Q _2974_/X _2204_/Y _2989_/X vssd1 vssd1 vccd1 vccd1 _3369_/D sky130_fd_sc_hd__o211a_1
XFILLER_61_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1941_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1942_/C sky130_fd_sc_hd__clkinv_4
X_1872_ _1872_/A vssd1 vssd1 vccd1 vccd1 _1873_/C sky130_fd_sc_hd__inv_4
XFILLER_9_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3473_ _3473_/CLK _3473_/D vssd1 vssd1 vccd1 vccd1 _3473_/Q sky130_fd_sc_hd__dfxtp_1
X_2424_ _3445_/Q _2411_/X _2423_/Y vssd1 vssd1 vccd1 vccd1 _2424_/X sky130_fd_sc_hd__o21a_1
X_2355_ _2459_/B vssd1 vssd1 vccd1 vccd1 _2355_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2286_ _1931_/C _2283_/X _2285_/Y vssd1 vssd1 vccd1 vccd1 _2286_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_56_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input214_A ram_dmem_response_put[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2597__A1 _2466_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output433_A _2114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2140_ _2169_/A _2967_/B _2140_/C vssd1 vssd1 vccd1 vccd1 _2140_/Y sky130_fd_sc_hd__nand3_1
XFILLER_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2071_ _2071_/A vssd1 vssd1 vccd1 vccd1 _2072_/C sky130_fd_sc_hd__inv_2
XFILLER_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2973_ _2973_/A vssd1 vssd1 vccd1 vccd1 _3037_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1924_ _1945_/A _1953_/B _1924_/C vssd1 vssd1 vccd1 vccd1 _1924_/Y sky130_fd_sc_hd__nand3_1
XFILLER_30_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1855_ _3275_/Q _1852_/X _1854_/Y vssd1 vssd1 vccd1 vccd1 _1855_/X sky130_fd_sc_hd__o21a_1
X_1786_ _2163_/A vssd1 vssd1 vccd1 vccd1 _2319_/A sky130_fd_sc_hd__buf_2
XFILLER_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3456_ _3456_/CLK _3456_/D vssd1 vssd1 vccd1 vccd1 _3456_/Q sky130_fd_sc_hd__dfxtp_1
X_2407_ _3439_/Q _2383_/X _2406_/Y vssd1 vssd1 vccd1 vccd1 _2407_/X sky130_fd_sc_hd__o21a_1
X_3387_ _3397_/CLK _3387_/D vssd1 vssd1 vccd1 vccd1 _3387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2338_ _2327_/X _2328_/X _2329_/X _2000_/C _2320_/X vssd1 vssd1 vccd1 vccd1 _2338_/Y
+ sky130_fd_sc_hd__o311ai_4
XFILLER_69_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2177__A _2177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2269_ _2298_/A vssd1 vssd1 vccd1 vccd1 _2269_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_84_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1512__C _1512_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2276__B1 _1920_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1554__A2 _1527_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input164_A fmc_dmem_response_put[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2087__A _2087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input25_A core_dmem_request_put[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_CLK clkbuf_2_0_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3485_/CLK sky130_fd_sc_hd__clkbuf_16
X_1640_ _2734_/B vssd1 vssd1 vccd1 vccd1 _1640_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output550_A _2390_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1571_ _1452_/C _1562_/X _1570_/Y vssd1 vssd1 vccd1 vccd1 _1571_/Y sky130_fd_sc_hd__o21ai_2
X_3310_ _3456_/CLK _3310_/D vssd1 vssd1 vccd1 vccd1 _3310_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _3241_/CLK _3241_/D vssd1 vssd1 vccd1 vccd1 _3241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3172_ _3247_/CLK _3172_/D vssd1 vssd1 vccd1 vccd1 _3172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2123_ _2123_/A vssd1 vssd1 vccd1 vccd1 _2124_/C sky130_fd_sc_hd__clkinv_2
XFILLER_39_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2258__B1 _1898_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2054_ _2054_/A _2062_/B _2054_/C vssd1 vssd1 vccd1 vccd1 _2054_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__2725__A _2725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2956_ _3350_/Q _2945_/X _2941_/X _2131_/Y vssd1 vssd1 vccd1 vccd1 _3350_/D sky130_fd_sc_hd__o211a_1
XFILLER_22_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2887_ _2887_/A _2895_/B vssd1 vssd1 vccd1 vccd1 _3313_/D sky130_fd_sc_hd__nand2_1
X_1907_ _3288_/Q _1892_/X _1906_/Y vssd1 vssd1 vccd1 vccd1 _1907_/X sky130_fd_sc_hd__o21a_2
XANTENNA__2981__A1 _1801_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1838_ _1951_/A vssd1 vssd1 vccd1 vccd1 _1869_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_35_CLK clkbuf_2_1_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3271_/CLK sky130_fd_sc_hd__clkbuf_16
X_1769_ _1769_/A _1644_/A vssd1 vssd1 vccd1 vccd1 _1769_/X sky130_fd_sc_hd__or2b_1
XFILLER_89_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3439_ _3447_/CLK _3439_/D vssd1 vssd1 vccd1 vccd1 _3439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1804__A _3116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_26_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3420_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__2370__A _2370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2972__A1 _3360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1775__A2 _2772_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1714__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput163 fmc_dmem_response_put[25] vssd1 vssd1 vccd1 vccd1 _3153_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput130 core_imem_request_put[24] vssd1 vssd1 vccd1 vccd1 _1511_/A sky130_fd_sc_hd__clkbuf_1
Xinput141 core_imem_request_put[5] vssd1 vssd1 vccd1 vccd1 _1442_/A sky130_fd_sc_hd__clkbuf_1
Xinput152 fmc_dmem_response_put[15] vssd1 vssd1 vccd1 vccd1 _3142_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput196 fmc_imem_response_put[26] vssd1 vssd1 vccd1 vccd1 _1756_/A2 sky130_fd_sc_hd__buf_2
Xinput174 fmc_dmem_response_put[6] vssd1 vssd1 vccd1 vccd1 _2503_/A2 sky130_fd_sc_hd__clkbuf_4
Xinput185 fmc_imem_response_put[16] vssd1 vssd1 vccd1 vccd1 _1717_/A2 sky130_fd_sc_hd__buf_2
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2545__A _2545_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2810_ _2868_/A vssd1 vssd1 vccd1 vccd1 _2810_/X sky130_fd_sc_hd__clkbuf_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2741_ _2743_/A _2741_/B vssd1 vssd1 vccd1 vccd1 _3233_/D sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_17_CLK clkbuf_2_3_0_CLK/X vssd1 vssd1 vccd1 vccd1 _3457_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2672_ _3188_/Q _1415_/A _1523_/Y vssd1 vssd1 vccd1 vccd1 _2673_/A sky130_fd_sc_hd__o21ai_1
Xoutput604 _1557_/X vssd1 vssd1 vccd1 vccd1 ram_imem_request_get[2] sky130_fd_sc_hd__buf_2
XANTENNA__2715__A1 _1503_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1623_ _1563_/A _1452_/B _3221_/Q vssd1 vssd1 vccd1 vccd1 _1623_/Y sky130_fd_sc_hd__o21ai_2
X_1554_ _1537_/X _1527_/B _3195_/Q vssd1 vssd1 vccd1 vccd1 _1554_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__2191__A2 _2186_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1485_ _3177_/Q _1478_/X _1484_/Y vssd1 vssd1 vccd1 vccd1 _1485_/X sky130_fd_sc_hd__o21a_2
XFILLER_86_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3224_ _3225_/CLK _3224_/D vssd1 vssd1 vccd1 vccd1 _3224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
.ends

